magic
tech gf180mcuD
magscale 1 10
timestamp 1754409076
<< metal1 >>
rect 340050 404350 340062 404402
rect 340114 404399 340126 404402
rect 343410 404399 343422 404402
rect 340114 404353 343422 404399
rect 340114 404350 340126 404353
rect 343410 404350 343422 404353
rect 343474 404350 343486 404402
rect 332434 261550 332446 261602
rect 332498 261550 332510 261602
rect 332449 261154 332495 261550
rect 332434 261102 332446 261154
rect 332498 261102 332510 261154
rect 38434 240718 38446 240770
rect 38498 240767 38510 240770
rect 40450 240767 40462 240770
rect 38498 240721 40462 240767
rect 38498 240718 38510 240721
rect 40450 240718 40462 240721
rect 40514 240718 40526 240770
rect 337810 240494 337822 240546
rect 337874 240494 337886 240546
rect 337825 240095 337871 240494
rect 337922 240095 337934 240098
rect 337825 240049 337934 240095
rect 337922 240046 337934 240049
rect 337986 240046 337998 240098
rect 301186 235790 301198 235842
rect 301250 235839 301262 235842
rect 301746 235839 301758 235842
rect 301250 235793 301758 235839
rect 301250 235790 301262 235793
rect 301746 235790 301758 235793
rect 301810 235790 301822 235842
rect 324370 209806 324382 209858
rect 324434 209855 324446 209858
rect 324706 209855 324718 209858
rect 324434 209809 324718 209855
rect 324434 209806 324446 209809
rect 324706 209806 324718 209809
rect 324770 209806 324782 209858
rect 285170 160638 285182 160690
rect 285234 160687 285246 160690
rect 287298 160687 287310 160690
rect 285234 160641 287310 160687
rect 285234 160638 285246 160641
rect 287298 160638 287310 160641
rect 287362 160638 287374 160690
rect 285058 160526 285070 160578
rect 285122 160575 285134 160578
rect 289090 160575 289102 160578
rect 285122 160529 289102 160575
rect 285122 160526 285134 160529
rect 289090 160526 289102 160529
rect 289154 160526 289166 160578
<< via1 >>
rect 340062 404350 340114 404402
rect 343422 404350 343474 404402
rect 332446 261550 332498 261602
rect 332446 261102 332498 261154
rect 38446 240718 38498 240770
rect 40462 240718 40514 240770
rect 337822 240494 337874 240546
rect 337934 240046 337986 240098
rect 301198 235790 301250 235842
rect 301758 235790 301810 235842
rect 324382 209806 324434 209858
rect 324718 209806 324770 209858
rect 285182 160638 285234 160690
rect 287310 160638 287362 160690
rect 285070 160526 285122 160578
rect 289102 160526 289154 160578
<< metal2 >>
rect 11032 595672 11256 597000
rect 11004 595560 11256 595672
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 33096 595560 33348 595672
rect 4956 587188 5012 587198
rect 4956 583828 5012 587132
rect 4956 583762 5012 583772
rect 4172 390404 4228 390414
rect 4172 333396 4228 390348
rect 4172 333330 4228 333340
rect 11004 296548 11060 595560
rect 33292 590548 33348 595560
rect 33292 590482 33348 590492
rect 55132 595560 55384 595672
rect 77224 595672 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 77224 595560 77476 595672
rect 99288 595560 99540 595672
rect 52892 573076 52948 573086
rect 52892 390628 52948 573020
rect 55132 414148 55188 595560
rect 77420 588868 77476 595560
rect 99484 590660 99540 595560
rect 99484 590594 99540 590604
rect 121324 595560 121576 595672
rect 143388 595560 143640 595672
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 165480 595560 165732 595672
rect 187544 595560 187796 595672
rect 77420 588802 77476 588812
rect 121324 582148 121380 595560
rect 143388 583940 143444 595560
rect 143388 583874 143444 583884
rect 152012 590660 152068 590670
rect 121324 582082 121380 582092
rect 94892 446068 94948 446078
rect 68572 417508 68628 417518
rect 66332 417060 66388 417070
rect 55132 414082 55188 414092
rect 64092 416948 64148 416958
rect 64092 413896 64148 416892
rect 66332 413896 66388 417004
rect 68572 413896 68628 417452
rect 85260 417508 85316 417518
rect 73052 417396 73108 417406
rect 70812 417284 70868 417294
rect 70812 413896 70868 417228
rect 73052 413896 73108 417340
rect 75292 417172 75348 417182
rect 75292 413896 75348 417116
rect 85036 417172 85092 417182
rect 77532 416836 77588 416846
rect 77532 413896 77588 416780
rect 79772 416724 79828 416734
rect 79772 413896 79828 416668
rect 62076 413476 62132 413486
rect 82236 413476 82292 413486
rect 61880 413420 62076 413476
rect 82040 413420 82236 413476
rect 62076 413410 62132 413420
rect 82236 413410 82292 413420
rect 84812 413476 84868 413486
rect 52892 390562 52948 390572
rect 59612 403732 59668 403742
rect 37996 390068 38052 390078
rect 11004 296482 11060 296492
rect 20860 388164 20916 388174
rect 4172 290836 4228 290846
rect 4172 239988 4228 290780
rect 4172 239922 4228 239932
rect 13244 227780 13300 227790
rect 11340 47908 11396 47918
rect 11340 480 11396 47852
rect 13244 480 13300 227724
rect 15372 4228 15428 4238
rect 15372 480 15428 4172
rect 17276 4228 17332 4238
rect 17276 480 17332 4172
rect 19180 4228 19236 4238
rect 19180 480 19236 4172
rect 11340 392 11592 480
rect 13244 392 13496 480
rect 11368 -960 11592 392
rect 13272 -960 13496 392
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18984 392 19236 480
rect 20860 480 20916 388108
rect 24332 384132 24388 384142
rect 24332 234388 24388 384076
rect 34412 384020 34468 384030
rect 34412 276724 34468 383964
rect 34412 276658 34468 276668
rect 37996 238532 38052 390012
rect 53116 389844 53172 389854
rect 38444 384916 38500 384926
rect 37996 238466 38052 238476
rect 38220 380212 38276 380222
rect 38220 238420 38276 380156
rect 38220 238354 38276 238364
rect 38332 379988 38388 379998
rect 38332 238196 38388 379932
rect 38444 240770 38500 384860
rect 40236 384804 40292 384814
rect 38444 240718 38446 240770
rect 38498 240718 38500 240770
rect 38444 240706 38500 240718
rect 40124 380100 40180 380110
rect 40124 238308 40180 380044
rect 40124 238242 40180 238252
rect 38332 238130 38388 238140
rect 40236 237972 40292 384748
rect 44492 379652 44548 379662
rect 44492 319060 44548 379596
rect 50652 364532 50708 364542
rect 50652 360920 50708 364476
rect 53116 364532 53172 389788
rect 59612 383908 59668 403676
rect 83356 391860 83412 391870
rect 59612 383842 59668 383852
rect 69692 388276 69748 388286
rect 53116 364466 53172 364476
rect 58268 379764 58324 379774
rect 54460 362964 54516 362974
rect 54460 360920 54516 362908
rect 58268 360920 58324 379708
rect 65884 363860 65940 363870
rect 62076 363748 62132 363758
rect 62076 360920 62132 363692
rect 65884 360920 65940 363804
rect 69692 360920 69748 388220
rect 73500 386484 73556 386494
rect 73500 360920 73556 386428
rect 81116 379876 81172 379886
rect 77308 363972 77364 363982
rect 77308 360920 77364 363916
rect 81116 360920 81172 379820
rect 83356 363972 83412 391804
rect 84812 385588 84868 413420
rect 85036 393988 85092 417116
rect 85260 397348 85316 417452
rect 90076 417284 90132 417294
rect 86828 417060 86884 417070
rect 85260 397282 85316 397292
rect 86492 416724 86548 416734
rect 85036 393922 85092 393932
rect 86492 385700 86548 416668
rect 86828 392308 86884 417004
rect 88284 416948 88340 416958
rect 87276 409108 87332 409118
rect 87276 407540 87332 409052
rect 87276 407474 87332 407484
rect 86828 392242 86884 392252
rect 88172 400372 88228 400382
rect 86492 385634 86548 385644
rect 86604 391636 86660 391646
rect 84812 385522 84868 385532
rect 83356 363906 83412 363916
rect 84924 379428 84980 379438
rect 84924 360920 84980 379372
rect 86604 372988 86660 391580
rect 88172 374612 88228 400316
rect 88284 394100 88340 416892
rect 88284 394034 88340 394044
rect 90076 392420 90132 417228
rect 93324 403284 93380 403294
rect 90076 392354 90132 392364
rect 93212 397460 93268 397470
rect 89852 391636 89908 391646
rect 88172 374546 88228 374556
rect 88956 374612 89012 374622
rect 86492 372932 86660 372988
rect 88956 373828 89012 374556
rect 86492 365428 86548 372932
rect 86492 362964 86548 365372
rect 86492 360388 86548 362908
rect 88732 363972 88788 363982
rect 88732 360920 88788 363916
rect 44492 318994 44548 319004
rect 46508 360332 46872 360388
rect 46508 314188 46564 360332
rect 86492 360322 86548 360332
rect 88956 359940 89012 373772
rect 88956 359874 89012 359884
rect 46508 314132 46900 314188
rect 46844 292404 46900 314132
rect 72156 293972 72212 293982
rect 46844 290948 46900 292348
rect 46312 290892 46900 290948
rect 59052 293188 59108 293198
rect 59052 290920 59108 293132
rect 72156 290948 72212 293916
rect 71848 290892 72212 290948
rect 84588 293972 84644 293982
rect 84588 290920 84644 293916
rect 40460 240772 40516 240782
rect 40460 240770 41160 240772
rect 40460 240718 40462 240770
rect 40514 240718 41160 240770
rect 40460 240716 41160 240718
rect 40460 240706 40516 240716
rect 48300 240660 48356 240670
rect 89852 240660 89908 391580
rect 91532 388500 91588 388510
rect 89964 360388 90020 360398
rect 89964 330932 90020 360332
rect 89964 330866 90020 330876
rect 89544 240604 89908 240660
rect 48300 240594 48356 240604
rect 60844 240548 60900 240558
rect 60844 240482 60900 240492
rect 44716 240436 44772 240446
rect 44716 240370 44772 240380
rect 53676 240324 53732 240334
rect 53676 240258 53732 240268
rect 50092 240212 50148 240222
rect 50092 240146 50148 240156
rect 66220 240100 66276 240110
rect 42924 238532 42980 240072
rect 42924 238466 42980 238476
rect 46508 238420 46564 240072
rect 46508 238354 46564 238364
rect 51884 238308 51940 240072
rect 51884 238242 51940 238252
rect 55468 238196 55524 240072
rect 57260 239876 57316 240072
rect 57260 239810 57316 239820
rect 55468 238130 55524 238140
rect 40236 237906 40292 237916
rect 59052 237972 59108 240072
rect 59052 237906 59108 237916
rect 38220 236180 38276 236190
rect 24332 234322 24388 234332
rect 36876 236068 36932 236078
rect 35196 232820 35252 232830
rect 22764 232708 22820 232718
rect 22764 480 22820 232652
rect 30380 222852 30436 222862
rect 26572 219268 26628 219278
rect 24668 212548 24724 212558
rect 24668 480 24724 212492
rect 26572 480 26628 219212
rect 30380 480 30436 222796
rect 34412 222740 34468 222750
rect 33516 214228 33572 214238
rect 33516 4900 33572 214172
rect 34412 8428 34468 222684
rect 33516 4834 33572 4844
rect 34300 8372 34468 8428
rect 32508 4340 32564 4350
rect 32508 480 32564 4284
rect 34300 4340 34356 8372
rect 35196 4676 35252 232764
rect 36092 213444 36148 213454
rect 36092 121492 36148 213388
rect 36092 121426 36148 121436
rect 36876 49588 36932 236012
rect 36876 49522 36932 49532
rect 37996 229460 38052 229470
rect 35196 4610 35252 4620
rect 34300 4274 34356 4284
rect 34412 4228 34468 4238
rect 34412 480 34468 4172
rect 37996 480 38052 229404
rect 38220 49700 38276 236124
rect 41356 234612 41412 234622
rect 40012 234500 40068 234510
rect 39788 227892 39844 227902
rect 39676 222964 39732 222974
rect 38556 219492 38612 219502
rect 38444 217700 38500 217710
rect 38220 49634 38276 49644
rect 38332 214340 38388 214350
rect 38332 5012 38388 214284
rect 38332 4946 38388 4956
rect 38444 4788 38500 217644
rect 38444 4722 38500 4732
rect 38556 4228 38612 219436
rect 39676 50820 39732 222908
rect 39676 50754 39732 50764
rect 39788 50148 39844 227836
rect 39788 50082 39844 50092
rect 39900 227668 39956 227678
rect 39900 50036 39956 227612
rect 40012 51268 40068 234444
rect 41244 234388 41300 234398
rect 41020 231140 41076 231150
rect 40908 219604 40964 219614
rect 40236 214452 40292 214462
rect 40012 51202 40068 51212
rect 40124 212660 40180 212670
rect 39900 49970 39956 49980
rect 40124 4564 40180 212604
rect 40124 4498 40180 4508
rect 40236 4340 40292 214396
rect 40908 50484 40964 219548
rect 40908 50418 40964 50428
rect 41020 49924 41076 231084
rect 41020 49858 41076 49868
rect 41132 231028 41188 231038
rect 41132 49812 41188 230972
rect 41244 50708 41300 234332
rect 41244 50642 41300 50652
rect 41356 50596 41412 234556
rect 62636 233380 62692 240072
rect 64428 238420 64484 240072
rect 66220 240034 66276 240044
rect 64428 238354 64484 238364
rect 68012 237748 68068 240072
rect 69804 237860 69860 240072
rect 69804 237794 69860 237804
rect 68012 237682 68068 237692
rect 71596 237636 71652 240072
rect 73388 237972 73444 240072
rect 75180 238196 75236 240072
rect 75180 238130 75236 238140
rect 73388 237906 73444 237916
rect 71596 237570 71652 237580
rect 76972 237636 77028 240072
rect 77308 239428 77364 239438
rect 77308 238420 77364 239372
rect 77308 238354 77364 238364
rect 78764 238084 78820 240072
rect 80556 238420 80612 240072
rect 80556 238354 80612 238364
rect 78764 238018 78820 238028
rect 82348 237748 82404 240072
rect 84140 238308 84196 240072
rect 85932 239764 85988 240072
rect 85932 239698 85988 239708
rect 87724 238532 87780 240072
rect 87724 238466 87780 238476
rect 84140 238242 84196 238252
rect 82348 237682 82404 237692
rect 76972 237570 77028 237580
rect 91532 237636 91588 388444
rect 93212 367108 93268 397404
rect 92428 359940 92484 359950
rect 92428 250628 92484 359884
rect 92428 250562 92484 250572
rect 92540 330932 92596 330942
rect 92540 242004 92596 330876
rect 93212 246372 93268 367052
rect 93324 320852 93380 403228
rect 94892 397460 94948 446012
rect 94892 397394 94948 397404
rect 152012 395780 152068 590604
rect 160412 590548 160468 590558
rect 153692 583828 153748 583838
rect 153692 407092 153748 583772
rect 155372 582148 155428 582158
rect 155372 407428 155428 582092
rect 155372 407362 155428 407372
rect 153692 407026 153748 407036
rect 152012 395714 152068 395724
rect 160412 394324 160468 590492
rect 165676 590548 165732 595560
rect 186172 590996 186228 591006
rect 165676 590482 165732 590492
rect 177212 590548 177268 590558
rect 165452 588868 165508 588878
rect 163660 407540 163716 407550
rect 163100 406644 163156 406654
rect 160412 394258 160468 394268
rect 162988 405076 163044 405086
rect 99932 390180 99988 390190
rect 95116 388724 95172 388734
rect 93324 254884 93380 320796
rect 94892 388612 94948 388622
rect 93436 284788 93492 284798
rect 93436 263396 93492 284732
rect 93436 263330 93492 263340
rect 93324 254818 93380 254828
rect 93212 246306 93268 246316
rect 93324 250628 93380 250638
rect 92540 241938 92596 241948
rect 93212 242004 93268 242014
rect 91532 237570 91588 237580
rect 62636 233314 62692 233324
rect 41356 50530 41412 50540
rect 41468 219380 41524 219390
rect 41132 49746 41188 49756
rect 40236 4274 40292 4284
rect 38556 4162 38612 4172
rect 39900 4228 39956 4238
rect 39900 480 39956 4172
rect 41468 4228 41524 219324
rect 93212 217588 93268 241948
rect 93324 224308 93380 250572
rect 93324 224242 93380 224252
rect 93436 246372 93492 246382
rect 93436 222628 93492 246316
rect 94892 238308 94948 388556
rect 95116 238420 95172 388668
rect 96572 387044 96628 387054
rect 95116 238354 95172 238364
rect 95340 386708 95396 386718
rect 94892 238242 94948 238252
rect 95340 238196 95396 386652
rect 95340 238130 95396 238140
rect 96572 237860 96628 386988
rect 96796 380324 96852 380334
rect 96796 238084 96852 380268
rect 99932 238532 99988 390124
rect 99932 238466 99988 238476
rect 103292 385140 103348 385150
rect 96796 238018 96852 238028
rect 96572 237794 96628 237804
rect 103292 237748 103348 385084
rect 113484 383572 113540 383582
rect 111692 382116 111748 382126
rect 104972 381556 105028 381566
rect 104972 239876 105028 381500
rect 106652 321748 106708 321758
rect 106652 267652 106708 321692
rect 106652 267586 106708 267596
rect 104972 239810 105028 239820
rect 111692 239764 111748 382060
rect 113372 381668 113428 381678
rect 113372 240436 113428 381612
rect 113484 361396 113540 383516
rect 160412 382004 160468 382014
rect 118412 381892 118468 381902
rect 113484 361330 113540 361340
rect 116732 381780 116788 381790
rect 113372 240370 113428 240380
rect 116732 240324 116788 381724
rect 118412 240660 118468 381836
rect 147756 320068 147812 320078
rect 139244 289044 139300 289054
rect 139244 285880 139300 288988
rect 147756 285880 147812 320012
rect 156268 294868 156324 294878
rect 156268 285880 156324 294812
rect 118412 240594 118468 240604
rect 116732 240258 116788 240268
rect 160412 240212 160468 381948
rect 162092 380436 162148 380446
rect 161308 346276 161364 346286
rect 160412 240146 160468 240156
rect 160524 318276 160580 318286
rect 111692 239698 111748 239708
rect 103292 237682 103348 237692
rect 93436 222562 93492 222572
rect 93212 217522 93268 217532
rect 154924 216804 154980 216814
rect 154924 209944 154980 216748
rect 160524 216804 160580 318220
rect 161308 284788 161364 346220
rect 161308 284722 161364 284732
rect 162092 237972 162148 380380
rect 162988 342916 163044 405020
rect 163100 346276 163156 406588
rect 163660 406644 163716 407484
rect 163660 406578 163716 406588
rect 163660 406196 163716 406206
rect 163660 405076 163716 406140
rect 163660 405010 163716 405020
rect 163100 346210 163156 346220
rect 163772 386820 163828 386830
rect 163044 342860 163268 342916
rect 162988 342850 163044 342860
rect 163100 341012 163156 341022
rect 163100 339444 163156 340956
rect 163100 320852 163156 339388
rect 163100 320786 163156 320796
rect 163212 259140 163268 342860
rect 163772 341012 163828 386764
rect 163772 340946 163828 340956
rect 165452 275716 165508 588812
rect 170492 583940 170548 583950
rect 168812 404180 168868 404190
rect 167132 397572 167188 397582
rect 165564 395892 165620 395902
rect 165564 323428 165620 395836
rect 166348 366212 166404 366222
rect 166348 365428 166404 366156
rect 167132 366212 167188 397516
rect 167132 366146 167188 366156
rect 168028 367108 168084 367118
rect 165564 323362 165620 323372
rect 165676 357476 165732 357486
rect 165676 294868 165732 357420
rect 166236 355236 166292 355246
rect 166124 328356 166180 328366
rect 165676 294802 165732 294812
rect 166012 324996 166068 325006
rect 165452 275650 165508 275660
rect 163212 259074 163268 259084
rect 162092 237906 162148 237916
rect 166012 229796 166068 324940
rect 166124 231364 166180 328300
rect 166124 231298 166180 231308
rect 166012 229730 166068 229740
rect 166236 224532 166292 355180
rect 166348 329476 166404 365372
rect 167804 354116 167860 354126
rect 166348 329410 166404 329420
rect 167692 345156 167748 345166
rect 167580 327236 167636 327246
rect 167580 233156 167636 327180
rect 167580 233090 167636 233100
rect 166236 224466 166292 224476
rect 167692 223076 167748 345100
rect 167804 228004 167860 354060
rect 167804 227938 167860 227948
rect 167916 347396 167972 347406
rect 167692 223010 167748 223020
rect 167916 220948 167972 347340
rect 168028 332836 168084 367052
rect 168812 367108 168868 404124
rect 168812 367042 168868 367052
rect 169596 346276 169652 346286
rect 168028 332770 168084 332780
rect 169372 342916 169428 342926
rect 169260 323876 169316 323886
rect 168812 296548 168868 296558
rect 168812 276836 168868 296492
rect 168812 276770 168868 276780
rect 169260 234836 169316 323820
rect 169260 234770 169316 234780
rect 167916 220882 167972 220892
rect 169372 217812 169428 342860
rect 169372 217746 169428 217756
rect 169484 341796 169540 341806
rect 160524 216738 160580 216748
rect 169484 216020 169540 341740
rect 169484 215954 169540 215964
rect 169596 215908 169652 346220
rect 170492 274596 170548 583884
rect 172956 578788 173012 578798
rect 172844 577108 172900 577118
rect 172172 407652 172228 407662
rect 171388 374612 171444 374622
rect 171388 373828 171444 374556
rect 172172 374612 172228 407596
rect 172172 374546 172228 374556
rect 171276 352996 171332 353006
rect 171164 344036 171220 344046
rect 170940 339556 170996 339566
rect 170492 274530 170548 274540
rect 170828 330596 170884 330606
rect 170828 226212 170884 330540
rect 170940 228116 170996 339500
rect 170940 228050 170996 228060
rect 171052 337316 171108 337326
rect 170828 226146 170884 226156
rect 171052 223188 171108 337260
rect 171164 224644 171220 343980
rect 171276 231252 171332 352940
rect 171388 336196 171444 373772
rect 172732 348516 172788 348526
rect 171388 336130 171444 336140
rect 172396 340676 172452 340686
rect 172284 335076 172340 335086
rect 172284 233044 172340 335020
rect 172396 234724 172452 340620
rect 172620 333956 172676 333966
rect 172396 234658 172452 234668
rect 172508 329476 172564 329486
rect 172284 232978 172340 232988
rect 171276 231186 171332 231196
rect 171164 224578 171220 224588
rect 172508 223300 172564 329420
rect 172620 224868 172676 333900
rect 172732 232932 172788 348460
rect 172844 267876 172900 577052
rect 172956 268996 173012 578732
rect 177212 397236 177268 590492
rect 180012 588868 180068 588878
rect 179676 583828 179732 583838
rect 177212 397170 177268 397180
rect 179564 570500 179620 570510
rect 178892 387156 178948 387166
rect 177212 386932 177268 386942
rect 176988 383460 177044 383470
rect 176988 363748 177044 383404
rect 177212 363972 177268 386876
rect 177212 363906 177268 363916
rect 177436 383348 177492 383358
rect 177436 363860 177492 383292
rect 177884 368676 177940 368686
rect 177772 367556 177828 367566
rect 177436 363794 177492 363804
rect 177660 365316 177716 365326
rect 176988 363682 177044 363692
rect 177212 356356 177268 356366
rect 176316 350756 176372 350766
rect 176204 338436 176260 338446
rect 174524 336196 174580 336206
rect 174412 326116 174468 326126
rect 172956 268930 173012 268940
rect 174300 322756 174356 322766
rect 172844 267810 172900 267820
rect 172732 232866 172788 232876
rect 172620 224802 172676 224812
rect 172508 223234 172564 223244
rect 171052 223122 171108 223132
rect 174300 219828 174356 322700
rect 174412 221172 174468 326060
rect 174524 229684 174580 336140
rect 174524 229618 174580 229628
rect 174636 332836 174692 332846
rect 174412 221106 174468 221116
rect 174300 219762 174356 219772
rect 174636 218036 174692 332780
rect 176092 321636 176148 321646
rect 176092 228340 176148 321580
rect 176204 231476 176260 338380
rect 176204 231410 176260 231420
rect 176092 228274 176148 228284
rect 176316 219716 176372 350700
rect 177212 320068 177268 356300
rect 177212 320002 177268 320012
rect 176316 219650 176372 219660
rect 177548 251076 177604 251086
rect 174636 217970 174692 217980
rect 169596 215842 169652 215852
rect 177548 213332 177604 251020
rect 177660 239540 177716 365260
rect 177660 239474 177716 239484
rect 177772 214564 177828 367500
rect 177884 216132 177940 368620
rect 177884 216066 177940 216076
rect 177996 366436 178052 366446
rect 177772 214498 177828 214508
rect 177548 213266 177604 213276
rect 177996 212884 178052 366380
rect 178892 240100 178948 387100
rect 178892 240034 178948 240044
rect 179116 383684 179172 383694
rect 179116 239428 179172 383628
rect 179452 349636 179508 349646
rect 179116 239362 179172 239372
rect 179340 331716 179396 331726
rect 179340 228228 179396 331660
rect 179340 228162 179396 228172
rect 179452 217924 179508 349580
rect 179564 272356 179620 570444
rect 179676 273476 179732 583772
rect 179676 273410 179732 273420
rect 179564 272290 179620 272300
rect 180012 270452 180068 588812
rect 184716 572964 184772 572974
rect 183036 536452 183092 536462
rect 182252 417396 182308 417406
rect 180572 416836 180628 416846
rect 180572 385812 180628 416780
rect 182252 388948 182308 417340
rect 182364 414148 182420 414158
rect 182364 408100 182420 414092
rect 182364 408034 182420 408044
rect 183036 390852 183092 536396
rect 184604 529284 184660 529294
rect 184492 514948 184548 514958
rect 183036 390786 183092 390796
rect 183932 412020 183988 412030
rect 182252 388882 182308 388892
rect 183932 385924 183988 411964
rect 184492 392532 184548 514892
rect 184604 396004 184660 529228
rect 184716 402836 184772 572908
rect 186172 404516 186228 590940
rect 186396 590772 186452 590782
rect 186172 404450 186228 404460
rect 186284 590548 186340 590558
rect 184716 402770 184772 402780
rect 184604 395938 184660 395948
rect 186284 394660 186340 590492
rect 186284 394594 186340 394604
rect 186396 394436 186452 590716
rect 187740 590212 187796 595560
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 187740 590146 187796 590156
rect 189532 591332 189588 591342
rect 189308 576548 189364 576558
rect 188972 575092 189028 575102
rect 187964 573076 188020 573086
rect 187740 567364 187796 567374
rect 187628 557956 187684 557966
rect 187628 399140 187684 557900
rect 187740 402500 187796 567308
rect 187740 402434 187796 402444
rect 187852 565124 187908 565134
rect 187852 400708 187908 565068
rect 187964 402948 188020 573020
rect 187964 402882 188020 402892
rect 188076 569604 188132 569614
rect 187852 400642 187908 400652
rect 187628 399074 187684 399084
rect 188076 398020 188132 569548
rect 188860 566132 188916 566142
rect 188860 409444 188916 566076
rect 188972 410004 189028 575036
rect 189196 569716 189252 569726
rect 188972 409938 189028 409948
rect 189084 567140 189140 567150
rect 188860 409378 188916 409388
rect 189084 401156 189140 567084
rect 189084 401090 189140 401100
rect 189196 400932 189252 569660
rect 189308 402724 189364 576492
rect 189308 402658 189364 402668
rect 189420 574980 189476 574990
rect 189196 400866 189252 400876
rect 189420 399476 189476 574924
rect 189532 410564 189588 591276
rect 189532 410498 189588 410508
rect 189644 591108 189700 591118
rect 189644 405748 189700 591052
rect 189644 405682 189700 405692
rect 189756 590436 189812 590446
rect 189756 403844 189812 590380
rect 209580 583828 209636 595560
rect 231644 590436 231700 595560
rect 231644 590370 231700 590380
rect 253708 590212 253764 595560
rect 253708 590146 253764 590156
rect 209580 583762 209636 583772
rect 200620 573860 200676 573870
rect 198268 573748 198324 573758
rect 193788 570388 193844 570398
rect 193788 567140 193844 570332
rect 198268 569940 198324 573692
rect 200620 570388 200676 573804
rect 275772 570500 275828 595560
rect 297836 591332 297892 595560
rect 297836 591266 297892 591276
rect 319900 591220 319956 595560
rect 319900 591154 319956 591164
rect 341964 590212 342020 595560
rect 364028 591108 364084 595560
rect 364028 591042 364084 591052
rect 341964 590146 342020 590156
rect 386092 587300 386148 595560
rect 408268 588868 408324 595560
rect 430220 590996 430276 595560
rect 430220 590930 430276 590940
rect 452284 590884 452340 595560
rect 452284 590818 452340 590828
rect 408268 588802 408324 588812
rect 386092 587234 386148 587244
rect 474348 578788 474404 595560
rect 496412 590772 496468 595560
rect 496412 590706 496468 590716
rect 518476 590660 518532 595560
rect 518476 590594 518532 590604
rect 474348 578722 474404 578732
rect 540540 577108 540596 595560
rect 562604 590548 562660 595560
rect 562604 590482 562660 590492
rect 584668 587188 584724 595560
rect 584668 587122 584724 587132
rect 540540 577042 540596 577052
rect 590828 576324 590884 576334
rect 530124 574980 530180 574990
rect 529676 573076 529732 573086
rect 275772 570434 275828 570444
rect 529340 572964 529396 572974
rect 200620 570322 200676 570332
rect 252028 570388 252084 570398
rect 198268 569874 198324 569884
rect 252028 568708 252084 570332
rect 252028 568642 252084 568652
rect 193788 567074 193844 567084
rect 194012 567364 194068 567374
rect 194012 567140 194068 567308
rect 194012 567074 194068 567084
rect 189868 567028 189924 567038
rect 189868 566132 189924 566972
rect 189868 566066 189924 566076
rect 529340 448084 529396 572908
rect 529564 569828 529620 569838
rect 529340 448018 529396 448028
rect 529452 567140 529508 567150
rect 529452 443380 529508 567084
rect 529564 452788 529620 569772
rect 529676 457044 529732 573020
rect 530012 569716 530068 569726
rect 529900 568372 529956 568382
rect 529788 568260 529844 568270
rect 529788 461972 529844 568204
rect 529900 476308 529956 568316
rect 530012 480452 530068 569660
rect 530124 485156 530180 574924
rect 590604 574644 590660 574654
rect 532924 573636 532980 573646
rect 532812 573188 532868 573198
rect 532700 571732 532756 571742
rect 531132 571508 531188 571518
rect 530908 569604 530964 569614
rect 530124 485090 530180 485100
rect 530236 567252 530292 567262
rect 530124 480452 530180 480462
rect 530012 480396 530124 480452
rect 530124 480386 530180 480396
rect 529900 476242 529956 476252
rect 529788 461906 529844 461916
rect 529676 456978 529732 456988
rect 529564 452722 529620 452732
rect 529452 443314 529508 443324
rect 530236 433412 530292 567196
rect 530236 433346 530292 433356
rect 530908 419300 530964 569548
rect 531020 567028 531076 567038
rect 531020 424004 531076 566972
rect 531132 438116 531188 571452
rect 532588 569940 532644 569950
rect 532588 536900 532644 569884
rect 532588 536834 532644 536844
rect 532700 471044 532756 571676
rect 532812 499268 532868 573132
rect 532924 503972 532980 573580
rect 533372 573524 533428 573534
rect 533260 573412 533316 573422
rect 533036 571620 533092 571630
rect 533036 513380 533092 571564
rect 533148 570052 533204 570062
rect 533148 518084 533204 569996
rect 533260 522788 533316 573356
rect 533372 527492 533428 573468
rect 533372 527426 533428 527436
rect 533484 571956 533540 571966
rect 533260 522722 533316 522732
rect 533148 518018 533204 518028
rect 533036 513314 533092 513324
rect 532924 503906 532980 503916
rect 532812 499202 532868 499212
rect 532700 470978 532756 470988
rect 531132 438050 531188 438060
rect 531020 423938 531076 423948
rect 530908 419234 530964 419244
rect 533484 414596 533540 571900
rect 590492 568036 590548 568046
rect 590492 417060 590548 567980
rect 590604 443492 590660 574588
rect 590716 571396 590772 571406
rect 590716 456708 590772 571340
rect 590828 522788 590884 576268
rect 591164 574756 591220 574766
rect 590828 522722 590884 522732
rect 590940 571284 590996 571294
rect 590940 483140 590996 571228
rect 591052 567924 591108 567934
rect 591052 535892 591108 567868
rect 591164 562436 591220 574700
rect 591164 562370 591220 562380
rect 591052 535826 591108 535836
rect 590940 483074 590996 483084
rect 590716 456642 590772 456652
rect 590604 443426 590660 443436
rect 590492 416994 590548 417004
rect 591276 430164 591332 430174
rect 533484 414530 533540 414540
rect 203756 410564 203812 410574
rect 189756 403778 189812 403788
rect 192332 410004 192388 410014
rect 189420 399410 189476 399420
rect 188076 397954 188132 397964
rect 186396 394370 186452 394380
rect 192332 392644 192388 409948
rect 192444 397572 192500 410088
rect 197484 407204 197540 407214
rect 197484 398132 197540 407148
rect 197596 404180 197652 410088
rect 200732 409780 200788 409790
rect 200732 409108 200788 409724
rect 200732 409042 200788 409052
rect 202524 409444 202580 409454
rect 197596 404114 197652 404124
rect 199052 406756 199108 406766
rect 197484 398066 197540 398076
rect 199052 397796 199108 406700
rect 202412 404516 202468 404526
rect 199052 397730 199108 397740
rect 200508 398132 200564 398142
rect 192444 397506 192500 397516
rect 192332 392578 192388 392588
rect 196364 395668 196420 395678
rect 184492 392466 184548 392476
rect 183932 385858 183988 385868
rect 180572 385746 180628 385756
rect 196364 379960 196420 395612
rect 200508 389060 200564 398076
rect 200508 388994 200564 389004
rect 201068 394660 201124 394670
rect 199724 382900 199780 382910
rect 198380 382340 198436 382350
rect 197036 382228 197092 382238
rect 197036 379960 197092 382172
rect 198156 382228 198212 382238
rect 198156 379988 198212 382172
rect 197736 379932 198212 379988
rect 198380 379960 198436 382284
rect 199052 382228 199108 382238
rect 199052 379960 199108 382172
rect 199724 379960 199780 382844
rect 199948 382228 200004 382238
rect 199948 379988 200004 382172
rect 199948 379932 200424 379988
rect 201068 379960 201124 394604
rect 201740 394436 201796 394446
rect 201740 379960 201796 394380
rect 202412 379960 202468 404460
rect 202524 394436 202580 409388
rect 202748 407652 202804 410088
rect 202748 407586 202804 407596
rect 203084 405748 203140 405758
rect 202524 394370 202580 394380
rect 202636 397796 202692 397806
rect 202636 387268 202692 397740
rect 202636 387202 202692 387212
rect 203084 379960 203140 405692
rect 203756 379960 203812 410508
rect 480508 410564 480564 410574
rect 480564 410508 480984 410564
rect 480508 410498 480564 410508
rect 352828 410452 352884 410462
rect 339388 410340 339444 410350
rect 238028 410116 238084 410126
rect 207452 410088 207928 410116
rect 207452 410060 207956 410088
rect 206556 409780 206612 409790
rect 204988 409108 205044 409118
rect 204428 403844 204484 403854
rect 204428 379960 204484 403788
rect 204988 398132 205044 409052
rect 204988 398066 205044 398076
rect 206556 407988 206612 409724
rect 205212 397236 205268 397246
rect 205212 396508 205268 397180
rect 205212 396452 205380 396508
rect 205324 379988 205380 396452
rect 205128 379932 205380 379988
rect 205772 395780 205828 395790
rect 205772 379960 205828 395724
rect 206444 394324 206500 394334
rect 206444 379960 206500 394268
rect 206556 382228 206612 407932
rect 206556 382162 206612 382172
rect 207116 390628 207172 390638
rect 207116 379960 207172 390572
rect 207452 388052 207508 410060
rect 207900 409780 207956 410060
rect 207900 409714 207956 409724
rect 213052 406196 213108 410088
rect 213052 405860 213108 406140
rect 213052 405794 213108 405804
rect 216636 406644 216692 406654
rect 207452 387986 207508 387996
rect 209132 397460 209188 397470
rect 208236 384244 208292 384254
rect 207788 383012 207844 383022
rect 207788 379960 207844 382956
rect 208236 379764 208292 384188
rect 208908 383124 208964 383134
rect 208908 380548 208964 383068
rect 208908 380482 208964 380492
rect 209132 379960 209188 397404
rect 212492 384132 212548 384142
rect 211820 384020 211876 384030
rect 209804 383908 209860 383918
rect 209804 379960 209860 383852
rect 210476 383572 210532 383582
rect 210476 379960 210532 383516
rect 211820 379960 211876 383964
rect 212492 379960 212548 384076
rect 214508 381444 214564 381454
rect 214508 379960 214564 381388
rect 216524 381444 216580 381454
rect 215852 379988 215908 379998
rect 216524 379960 216580 381388
rect 216636 380660 216692 406588
rect 218204 406644 218260 410088
rect 218204 406578 218260 406588
rect 223356 396452 223412 410088
rect 228508 398132 228564 410088
rect 233660 407316 233716 410088
rect 233660 407250 233716 407260
rect 228508 398066 228564 398076
rect 223356 395780 223412 396396
rect 223356 395714 223412 395724
rect 229404 394436 229460 394446
rect 227612 392644 227668 392654
rect 219884 390068 219940 390078
rect 217532 389060 217588 389070
rect 217532 384692 217588 389004
rect 217532 384626 217588 384636
rect 218204 387268 218260 387278
rect 216636 380594 216692 380604
rect 217868 382676 217924 382686
rect 217868 379960 217924 382620
rect 218204 382564 218260 387212
rect 218204 382498 218260 382508
rect 219212 384916 219268 384926
rect 219212 379960 219268 384860
rect 219884 379960 219940 390012
rect 225932 384804 225988 384814
rect 225148 384692 225204 384702
rect 225148 382676 225204 384636
rect 225148 382610 225204 382620
rect 222572 382004 222628 382014
rect 221900 381892 221956 381902
rect 220556 381668 220612 381678
rect 220556 379960 220612 381612
rect 221228 380212 221284 380222
rect 221228 379960 221284 380156
rect 221900 379960 221956 381836
rect 222572 379960 222628 381948
rect 223916 381780 223972 381790
rect 223244 380548 223300 380558
rect 223244 379960 223300 380492
rect 223916 379960 223972 381724
rect 225260 381556 225316 381566
rect 224140 380100 224196 380110
rect 224140 379988 224196 380044
rect 224140 379932 224616 379988
rect 225260 379960 225316 381500
rect 225932 379960 225988 384748
rect 227612 384020 227668 392588
rect 227612 383954 227668 383964
rect 228620 387156 228676 387166
rect 227276 383796 227332 383806
rect 226604 383236 226660 383246
rect 226604 379960 226660 383180
rect 227276 379960 227332 383740
rect 227948 383684 228004 383694
rect 227948 379960 228004 383628
rect 228620 379960 228676 387100
rect 229292 385028 229348 385038
rect 229292 379960 229348 384972
rect 229404 382788 229460 394380
rect 229628 392532 229684 392542
rect 229628 382900 229684 392476
rect 237356 391636 237412 391646
rect 229852 390740 229908 390750
rect 229852 383012 229908 390684
rect 236684 390180 236740 390190
rect 233996 388724 234052 388734
rect 232652 388500 232708 388510
rect 229852 382946 229908 382956
rect 229964 387044 230020 387054
rect 229628 382834 229684 382844
rect 229404 382722 229460 382732
rect 229964 379960 230020 386988
rect 231980 386708 232036 386718
rect 230636 386596 230692 386606
rect 230636 379960 230692 386540
rect 231308 380436 231364 380446
rect 231308 379960 231364 380380
rect 231980 379960 232036 386652
rect 232652 379960 232708 388444
rect 233324 380324 233380 380334
rect 233324 379960 233380 380268
rect 233996 379960 234052 388668
rect 235340 388612 235396 388622
rect 234668 385140 234724 385150
rect 234668 379960 234724 385084
rect 235340 379960 235396 388556
rect 236012 382116 236068 382126
rect 236012 379960 236068 382060
rect 236684 379960 236740 390124
rect 237356 379960 237412 391580
rect 238028 379960 238084 410060
rect 238812 409332 238868 410088
rect 238812 409266 238868 409276
rect 238700 409220 238756 409230
rect 238700 379960 238756 409164
rect 243964 406532 244020 410088
rect 249116 409444 249172 410088
rect 249116 409378 249172 409388
rect 249788 409444 249844 409454
rect 249788 407652 249844 409388
rect 249788 407586 249844 407596
rect 253484 407540 253540 407550
rect 243964 406466 244020 406476
rect 252812 406756 252868 406766
rect 252140 404740 252196 404750
rect 242060 404516 242116 404526
rect 240716 402388 240772 402398
rect 240044 398020 240100 398030
rect 239372 382340 239428 382350
rect 239372 379960 239428 382284
rect 240044 379960 240100 397964
rect 240716 379960 240772 402332
rect 241388 401156 241444 401166
rect 241388 379960 241444 401100
rect 242060 379960 242116 404460
rect 244076 403956 244132 403966
rect 243404 383908 243460 383918
rect 242732 382004 242788 382014
rect 242732 379960 242788 381948
rect 243404 379960 243460 383852
rect 244076 379960 244132 403900
rect 250796 402948 250852 402958
rect 248108 402836 248164 402846
rect 246764 402500 246820 402510
rect 244748 399140 244804 399150
rect 244748 379960 244804 399084
rect 245420 397908 245476 397918
rect 245420 379960 245476 397852
rect 246092 382116 246148 382126
rect 246092 379960 246148 382060
rect 246764 379960 246820 402444
rect 247436 402500 247492 402510
rect 247436 379960 247492 402444
rect 248108 379960 248164 402780
rect 249452 401044 249508 401054
rect 248780 392532 248836 392542
rect 248780 379960 248836 392476
rect 249452 379960 249508 400988
rect 250124 395892 250180 395902
rect 250124 379960 250180 395836
rect 250796 379960 250852 402892
rect 251468 382900 251524 382910
rect 251468 379960 251524 382844
rect 252140 379960 252196 404684
rect 252812 379960 252868 406700
rect 253484 379960 253540 407484
rect 253708 407540 253764 407550
rect 253708 407204 253764 407484
rect 254268 407540 254324 410088
rect 259420 409556 259476 410088
rect 259420 409332 259476 409500
rect 259420 409266 259476 409276
rect 261996 409332 262052 409342
rect 261548 407876 261604 407886
rect 254268 407474 254324 407484
rect 254828 407764 254884 407774
rect 253708 407138 253764 407148
rect 254156 382788 254212 382798
rect 254156 379960 254212 382732
rect 254828 379960 254884 407708
rect 255500 404740 255556 404750
rect 255500 379960 255556 404684
rect 256172 404628 256228 404638
rect 256172 379960 256228 404572
rect 259532 404628 259588 404638
rect 257516 400932 257572 400942
rect 256844 392644 256900 392654
rect 256844 379960 256900 392588
rect 257516 379960 257572 400876
rect 258860 399476 258916 399486
rect 258188 392756 258244 392766
rect 258188 379960 258244 392700
rect 258860 379960 258916 399420
rect 259532 379960 259588 404572
rect 260204 402724 260260 402734
rect 260204 379960 260260 402668
rect 260876 381668 260932 381678
rect 260876 379960 260932 381612
rect 261548 379960 261604 407820
rect 261996 407764 262052 409276
rect 264572 407988 264628 410088
rect 268828 410060 269752 410116
rect 264572 407922 264628 407932
rect 264908 409108 264964 409118
rect 261996 407698 262052 407708
rect 264236 404852 264292 404862
rect 262892 404068 262948 404078
rect 262220 382004 262276 382014
rect 262220 379960 262276 381948
rect 262892 379960 262948 404012
rect 263564 382564 263620 382574
rect 263564 379960 263620 382508
rect 264236 379960 264292 404796
rect 264908 379960 264964 409052
rect 268716 404964 268772 404974
rect 268828 404964 268884 410060
rect 273756 410004 273812 410014
rect 273756 407988 273812 409948
rect 273756 407922 273812 407932
rect 274652 409668 274708 409678
rect 268772 404908 268884 404964
rect 271628 405748 271684 405758
rect 267596 404068 267652 404078
rect 265580 400820 265636 400830
rect 265580 379960 265636 400764
rect 266924 396004 266980 396014
rect 266252 384020 266308 384030
rect 266252 379960 266308 383964
rect 266924 379960 266980 395948
rect 267596 379960 267652 404012
rect 268716 386036 268772 404908
rect 268716 385970 268772 385980
rect 269612 404404 269668 404414
rect 268940 382676 268996 382686
rect 268268 382452 268324 382462
rect 268268 379960 268324 382396
rect 268940 379960 268996 382620
rect 269612 379960 269668 404348
rect 270956 399364 271012 399374
rect 270284 382452 270340 382462
rect 270284 379960 270340 382396
rect 270956 379960 271012 399308
rect 271628 379960 271684 405692
rect 272972 405300 273028 405310
rect 272300 397796 272356 397806
rect 272300 379960 272356 397740
rect 272972 379960 273028 405244
rect 273644 404180 273700 404190
rect 273644 379960 273700 404124
rect 274316 397460 274372 397470
rect 274316 379960 274372 397404
rect 274652 383236 274708 409612
rect 274876 409668 274932 410088
rect 274876 409602 274932 409612
rect 277228 407428 277284 407438
rect 274652 380660 274708 383180
rect 274652 380594 274708 380604
rect 274988 404292 275044 404302
rect 274988 379960 275044 404236
rect 276332 397684 276388 397694
rect 275660 396004 275716 396014
rect 275660 379960 275716 395948
rect 276332 379960 276388 397628
rect 277228 396508 277284 407372
rect 280028 407428 280084 410088
rect 280028 407362 280084 407372
rect 284732 410060 285208 410116
rect 289884 410060 290360 410116
rect 294812 410060 295512 410116
rect 299964 410060 300664 410116
rect 310968 410088 311668 410116
rect 284732 408100 284788 410060
rect 284396 402724 284452 402734
rect 281708 402612 281764 402622
rect 277676 400708 277732 400718
rect 277228 396452 277396 396508
rect 277228 394548 277284 394558
rect 277228 387268 277284 394492
rect 277340 390852 277396 396452
rect 277340 390516 277396 390796
rect 277340 390450 277396 390460
rect 277228 387202 277284 387212
rect 277004 382564 277060 382574
rect 277004 379960 277060 382508
rect 277676 379960 277732 400652
rect 280364 399252 280420 399262
rect 279020 397572 279076 397582
rect 278012 390852 278068 390862
rect 278012 380660 278068 390796
rect 278012 380594 278068 380604
rect 278796 382004 278852 382014
rect 278796 379988 278852 381948
rect 278376 379932 278852 379988
rect 279020 379960 279076 397516
rect 279692 397572 279748 397582
rect 279692 379960 279748 397516
rect 280364 379960 280420 399196
rect 281036 396116 281092 396126
rect 281036 379960 281092 396060
rect 281708 379960 281764 402556
rect 283724 402612 283780 402622
rect 283052 396228 283108 396238
rect 283052 379960 283108 396172
rect 283724 379960 283780 402556
rect 284396 379960 284452 402668
rect 284732 390628 284788 408044
rect 286412 408884 286468 408894
rect 284732 390562 284788 390572
rect 285068 404404 285124 404414
rect 285068 379960 285124 404348
rect 285740 399252 285796 399262
rect 285740 379960 285796 399196
rect 286412 379960 286468 408828
rect 289772 408436 289828 408446
rect 289100 399476 289156 399486
rect 287756 396340 287812 396350
rect 287084 389060 287140 389070
rect 287084 379960 287140 389004
rect 287756 379960 287812 396284
rect 288428 389172 288484 389182
rect 288428 379960 288484 389116
rect 289100 379960 289156 399420
rect 289772 379960 289828 408380
rect 289884 407092 289940 410060
rect 289884 394324 289940 407036
rect 291788 409108 291844 409118
rect 291116 402948 291172 402958
rect 289884 394258 289940 394268
rect 290444 396452 290500 396462
rect 290444 379960 290500 396396
rect 291116 379960 291172 402892
rect 291788 379960 291844 409052
rect 294812 407988 294868 410060
rect 293804 404180 293860 404190
rect 292460 392980 292516 392990
rect 292460 379960 292516 392924
rect 293132 381444 293188 381454
rect 293132 379960 293188 381388
rect 293804 379960 293860 404124
rect 294812 386148 294868 407932
rect 299964 407876 300020 410060
rect 299180 407204 299236 407214
rect 296492 405076 296548 405086
rect 294812 386082 294868 386092
rect 295148 392868 295204 392878
rect 294476 381668 294532 381678
rect 294476 379960 294532 381612
rect 295148 379960 295204 392812
rect 295820 389284 295876 389294
rect 295820 379960 295876 389228
rect 296492 379960 296548 405020
rect 297836 399588 297892 399598
rect 297164 382004 297220 382014
rect 297164 379960 297220 381948
rect 297836 379960 297892 399532
rect 298956 382004 299012 382014
rect 298956 379988 299012 381948
rect 298536 379932 299012 379988
rect 299180 379960 299236 407148
rect 299852 399700 299908 399710
rect 299852 379960 299908 399644
rect 299964 390740 300020 407820
rect 299964 390674 300020 390684
rect 302540 408660 302596 408670
rect 301196 382116 301252 382126
rect 300524 382004 300580 382014
rect 300524 379960 300580 381948
rect 301196 379960 301252 382060
rect 302204 382004 302260 382014
rect 302204 379988 302260 381948
rect 301896 379932 302260 379988
rect 302540 379960 302596 408604
rect 305788 408100 305844 410088
rect 310940 410060 311668 410088
rect 310940 409892 310996 410060
rect 310940 409826 310996 409836
rect 305788 406644 305844 408044
rect 305788 406578 305844 406588
rect 306796 406644 306852 406654
rect 305228 389844 305284 389854
rect 303212 382116 303268 382126
rect 303212 379960 303268 382060
rect 303884 382004 303940 382014
rect 303884 379960 303940 381948
rect 304556 381668 304612 381678
rect 304556 379960 304612 381612
rect 305228 379960 305284 389788
rect 306796 384020 306852 406588
rect 309260 391860 309316 391870
rect 306796 383954 306852 383964
rect 307916 388276 307972 388286
rect 306572 383460 306628 383470
rect 306572 379960 306628 383404
rect 307244 383348 307300 383358
rect 307244 379960 307300 383292
rect 307916 379960 307972 388220
rect 308588 386484 308644 386494
rect 308588 379960 308644 386428
rect 309260 379960 309316 391804
rect 311276 386932 311332 386942
rect 311276 379960 311332 386876
rect 311612 380772 311668 410060
rect 315308 397348 315364 397358
rect 313964 394100 314020 394110
rect 311612 380706 311668 380716
rect 311948 387268 312004 387278
rect 311948 379960 312004 387212
rect 312620 385924 312676 385934
rect 312620 379960 312676 385868
rect 313292 382004 313348 382014
rect 313292 379960 313348 381948
rect 313964 379960 314020 394044
rect 314636 392308 314692 392318
rect 314636 379960 314692 392252
rect 315308 379960 315364 397292
rect 315980 392420 316036 392430
rect 315980 379960 316036 392364
rect 316092 388276 316148 410088
rect 321244 396508 321300 410088
rect 321244 396452 321748 396508
rect 317324 393988 317380 393998
rect 316092 388210 316148 388220
rect 316652 388948 316708 388958
rect 316652 379960 316708 388892
rect 317324 379960 317380 393932
rect 321692 390404 321748 396452
rect 317996 385812 318052 385822
rect 317996 379960 318052 385756
rect 318668 385700 318724 385710
rect 318668 379960 318724 385644
rect 319340 385588 319396 385598
rect 319340 379960 319396 385532
rect 321692 380884 321748 390348
rect 326396 385252 326452 410088
rect 326396 385186 326452 385196
rect 329644 399924 329700 399934
rect 321692 380818 321748 380828
rect 215852 379922 215908 379932
rect 309932 379876 309988 379886
rect 309932 379810 309988 379820
rect 305900 379764 305956 379774
rect 208236 379708 208488 379764
rect 305900 379698 305956 379708
rect 211148 379652 211204 379662
rect 211148 379586 211204 379596
rect 218540 379652 218596 379662
rect 218540 379586 218596 379596
rect 190764 379540 190820 379550
rect 191324 379540 191380 379550
rect 192108 379540 192164 379550
rect 192668 379540 192724 379550
rect 190344 379484 190764 379540
rect 191016 379484 191324 379540
rect 191688 379484 192108 379540
rect 192360 379484 192668 379540
rect 190764 379474 190820 379484
rect 191324 379474 191380 379484
rect 192108 379474 192164 379484
rect 192668 379474 192724 379484
rect 193340 379540 193396 379550
rect 194684 379540 194740 379550
rect 193396 379484 193704 379540
rect 194376 379484 194684 379540
rect 193340 379474 193396 379484
rect 194684 379474 194740 379484
rect 195244 379540 195300 379550
rect 282380 379540 282436 379550
rect 195300 379484 195720 379540
rect 195244 379474 195300 379484
rect 282380 379474 282436 379484
rect 310604 379428 310660 379438
rect 310604 379362 310660 379372
rect 193004 379316 193060 379326
rect 193004 379250 193060 379260
rect 195020 379316 195076 379326
rect 195020 379250 195076 379260
rect 213164 379316 213220 379326
rect 213164 379250 213220 379260
rect 213836 379316 213892 379326
rect 213836 379250 213892 379260
rect 215180 379316 215236 379326
rect 215180 379250 215236 379260
rect 217196 379316 217252 379326
rect 217196 379250 217252 379260
rect 329532 366324 329588 366334
rect 329420 362964 329476 362974
rect 180012 270386 180068 270396
rect 180124 351316 180180 351326
rect 180124 229572 180180 351260
rect 180124 229506 180180 229516
rect 180236 293076 180292 293086
rect 179452 217858 179508 217868
rect 180236 212996 180292 293020
rect 329420 259588 329476 362908
rect 329532 308420 329588 366268
rect 329532 308354 329588 308364
rect 329644 295652 329700 399868
rect 330988 398244 331044 398254
rect 330316 395780 330372 395790
rect 330092 386036 330148 386046
rect 329756 346612 329812 346622
rect 329756 325948 329812 346556
rect 329756 325892 330036 325948
rect 329980 308980 330036 325892
rect 329980 308914 330036 308924
rect 329980 307972 330036 307982
rect 329644 295586 329700 295596
rect 329756 307412 329812 307422
rect 329420 259522 329476 259532
rect 329532 270564 329588 270574
rect 329420 242004 329476 242014
rect 327964 240548 328020 240558
rect 184940 240100 184996 240110
rect 184940 238532 184996 240044
rect 184940 238466 184996 238476
rect 185836 227780 185892 240072
rect 186396 238532 186452 238542
rect 186396 229348 186452 238476
rect 186732 232708 186788 240072
rect 186732 232642 186788 232652
rect 186396 229282 186452 229292
rect 185836 227714 185892 227724
rect 187628 222852 187684 240072
rect 188524 229460 188580 240072
rect 188524 229394 188580 229404
rect 189420 222964 189476 240072
rect 189420 222898 189476 222908
rect 187628 222786 187684 222796
rect 190316 219604 190372 240072
rect 191212 232820 191268 240072
rect 191212 232754 191268 232764
rect 190316 219538 190372 219548
rect 180236 212930 180292 212940
rect 177996 212818 178052 212828
rect 192108 212660 192164 240072
rect 193004 214452 193060 240072
rect 193900 227892 193956 240072
rect 194796 231140 194852 240072
rect 195692 234500 195748 240072
rect 196588 234612 196644 240072
rect 196588 234546 196644 234556
rect 195692 234434 195748 234444
rect 197484 234388 197540 240072
rect 198380 236180 198436 240072
rect 198380 236114 198436 236124
rect 199276 236068 199332 240072
rect 199276 236002 199332 236012
rect 200172 234500 200228 240072
rect 200172 234434 200228 234444
rect 197484 234322 197540 234332
rect 194796 231074 194852 231084
rect 193900 227826 193956 227836
rect 201068 225092 201124 240072
rect 201964 233380 202020 240072
rect 202860 233492 202916 240072
rect 202860 233426 202916 233436
rect 201964 233314 202020 233324
rect 203756 230020 203812 240072
rect 203756 229954 203812 229964
rect 201068 225026 201124 225036
rect 204652 217476 204708 240072
rect 205548 221620 205604 240072
rect 206444 224196 206500 240072
rect 207340 230132 207396 240072
rect 208236 232596 208292 240072
rect 208236 232530 208292 232540
rect 209132 231812 209188 240072
rect 209132 231746 209188 231756
rect 207340 230066 207396 230076
rect 210028 227892 210084 240072
rect 210924 228452 210980 240072
rect 210924 228386 210980 228396
rect 210028 227826 210084 227836
rect 211820 227780 211876 240072
rect 212716 229236 212772 240072
rect 213612 234612 213668 240072
rect 213612 234546 213668 234556
rect 214508 230916 214564 240072
rect 214508 230850 214564 230860
rect 212716 229170 212772 229180
rect 211820 227714 211876 227724
rect 206444 224130 206500 224140
rect 205548 221554 205604 221564
rect 204652 217410 204708 217420
rect 193004 214386 193060 214396
rect 192108 212594 192164 212604
rect 215404 212548 215460 240072
rect 216300 222740 216356 240072
rect 216300 222674 216356 222684
rect 217196 219492 217252 240072
rect 217196 219426 217252 219436
rect 218092 214340 218148 240072
rect 218092 214274 218148 214284
rect 218988 214228 219044 240072
rect 219884 217700 219940 240072
rect 220780 224420 220836 240072
rect 220780 224354 220836 224364
rect 221676 219380 221732 240072
rect 222572 227668 222628 240072
rect 223468 231028 223524 240072
rect 224364 235060 224420 240072
rect 225260 235172 225316 240072
rect 226184 240044 226772 240100
rect 226716 236964 226772 240044
rect 226716 236898 226772 236908
rect 225260 235106 225316 235116
rect 224364 234994 224420 235004
rect 223468 230962 223524 230972
rect 227052 231028 227108 240072
rect 227052 230962 227108 230972
rect 222572 227602 222628 227612
rect 227948 227556 228004 240072
rect 228844 227668 228900 240072
rect 228844 227602 228900 227612
rect 227948 227490 228004 227500
rect 229740 221732 229796 240072
rect 230636 234276 230692 240072
rect 231560 240044 231812 240100
rect 231756 236964 231812 240044
rect 231756 236898 231812 236908
rect 230636 234210 230692 234220
rect 232428 224420 232484 240072
rect 233324 236964 233380 240072
rect 234220 237076 234276 240072
rect 235116 237188 235172 240072
rect 236012 238084 236068 240072
rect 236012 238018 236068 238028
rect 235116 237122 235172 237132
rect 234220 237010 234276 237020
rect 233324 236898 233380 236908
rect 232428 224354 232484 224364
rect 229740 221666 229796 221676
rect 221676 219314 221732 219324
rect 219884 217634 219940 217644
rect 218988 214162 219044 214172
rect 236908 213108 236964 240072
rect 237804 238196 237860 240072
rect 237804 238130 237860 238140
rect 238700 237748 238756 240072
rect 239596 238420 239652 240072
rect 239596 238354 239652 238364
rect 240492 237860 240548 240072
rect 240492 237794 240548 237804
rect 238700 237682 238756 237692
rect 236908 213042 236964 213052
rect 215404 212482 215460 212492
rect 241388 210084 241444 240072
rect 242284 237972 242340 240072
rect 243180 238308 243236 240072
rect 243180 238242 243236 238252
rect 242284 237906 242340 237916
rect 244076 216692 244132 240072
rect 244972 217700 245028 240072
rect 244972 217634 245028 217644
rect 244076 216626 244132 216636
rect 245868 212548 245924 240072
rect 246764 214228 246820 240072
rect 247660 222740 247716 240072
rect 247660 222674 247716 222684
rect 248556 214340 248612 240072
rect 248556 214274 248612 214284
rect 246764 214162 246820 214172
rect 245868 212482 245924 212492
rect 249452 211204 249508 240072
rect 250348 222516 250404 240072
rect 251244 238532 251300 240072
rect 251244 238466 251300 238476
rect 252140 237636 252196 240072
rect 252140 237570 252196 237580
rect 250348 222450 250404 222460
rect 253036 211316 253092 240072
rect 253932 213220 253988 240072
rect 253932 213154 253988 213164
rect 254828 211428 254884 240072
rect 255724 213332 255780 240072
rect 256620 215796 256676 240072
rect 256620 215730 256676 215740
rect 255724 213266 255780 213276
rect 257516 211652 257572 240072
rect 258412 219380 258468 240072
rect 258412 219314 258468 219324
rect 257516 211586 257572 211596
rect 254828 211362 254884 211372
rect 253036 211250 253092 211260
rect 249452 211138 249508 211148
rect 259308 210756 259364 240072
rect 260204 219492 260260 240072
rect 260204 219426 260260 219436
rect 261100 212436 261156 240072
rect 261996 219156 262052 240072
rect 261996 219090 262052 219100
rect 261100 212370 261156 212380
rect 262892 211540 262948 240072
rect 263816 240044 264516 240100
rect 264712 240044 265412 240100
rect 265608 240044 266308 240100
rect 266504 240044 267092 240100
rect 267400 240044 268100 240100
rect 268296 240044 268660 240100
rect 269192 240044 269892 240100
rect 270088 240044 270340 240100
rect 264460 237076 264516 240044
rect 264460 237010 264516 237020
rect 265356 236964 265412 240044
rect 265356 236898 265412 236908
rect 266252 236964 266308 240044
rect 266252 236898 266308 236908
rect 267036 236964 267092 240044
rect 268044 237076 268100 240044
rect 268044 237010 268100 237020
rect 267036 236898 267092 236908
rect 268604 236964 268660 240044
rect 269836 237076 269892 240044
rect 269836 237010 269892 237020
rect 270172 239876 270228 239886
rect 268604 236898 268660 236908
rect 270172 235060 270228 239820
rect 270284 236964 270340 240044
rect 270284 236898 270340 236908
rect 270620 238196 270676 238206
rect 270172 234994 270228 235004
rect 268940 228452 268996 228462
rect 268828 227892 268884 227902
rect 262892 211474 262948 211484
rect 267932 211652 267988 211662
rect 267932 211428 267988 211596
rect 267932 211362 267988 211372
rect 259308 210690 259364 210700
rect 241388 210018 241444 210028
rect 98924 50708 98980 50718
rect 87500 50596 87556 50606
rect 53228 50484 53284 50494
rect 45612 50372 45668 50382
rect 41468 4162 41524 4172
rect 41804 5012 41860 5022
rect 41804 480 41860 4956
rect 45612 480 45668 50316
rect 49420 41188 49476 41198
rect 47516 5012 47572 5022
rect 47516 480 47572 4956
rect 49420 480 49476 41132
rect 53228 480 53284 50428
rect 76076 50148 76132 50158
rect 74172 48132 74228 48142
rect 68460 41524 68516 41534
rect 62748 41412 62804 41422
rect 57148 41300 57204 41310
rect 55132 4900 55188 4910
rect 55132 480 55188 4844
rect 57148 480 57204 41244
rect 60844 4788 60900 4798
rect 58940 4676 58996 4686
rect 58940 480 58996 4620
rect 60844 480 60900 4732
rect 62748 480 62804 41356
rect 64652 4564 64708 4574
rect 64652 480 64708 4508
rect 66556 4452 66612 4462
rect 66556 480 66612 4396
rect 68460 480 68516 41468
rect 70364 4340 70420 4350
rect 70364 480 70420 4284
rect 72268 4228 72324 4238
rect 72268 480 72324 4172
rect 74172 480 74228 48076
rect 76076 480 76132 50092
rect 77980 50036 78036 50046
rect 77980 480 78036 49980
rect 81788 49924 81844 49934
rect 79884 41636 79940 41646
rect 79884 480 79940 41580
rect 81788 480 81844 49868
rect 83692 49812 83748 49822
rect 83692 480 83748 49756
rect 85708 41748 85764 41758
rect 85708 480 85764 41692
rect 87500 480 87556 50540
rect 89404 50596 89460 50606
rect 89404 480 89460 50540
rect 93212 50484 93268 50494
rect 91308 48020 91364 48030
rect 91308 480 91364 47964
rect 93212 480 93268 50428
rect 97356 48692 97412 50120
rect 97020 48244 97076 48254
rect 95116 42868 95172 42878
rect 95116 480 95172 42812
rect 97020 480 97076 48188
rect 97356 47908 97412 48636
rect 97356 47842 97412 47852
rect 98924 480 98980 50652
rect 137004 50708 137060 50718
rect 104636 49700 104692 49710
rect 102732 47908 102788 47918
rect 100828 46228 100884 46238
rect 100828 480 100884 46172
rect 102732 480 102788 47852
rect 104636 480 104692 49644
rect 110348 49588 110404 49598
rect 108444 44548 108500 44558
rect 106540 42980 106596 42990
rect 106540 480 106596 42924
rect 108444 480 108500 44492
rect 110348 480 110404 49532
rect 114268 49588 114324 49598
rect 112252 43204 112308 43214
rect 112252 480 112308 43148
rect 114268 480 114324 49532
rect 125580 44884 125636 44894
rect 119868 44660 119924 44670
rect 116060 43092 116116 43102
rect 116060 480 116116 43036
rect 117964 39508 118020 39518
rect 117964 480 118020 39452
rect 119868 480 119924 44604
rect 123676 39620 123732 39630
rect 121772 32788 121828 32798
rect 121772 480 121828 32732
rect 123676 480 123732 39564
rect 125580 480 125636 44828
rect 131292 44772 131348 44782
rect 129388 36148 129444 36158
rect 127484 32900 127540 32910
rect 127484 480 127540 32844
rect 129388 480 129444 36092
rect 131292 480 131348 44716
rect 135100 39732 135156 39742
rect 133196 33012 133252 33022
rect 133196 480 133252 32956
rect 135100 480 135156 39676
rect 137004 480 137060 50652
rect 173180 50596 173236 50606
rect 167468 49924 167524 49934
rect 152236 49812 152292 49822
rect 150332 46340 150388 46350
rect 148428 44996 148484 45006
rect 144620 43316 144676 43326
rect 140812 36260 140868 36270
rect 138908 33124 138964 33134
rect 138908 480 138964 33068
rect 140812 480 140868 36204
rect 142828 29428 142884 29438
rect 142828 480 142884 29372
rect 144620 480 144676 43260
rect 146524 36372 146580 36382
rect 146524 480 146580 36316
rect 148428 480 148484 44940
rect 150332 480 150388 46284
rect 152236 480 152292 49756
rect 156044 49700 156100 49710
rect 154140 45108 154196 45118
rect 154140 480 154196 45052
rect 156044 480 156100 49644
rect 159852 48356 159908 48366
rect 158172 7588 158228 7598
rect 158172 480 158228 7532
rect 20860 392 21112 480
rect 22764 392 23016 480
rect 24668 392 24920 480
rect 26572 392 26824 480
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 480
rect 30380 392 30632 480
rect 30408 -960 30632 392
rect 32312 392 32564 480
rect 34216 392 34468 480
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 480
rect 37996 392 38248 480
rect 39900 392 40152 480
rect 41804 392 42056 480
rect 38024 -960 38248 392
rect 39928 -960 40152 392
rect 41832 -960 42056 392
rect 43736 -960 43960 480
rect 45612 392 45864 480
rect 47516 392 47768 480
rect 49420 392 49672 480
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 480
rect 53228 392 53480 480
rect 55132 392 55384 480
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58940 392 59192 480
rect 60844 392 61096 480
rect 62748 392 63000 480
rect 64652 392 64904 480
rect 66556 392 66808 480
rect 68460 392 68712 480
rect 70364 392 70616 480
rect 72268 392 72520 480
rect 74172 392 74424 480
rect 76076 392 76328 480
rect 77980 392 78232 480
rect 79884 392 80136 480
rect 81788 392 82040 480
rect 83692 392 83944 480
rect 58968 -960 59192 392
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 392
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 -960 85848 480
rect 87500 392 87752 480
rect 89404 392 89656 480
rect 91308 392 91560 480
rect 93212 392 93464 480
rect 95116 392 95368 480
rect 97020 392 97272 480
rect 98924 392 99176 480
rect 100828 392 101080 480
rect 102732 392 102984 480
rect 104636 392 104888 480
rect 106540 392 106792 480
rect 108444 392 108696 480
rect 110348 392 110600 480
rect 112252 392 112504 480
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 392
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 480
rect 116060 392 116312 480
rect 117964 392 118216 480
rect 119868 392 120120 480
rect 121772 392 122024 480
rect 123676 392 123928 480
rect 125580 392 125832 480
rect 127484 392 127736 480
rect 129388 392 129640 480
rect 131292 392 131544 480
rect 133196 392 133448 480
rect 135100 392 135352 480
rect 137004 392 137256 480
rect 138908 392 139160 480
rect 140812 392 141064 480
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 392
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 146524 392 146776 480
rect 148428 392 148680 480
rect 150332 392 150584 480
rect 152236 392 152488 480
rect 154140 392 154392 480
rect 156044 392 156296 480
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 392
rect 157976 392 158228 480
rect 159852 480 159908 48300
rect 161756 46452 161812 46462
rect 161756 480 161812 46396
rect 165564 26068 165620 26078
rect 163884 9268 163940 9278
rect 163884 480 163940 9212
rect 159852 392 160104 480
rect 161756 392 162008 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 392 163940 480
rect 165564 480 165620 26012
rect 167468 480 167524 49868
rect 171388 45220 171444 45230
rect 169596 4228 169652 4238
rect 169596 480 169652 4172
rect 171388 480 171444 45164
rect 173180 480 173236 50540
rect 178892 50596 178948 50606
rect 175084 41860 175140 41870
rect 175084 480 175140 41804
rect 176988 37828 177044 37838
rect 176988 480 177044 37772
rect 178892 480 178948 50540
rect 268828 50596 268884 227836
rect 268828 50530 268884 50540
rect 184604 50484 184660 50494
rect 182700 26180 182756 26190
rect 180796 19348 180852 19358
rect 180796 480 180852 19292
rect 182700 480 182756 26124
rect 184604 480 184660 50428
rect 268940 50484 268996 228396
rect 269836 222740 269892 222750
rect 269612 222516 269668 222526
rect 268940 50418 268996 50428
rect 269052 212996 269108 213006
rect 190316 50372 190372 50382
rect 188412 47684 188468 47694
rect 186508 34468 186564 34478
rect 186508 480 186564 34412
rect 188412 480 188468 47628
rect 190316 480 190372 50316
rect 196028 50372 196084 50382
rect 194124 45332 194180 45342
rect 192220 15988 192276 15998
rect 192220 480 192276 15932
rect 194124 480 194180 45276
rect 196028 480 196084 50316
rect 201740 50372 201796 50382
rect 199948 41972 200004 41982
rect 198156 4340 198212 4350
rect 198156 480 198212 4284
rect 199948 480 200004 41916
rect 201740 480 201796 50316
rect 209356 50372 209412 50382
rect 207452 48580 207508 48590
rect 205548 44436 205604 44446
rect 203644 43428 203700 43438
rect 203644 480 203700 43372
rect 205548 480 205604 44380
rect 207452 480 207508 48524
rect 209356 480 209412 50316
rect 212268 47796 212324 50120
rect 212268 47730 212324 47740
rect 269052 47796 269108 212940
rect 269500 209860 269556 209870
rect 269500 207620 269556 209804
rect 269500 207554 269556 207564
rect 269612 108724 269668 222460
rect 269836 137788 269892 222684
rect 270508 213108 270564 213118
rect 269836 137732 270004 137788
rect 269948 113540 270004 137732
rect 269948 113474 270004 113484
rect 269612 108658 269668 108668
rect 269052 47730 269108 47740
rect 211260 37940 211316 37950
rect 211260 480 211316 37884
rect 270508 4228 270564 213052
rect 270620 41860 270676 238140
rect 270844 229236 270900 229246
rect 270620 41794 270676 41804
rect 270732 221732 270788 221742
rect 270732 39620 270788 221676
rect 270844 51604 270900 229180
rect 270956 137732 271012 240072
rect 271880 240044 272132 240100
rect 272076 236964 272132 240044
rect 272076 236898 272132 236908
rect 272188 238420 272244 238430
rect 271516 234612 271572 234622
rect 271404 230916 271460 230926
rect 270956 137666 271012 137676
rect 271068 227780 271124 227790
rect 270844 51538 270900 51548
rect 271068 51492 271124 227724
rect 271292 210644 271348 210654
rect 271292 108388 271348 210588
rect 271404 190708 271460 230860
rect 271516 197428 271572 234556
rect 271516 197362 271572 197372
rect 271404 190642 271460 190652
rect 271292 108322 271348 108332
rect 271068 51426 271124 51436
rect 270732 39554 270788 39564
rect 272188 34468 272244 238364
rect 272636 237748 272692 237758
rect 272300 232820 272356 232830
rect 272300 199220 272356 232764
rect 272300 199154 272356 199164
rect 272524 210532 272580 210542
rect 272300 197428 272356 197438
rect 272300 51716 272356 197372
rect 272300 51650 272356 51660
rect 272412 190708 272468 190718
rect 272412 48580 272468 190652
rect 272524 148820 272580 210476
rect 272636 186452 272692 237692
rect 272748 211316 272804 240072
rect 273644 211652 273700 240072
rect 274568 240044 275268 240100
rect 273644 211586 273700 211596
rect 273868 237860 273924 237870
rect 272748 211250 272804 211260
rect 273196 209860 273252 209870
rect 272636 186386 272692 186396
rect 272748 209524 272804 209534
rect 272748 163380 272804 209468
rect 272860 209412 272916 209422
rect 272860 166292 272916 209356
rect 273084 209188 273140 209198
rect 272972 206388 273028 206398
rect 272972 190708 273028 206332
rect 272972 190642 273028 190652
rect 272860 166226 272916 166236
rect 272972 186004 273028 186014
rect 272748 163314 272804 163324
rect 272524 148754 272580 148764
rect 272860 121828 272916 121838
rect 272860 119700 272916 121772
rect 272860 119634 272916 119644
rect 272860 58548 272916 58558
rect 272860 51940 272916 58492
rect 272860 51874 272916 51884
rect 272972 49924 273028 185948
rect 273084 169204 273140 209132
rect 273196 175028 273252 209804
rect 273196 174962 273252 174972
rect 273420 176372 273476 176382
rect 273084 169138 273140 169148
rect 273196 143444 273252 143454
rect 273084 139076 273140 139086
rect 273084 76020 273140 139020
rect 273196 134260 273252 143388
rect 273420 143444 273476 176316
rect 273420 143378 273476 143388
rect 273196 134194 273252 134204
rect 273084 75954 273140 75964
rect 273196 91588 273252 91598
rect 273196 73108 273252 91532
rect 273196 73042 273252 73052
rect 273308 86548 273364 86558
rect 273308 70196 273364 86492
rect 273420 83188 273476 83198
rect 273420 78932 273476 83132
rect 273420 78866 273476 78876
rect 273308 70130 273364 70140
rect 273084 67284 273140 67294
rect 273084 52052 273140 67228
rect 273084 51986 273140 51996
rect 273196 64372 273252 64382
rect 273196 50372 273252 64316
rect 273196 50306 273252 50316
rect 272972 49858 273028 49868
rect 272412 48514 272468 48524
rect 272188 34402 272244 34412
rect 273868 15988 273924 237804
rect 274764 237636 274820 237646
rect 274092 233492 274148 233502
rect 273868 15922 273924 15932
rect 273980 208964 274036 208974
rect 273980 4340 274036 208908
rect 274092 33012 274148 233436
rect 274092 32946 274148 32956
rect 274204 225092 274260 225102
rect 274204 32788 274260 225036
rect 274316 224420 274372 224430
rect 274316 36260 274372 224364
rect 274428 221620 274484 221630
rect 274428 46340 274484 221564
rect 274652 211428 274708 211438
rect 274652 103348 274708 211372
rect 274764 125188 274820 237580
rect 275212 237076 275268 240044
rect 275212 237010 275268 237020
rect 275436 236964 275492 240072
rect 276360 240044 277060 240100
rect 277256 240044 277956 240100
rect 278152 240044 278740 240100
rect 275884 238308 275940 238318
rect 275436 236898 275492 236908
rect 275660 237972 275716 237982
rect 275548 233380 275604 233390
rect 274876 211652 274932 211662
rect 274876 147588 274932 211596
rect 274876 147522 274932 147532
rect 274764 125122 274820 125132
rect 274652 103282 274708 103292
rect 274652 99092 274708 99102
rect 274652 81844 274708 99036
rect 274652 81778 274708 81788
rect 274428 46274 274484 46284
rect 274316 36194 274372 36204
rect 275548 32900 275604 233324
rect 275660 43428 275716 237916
rect 275660 43362 275716 43372
rect 275772 234500 275828 234510
rect 275772 43092 275828 234444
rect 275884 51828 275940 238252
rect 277004 236964 277060 240044
rect 277900 237076 277956 240044
rect 277900 237010 277956 237020
rect 277004 236898 277060 236908
rect 278684 236964 278740 240044
rect 278684 236898 278740 236908
rect 277452 232596 277508 232606
rect 275996 231700 276052 231710
rect 275996 178500 276052 231644
rect 277228 229348 277284 229358
rect 276332 224308 276388 224318
rect 276332 204148 276388 224252
rect 276332 204082 276388 204092
rect 276444 217700 276500 217710
rect 275996 178434 276052 178444
rect 276332 197764 276388 197774
rect 275884 51762 275940 51772
rect 275772 43026 275828 43036
rect 276332 41972 276388 197708
rect 276444 106820 276500 217644
rect 276780 211204 276836 211214
rect 276444 106754 276500 106764
rect 276556 210980 276612 210990
rect 276556 103460 276612 210924
rect 276780 103908 276836 211148
rect 276780 103842 276836 103852
rect 276556 103394 276612 103404
rect 276444 61460 276500 61470
rect 276444 50260 276500 61404
rect 276444 50194 276500 50204
rect 277228 48692 277284 229292
rect 277228 48626 277284 48636
rect 277340 217476 277396 217486
rect 277340 43316 277396 217420
rect 277452 186004 277508 232540
rect 278908 230020 278964 230030
rect 278124 219492 278180 219502
rect 277452 185938 277508 185948
rect 278012 214340 278068 214350
rect 278012 104020 278068 214284
rect 278124 110292 278180 219436
rect 278348 219380 278404 219390
rect 278124 110226 278180 110236
rect 278236 213220 278292 213230
rect 278012 103954 278068 103964
rect 278236 103684 278292 213164
rect 278348 110516 278404 219324
rect 278684 211316 278740 211326
rect 278348 110450 278404 110460
rect 278460 210756 278516 210766
rect 278460 103796 278516 210700
rect 278684 148932 278740 211260
rect 278684 148866 278740 148876
rect 278460 103730 278516 103740
rect 278236 103618 278292 103628
rect 277340 43250 277396 43260
rect 276332 41906 276388 41916
rect 278908 33124 278964 229964
rect 279020 142772 279076 240072
rect 279020 142706 279076 142716
rect 279132 224196 279188 224206
rect 279132 49700 279188 224140
rect 279692 219156 279748 219166
rect 279692 108500 279748 219100
rect 279692 108434 279748 108444
rect 279804 213332 279860 213342
rect 279804 103572 279860 213276
rect 279916 160356 279972 240072
rect 280364 237972 280420 237982
rect 279916 160290 279972 160300
rect 280028 215796 280084 215806
rect 280028 110628 280084 215740
rect 280364 147028 280420 237916
rect 280476 237188 280532 237198
rect 280476 147140 280532 237132
rect 280476 147074 280532 147084
rect 280588 235956 280644 235966
rect 280364 146962 280420 146972
rect 280028 110562 280084 110572
rect 279804 103506 279860 103516
rect 280588 93492 280644 235900
rect 280812 145796 280868 240072
rect 280812 145730 280868 145740
rect 281372 239540 281428 239550
rect 280588 93426 280644 93436
rect 279132 49634 279188 49644
rect 278908 33058 278964 33068
rect 275548 32834 275604 32844
rect 274204 32722 274260 32732
rect 281372 26180 281428 239484
rect 281596 233268 281652 233278
rect 281484 231588 281540 231598
rect 281484 45332 281540 231532
rect 281484 45266 281540 45276
rect 281372 26114 281428 26124
rect 281596 26068 281652 233212
rect 281708 145684 281764 240072
rect 281708 145618 281764 145628
rect 281820 238532 281876 238542
rect 281820 128548 281876 238476
rect 282044 238196 282100 238206
rect 282044 148708 282100 238140
rect 282044 148642 282100 148652
rect 282156 237076 282212 237086
rect 282156 141988 282212 237020
rect 282156 141922 282212 141932
rect 282268 230132 282324 230142
rect 281820 128482 281876 128492
rect 282156 94052 282212 94062
rect 282156 93492 282212 93996
rect 282156 93426 282212 93436
rect 282268 46452 282324 230076
rect 282268 46386 282324 46396
rect 282380 221508 282436 221518
rect 282380 44436 282436 221452
rect 282604 145572 282660 240072
rect 282604 145506 282660 145516
rect 283052 214228 283108 214238
rect 283052 104132 283108 214172
rect 283388 199444 283444 199454
rect 283388 157556 283444 199388
rect 283388 157490 283444 157500
rect 283500 145460 283556 240072
rect 283836 236964 283892 236974
rect 283612 199668 283668 199678
rect 283612 157780 283668 199612
rect 283612 157714 283668 157724
rect 283724 199556 283780 199566
rect 283724 157332 283780 199500
rect 283724 157266 283780 157276
rect 283836 147476 283892 236908
rect 284396 152404 284452 240072
rect 284732 239764 284788 239774
rect 284620 199780 284676 199790
rect 284620 157892 284676 199724
rect 284620 157826 284676 157836
rect 284396 152338 284452 152348
rect 283836 147410 283892 147420
rect 283500 145394 283556 145404
rect 283052 104066 283108 104076
rect 284732 45108 284788 239708
rect 285068 234276 285124 234286
rect 284956 210980 285012 210990
rect 284956 160580 285012 210924
rect 284956 160514 285012 160524
rect 285068 160578 285124 234220
rect 285180 234164 285236 234174
rect 285180 160690 285236 234108
rect 285180 160638 285182 160690
rect 285234 160638 285236 160690
rect 285180 160626 285236 160638
rect 285068 160526 285070 160578
rect 285122 160526 285124 160578
rect 285068 160514 285124 160526
rect 285292 154084 285348 240072
rect 285628 240044 286216 240100
rect 285628 237636 285684 240044
rect 285404 237580 285684 237636
rect 285404 155540 285460 237580
rect 285404 155474 285460 155484
rect 285516 237412 285572 237422
rect 285292 154018 285348 154028
rect 285516 147252 285572 237356
rect 287084 237076 287140 240072
rect 287308 238756 287364 238766
rect 287308 237860 287364 238700
rect 287308 237794 287364 237804
rect 287980 237188 288036 240072
rect 287980 237122 288036 237132
rect 287084 237010 287140 237020
rect 288876 236964 288932 240072
rect 289800 240044 290500 240100
rect 288876 236898 288932 236908
rect 290444 236964 290500 240044
rect 290668 237412 290724 240072
rect 291564 237972 291620 240072
rect 291564 237906 291620 237916
rect 292460 237748 292516 240072
rect 293384 240044 293860 240100
rect 292460 237682 292516 237692
rect 290668 237346 290724 237356
rect 290444 236898 290500 236908
rect 293804 236964 293860 240044
rect 294252 238084 294308 240072
rect 295176 240044 295428 240100
rect 294252 238018 294308 238028
rect 293804 236898 293860 236908
rect 295372 236964 295428 240044
rect 296044 237972 296100 240072
rect 296044 237906 296100 237916
rect 296940 237076 296996 240072
rect 297836 238196 297892 240072
rect 298760 240044 299012 240100
rect 297836 238130 297892 238140
rect 296940 237010 296996 237020
rect 295372 236898 295428 236908
rect 298956 236964 299012 240044
rect 298956 236898 299012 236908
rect 285964 235060 286020 235070
rect 285516 147186 285572 147196
rect 285852 216692 285908 216702
rect 285852 106932 285908 216636
rect 285852 106866 285908 106876
rect 284732 45042 284788 45052
rect 282380 44370 282436 44380
rect 285964 41636 286020 235004
rect 290444 234836 290500 234846
rect 288204 228340 288260 228350
rect 288204 199864 288260 228284
rect 289324 219828 289380 219838
rect 289324 199864 289380 219772
rect 290444 199864 290500 234780
rect 293804 233156 293860 233166
rect 291564 229796 291620 229806
rect 291564 199864 291620 229740
rect 292684 221172 292740 221182
rect 292684 199864 292740 221116
rect 293804 199864 293860 233100
rect 294924 231364 294980 231374
rect 294924 199864 294980 231308
rect 298284 228228 298340 228238
rect 297164 226212 297220 226222
rect 296044 223300 296100 223310
rect 296044 199864 296100 223244
rect 297164 199864 297220 226156
rect 298284 199864 298340 228172
rect 299404 218036 299460 218046
rect 299404 199864 299460 217980
rect 299628 200004 299684 240072
rect 300300 240044 300552 240100
rect 300300 200116 300356 240044
rect 301420 238588 301476 240072
rect 301756 240044 302344 240100
rect 301420 238532 301588 238588
rect 301196 235842 301252 235854
rect 301196 235790 301198 235842
rect 301250 235790 301252 235842
rect 300300 200050 300356 200060
rect 300412 224868 300468 224878
rect 299628 199938 299684 199948
rect 300412 199892 300468 224812
rect 301196 200004 301252 235790
rect 301532 220108 301588 238532
rect 301756 235842 301812 240044
rect 301756 235790 301758 235842
rect 301810 235790 301812 235842
rect 301756 235778 301812 235790
rect 301196 199938 301252 199948
rect 301420 220052 301588 220108
rect 301644 233044 301700 233054
rect 301420 200004 301476 220052
rect 301420 199938 301476 199948
rect 300412 199836 300552 199892
rect 301644 199864 301700 232988
rect 302764 229684 302820 229694
rect 302764 199864 302820 229628
rect 303212 199444 303268 240072
rect 304108 238196 304164 240072
rect 305032 240044 305732 240100
rect 304108 238130 304164 238140
rect 305676 236964 305732 240044
rect 305900 238308 305956 240072
rect 305900 238242 305956 238252
rect 305676 236898 305732 236908
rect 305004 231476 305060 231486
rect 303884 223188 303940 223198
rect 303884 199864 303940 223132
rect 305004 199864 305060 231420
rect 306124 228116 306180 228126
rect 306124 199864 306180 228060
rect 306796 202692 306852 240072
rect 307692 238420 307748 240072
rect 307692 238354 307748 238364
rect 306796 202626 306852 202636
rect 307244 234724 307300 234734
rect 307244 199864 307300 234668
rect 308364 216020 308420 216030
rect 308364 199864 308420 215964
rect 303212 199378 303268 199388
rect 308588 199444 308644 240072
rect 309372 217812 309428 217822
rect 309372 199892 309428 217756
rect 309484 202804 309540 240072
rect 309484 202738 309540 202748
rect 309372 199836 309512 199892
rect 308588 199378 308644 199388
rect 310380 199444 310436 240072
rect 311304 240044 311892 240100
rect 310604 224644 310660 224654
rect 310604 199864 310660 224588
rect 311724 223076 311780 223086
rect 311724 199864 311780 223020
rect 310380 199378 310436 199388
rect 311836 199444 311892 240044
rect 312172 210980 312228 240072
rect 313068 234164 313124 240072
rect 313964 234276 314020 240072
rect 313964 234210 314020 234220
rect 313068 234098 313124 234108
rect 313964 220948 314020 220958
rect 312172 210914 312228 210924
rect 312844 215908 312900 215918
rect 312844 199864 312900 215852
rect 313964 199864 314020 220892
rect 314860 199780 314916 240072
rect 315084 232932 315140 232942
rect 315084 199864 315140 232876
rect 314860 199714 314916 199724
rect 315756 199668 315812 240072
rect 316204 217924 316260 217934
rect 316204 199864 316260 217868
rect 315756 199602 315812 199612
rect 316652 199556 316708 240072
rect 317324 219716 317380 219726
rect 317324 199864 317380 219660
rect 316652 199490 316708 199500
rect 311836 199378 311892 199388
rect 317548 199444 317604 240072
rect 318444 238084 318500 240072
rect 318444 238018 318500 238028
rect 318444 229572 318500 229582
rect 318444 199864 318500 229516
rect 319340 199556 319396 240072
rect 319564 231252 319620 231262
rect 319564 199864 319620 231196
rect 320236 200004 320292 240072
rect 321132 237636 321188 240072
rect 321132 237570 321188 237580
rect 320236 199938 320292 199948
rect 320684 228004 320740 228014
rect 320684 199864 320740 227948
rect 321804 224532 321860 224542
rect 321804 199864 321860 224476
rect 322028 200004 322084 240072
rect 322924 237524 322980 240072
rect 322924 237458 322980 237468
rect 322028 199938 322084 199948
rect 323820 199668 323876 240072
rect 324268 240044 324744 240100
rect 324268 236964 324324 240044
rect 325388 238420 325444 238430
rect 325164 238196 325220 238206
rect 323820 199602 323876 199612
rect 324156 236908 324324 236964
rect 324492 238084 324548 238094
rect 319340 199490 319396 199500
rect 317548 199378 317604 199388
rect 324156 198324 324212 236908
rect 324380 236516 324436 236526
rect 324380 209858 324436 236460
rect 324380 209806 324382 209858
rect 324434 209806 324436 209858
rect 324380 209794 324436 209806
rect 324492 200452 324548 238028
rect 324940 237972 324996 237982
rect 324268 200396 324548 200452
rect 324716 209858 324772 209870
rect 324716 209806 324718 209858
rect 324770 209806 324772 209858
rect 324268 199948 324324 200396
rect 324268 199892 324548 199948
rect 324156 198258 324212 198268
rect 324268 199780 324324 199790
rect 287308 160692 287364 160702
rect 287308 160690 288008 160692
rect 287308 160638 287310 160690
rect 287362 160638 288008 160690
rect 287308 160636 288008 160638
rect 287308 160626 287364 160636
rect 286188 160580 286244 160590
rect 286188 160514 286244 160524
rect 289100 160580 289156 160590
rect 289100 160578 289800 160580
rect 289100 160526 289102 160578
rect 289154 160526 289800 160578
rect 289100 160524 289800 160526
rect 289100 160514 289156 160524
rect 298060 160356 298116 160366
rect 298116 160300 298760 160356
rect 298060 160290 298116 160300
rect 307692 160244 307748 160254
rect 307692 160178 307748 160188
rect 304108 160132 304164 160142
rect 291564 157892 291620 160104
rect 291564 157826 291620 157836
rect 293356 157780 293412 160104
rect 293356 157714 293412 157724
rect 295148 157332 295204 160104
rect 296940 157556 296996 160104
rect 296940 157490 296996 157500
rect 295148 157266 295204 157276
rect 300524 157220 300580 160104
rect 302316 157780 302372 160104
rect 304108 160066 304164 160076
rect 302316 157714 302372 157724
rect 305900 157668 305956 160104
rect 309484 157892 309540 160104
rect 311276 159236 311332 160104
rect 311276 159170 311332 159180
rect 309484 157826 309540 157836
rect 305900 157602 305956 157612
rect 300524 157154 300580 157164
rect 313068 156100 313124 160104
rect 313068 156034 313124 156044
rect 314860 155988 314916 160104
rect 316652 157556 316708 160104
rect 316652 157490 316708 157500
rect 318444 156772 318500 160104
rect 320236 157444 320292 160104
rect 320236 157378 320292 157388
rect 322028 157108 322084 160104
rect 323820 157332 323876 160104
rect 324268 157780 324324 199724
rect 324380 198324 324436 198334
rect 324380 195188 324436 198268
rect 324380 195122 324436 195132
rect 324268 157714 324324 157724
rect 324492 159236 324548 199892
rect 323820 157266 323876 157276
rect 322028 157042 322084 157052
rect 324492 156996 324548 159180
rect 324604 199892 324660 199902
rect 324604 157668 324660 199836
rect 324716 192276 324772 209806
rect 324716 192210 324772 192220
rect 324604 157602 324660 157612
rect 324492 156930 324548 156940
rect 318444 156706 318500 156716
rect 314860 155922 314916 155932
rect 324940 151060 324996 237916
rect 324940 150994 324996 151004
rect 325052 212548 325108 212558
rect 324156 144116 324212 144126
rect 318556 142660 318612 142670
rect 318332 142436 318388 142446
rect 309932 142324 309988 142334
rect 308252 138852 308308 138862
rect 287756 128660 287812 128670
rect 287756 122612 287812 128604
rect 287756 122546 287812 122556
rect 308252 108052 308308 138796
rect 308252 107986 308308 107996
rect 309932 87668 309988 142268
rect 309932 87602 309988 87612
rect 311612 139188 311668 139198
rect 311612 84756 311668 139132
rect 318332 90580 318388 142380
rect 318556 96404 318612 142604
rect 323372 142548 323428 142558
rect 323372 105140 323428 142492
rect 323372 105074 323428 105084
rect 323484 122724 323540 122734
rect 318556 96338 318612 96348
rect 323484 91588 323540 122668
rect 324156 122724 324212 144060
rect 324156 122658 324212 122668
rect 325052 103236 325108 212492
rect 325164 140644 325220 238140
rect 325388 142100 325444 238364
rect 325836 237972 325892 237982
rect 325836 144452 325892 237916
rect 326732 237860 326788 237870
rect 326060 237636 326116 237646
rect 325948 237524 326004 237534
rect 325948 160244 326004 237468
rect 325948 160178 326004 160188
rect 326060 160132 326116 237580
rect 326060 160066 326116 160076
rect 326284 199668 326340 199678
rect 326284 157892 326340 199612
rect 326284 157826 326340 157836
rect 326508 199556 326564 199566
rect 326508 157220 326564 199500
rect 326508 157154 326564 157164
rect 326732 152292 326788 237804
rect 327516 237860 327572 237870
rect 327404 237748 327460 237758
rect 326844 236404 326900 236414
rect 326844 217588 326900 236348
rect 327404 231868 327460 237692
rect 327516 234948 327572 237804
rect 327516 234882 327572 234892
rect 327852 237636 327908 237646
rect 327404 231812 327572 231868
rect 326844 217522 326900 217532
rect 326956 222628 327012 222638
rect 326732 152226 326788 152236
rect 326844 198884 326900 198894
rect 326844 148820 326900 198828
rect 326956 198100 327012 222572
rect 326956 198034 327012 198044
rect 326844 148754 326900 148764
rect 327404 186452 327460 186462
rect 327404 185332 327460 186396
rect 325836 144386 325892 144396
rect 325388 142034 325444 142044
rect 325164 140578 325220 140588
rect 325052 103170 325108 103180
rect 326732 117572 326788 117582
rect 326732 116788 326788 117516
rect 327404 117572 327460 185276
rect 327516 158564 327572 231812
rect 327516 158498 327572 158508
rect 327628 188916 327684 188926
rect 327628 144116 327684 188860
rect 327852 188916 327908 237580
rect 327964 233492 328020 240492
rect 329196 240324 329252 240334
rect 329084 238756 329140 238766
rect 328972 237636 329028 237646
rect 327964 233426 328020 233436
rect 328860 237300 328916 237310
rect 328636 230244 328692 230254
rect 327852 188850 327908 188860
rect 328524 191604 328580 191614
rect 327628 144050 327684 144060
rect 328412 188132 328468 188142
rect 327404 117506 327460 117516
rect 323484 91522 323540 91532
rect 318332 90514 318388 90524
rect 326732 86548 326788 116732
rect 326732 86482 326788 86492
rect 311612 84690 311668 84700
rect 288092 55636 288148 55646
rect 288092 51828 288148 55580
rect 288092 51762 288148 51772
rect 288988 52724 289044 52734
rect 288988 51716 289044 52668
rect 288988 51650 289044 51660
rect 293580 48692 293636 50120
rect 293580 48626 293636 48636
rect 300748 47796 300804 50120
rect 307916 48468 307972 50120
rect 307916 48402 307972 48412
rect 315084 48356 315140 50120
rect 322252 48580 322308 50120
rect 322252 48514 322308 48524
rect 315084 48290 315140 48300
rect 300748 47730 300804 47740
rect 285964 41570 286020 41580
rect 281596 26002 281652 26012
rect 328412 21812 328468 188076
rect 328524 143668 328580 191548
rect 328636 186452 328692 230188
rect 328636 186386 328692 186396
rect 328524 143602 328580 143612
rect 328860 142324 328916 237244
rect 328972 236964 329028 237580
rect 328972 236898 329028 236908
rect 328860 142258 328916 142268
rect 328972 235956 329028 235966
rect 328972 138964 329028 235900
rect 328972 138898 329028 138908
rect 329084 134372 329140 238700
rect 329084 134306 329140 134316
rect 329196 23044 329252 240268
rect 329420 239876 329476 241948
rect 329420 239810 329476 239820
rect 329532 231588 329588 270508
rect 329532 231522 329588 231532
rect 329756 149492 329812 307356
rect 329980 290668 330036 307916
rect 329756 149426 329812 149436
rect 329868 290612 330036 290668
rect 329868 137620 329924 290612
rect 330092 289044 330148 385980
rect 330204 380660 330260 380670
rect 330204 301924 330260 380604
rect 330316 319172 330372 395724
rect 330652 380884 330708 380894
rect 330428 380772 330484 380782
rect 330428 341012 330484 380716
rect 330652 353892 330708 380828
rect 330652 353826 330708 353836
rect 330428 340946 330484 340956
rect 330316 319106 330372 319116
rect 330540 309204 330596 309214
rect 330204 301858 330260 301868
rect 330428 308308 330484 308318
rect 330092 288978 330148 288988
rect 330428 287364 330484 308252
rect 330428 287298 330484 287308
rect 330316 285684 330372 285694
rect 330092 260932 330148 260942
rect 330092 237748 330148 260876
rect 330092 237682 330148 237692
rect 330204 256116 330260 256126
rect 330092 236628 330148 236638
rect 329980 197876 330036 197886
rect 329980 140868 330036 197820
rect 329980 140802 330036 140812
rect 329868 137554 329924 137564
rect 330092 48020 330148 236572
rect 330204 232820 330260 256060
rect 330316 246932 330372 285628
rect 330540 277620 330596 309148
rect 330540 277554 330596 277564
rect 330652 308196 330708 308206
rect 330540 267204 330596 267214
rect 330540 263844 330596 267148
rect 330540 263778 330596 263788
rect 330316 246866 330372 246876
rect 330428 252084 330484 252094
rect 330204 232754 330260 232764
rect 330428 160132 330484 252028
rect 330428 160066 330484 160076
rect 330540 250404 330596 250414
rect 330540 138852 330596 250348
rect 330652 160020 330708 308140
rect 330988 294308 331044 398188
rect 331100 388164 331156 388174
rect 331100 308308 331156 388108
rect 331548 388052 331604 410088
rect 336588 407428 336644 407438
rect 335356 394324 335412 394334
rect 335244 390628 335300 390638
rect 331548 387986 331604 387996
rect 332556 388052 332612 388062
rect 332108 386148 332164 386158
rect 331884 382228 331940 382238
rect 331212 365092 331268 365102
rect 331212 309204 331268 365036
rect 331212 309138 331268 309148
rect 331772 361508 331828 361518
rect 331100 308242 331156 308252
rect 330988 294242 331044 294252
rect 331548 299236 331604 299246
rect 330876 289156 330932 289166
rect 330876 273364 330932 289100
rect 330988 287364 331044 287374
rect 330988 274596 331044 287308
rect 330988 274530 331044 274540
rect 330876 273298 330932 273308
rect 331548 268772 331604 299180
rect 331548 268706 331604 268716
rect 330764 263844 330820 263854
rect 330764 250740 330820 263788
rect 330876 258692 330932 258702
rect 330876 255388 330932 258636
rect 331212 257012 331268 257022
rect 330876 255332 331156 255388
rect 330764 250674 330820 250684
rect 331100 243628 331156 255332
rect 331212 248724 331268 256956
rect 331212 248658 331268 248668
rect 331660 250516 331716 250526
rect 331548 245252 331604 245262
rect 331100 243572 331268 243628
rect 330988 242116 331044 242126
rect 330988 232932 331044 242060
rect 331212 240324 331268 243572
rect 331212 240258 331268 240268
rect 331548 238644 331604 245196
rect 331660 239540 331716 250460
rect 331660 239474 331716 239484
rect 331548 238578 331604 238588
rect 330988 232866 331044 232876
rect 330652 159954 330708 159964
rect 330988 231140 331044 231150
rect 330988 142660 331044 231084
rect 330988 142594 331044 142604
rect 330540 138786 330596 138796
rect 331772 135940 331828 361452
rect 331884 297556 331940 382172
rect 331884 297490 331940 297500
rect 331996 349860 332052 349870
rect 331884 265524 331940 265534
rect 331884 256452 331940 265468
rect 331884 256386 331940 256396
rect 331772 135874 331828 135884
rect 331884 246932 331940 246942
rect 330092 47954 330148 47964
rect 329196 22978 329252 22988
rect 328412 21746 328468 21756
rect 331884 21700 331940 246876
rect 331996 157668 332052 349804
rect 332108 321412 332164 386092
rect 332556 366884 332612 387996
rect 335132 383236 335188 383246
rect 332556 366818 332612 366828
rect 334908 383124 334964 383134
rect 334572 360612 334628 360622
rect 333228 359716 333284 359726
rect 332108 321346 332164 321356
rect 332220 348068 332276 348078
rect 332108 308420 332164 308430
rect 332108 159012 332164 308364
rect 332108 158946 332164 158956
rect 331996 157602 332052 157612
rect 332220 156884 332276 348012
rect 333004 340900 333060 340910
rect 332332 338212 332388 338222
rect 332332 305620 332388 338156
rect 332332 305554 332388 305564
rect 332556 317044 332612 317054
rect 332556 298564 332612 316988
rect 332556 298498 332612 298508
rect 332668 308308 332724 308318
rect 332444 297444 332500 297454
rect 332444 283780 332500 297388
rect 332444 283714 332500 283724
rect 332556 296548 332612 296558
rect 332444 271012 332500 271022
rect 332332 264180 332388 264190
rect 332332 261492 332388 264124
rect 332444 261602 332500 270956
rect 332556 263844 332612 296492
rect 332668 288932 332724 308252
rect 332780 308084 332836 308094
rect 332780 290724 332836 308028
rect 332780 290658 332836 290668
rect 332668 288866 332724 288876
rect 332780 268324 332836 268334
rect 332780 264068 332836 268268
rect 332780 264002 332836 264012
rect 332556 263788 332836 263844
rect 332444 261550 332446 261602
rect 332498 261550 332500 261602
rect 332444 261538 332500 261550
rect 332668 262052 332724 262062
rect 332332 261426 332388 261436
rect 332556 261380 332612 261390
rect 332444 261154 332500 261166
rect 332444 261102 332446 261154
rect 332498 261102 332500 261154
rect 332332 259476 332388 259486
rect 332332 243684 332388 259420
rect 332444 254660 332500 261102
rect 332444 254594 332500 254604
rect 332556 251636 332612 261324
rect 332668 257012 332724 261996
rect 332780 258916 332836 263788
rect 332780 258850 332836 258860
rect 332668 256946 332724 256956
rect 332780 258468 332836 258478
rect 332556 251580 332724 251636
rect 332668 249956 332724 251580
rect 332668 246988 332724 249900
rect 332780 249508 332836 258412
rect 332780 249442 332836 249452
rect 332332 243618 332388 243628
rect 332556 246932 332724 246988
rect 332780 248612 332836 248622
rect 332556 242004 332612 246932
rect 332780 243460 332836 248556
rect 332780 243394 332836 243404
rect 332556 241948 332724 242004
rect 332444 240324 332500 240334
rect 332444 235956 332500 240268
rect 332668 238756 332724 241948
rect 332668 238690 332724 238700
rect 332668 238532 332724 238542
rect 332668 236516 332724 238476
rect 332668 236450 332724 236460
rect 332444 235890 332500 235900
rect 333004 157444 333060 340844
rect 333004 157378 333060 157388
rect 333116 339108 333172 339118
rect 333116 157556 333172 339052
rect 333228 307972 333284 359660
rect 333452 354340 333508 354350
rect 333340 346276 333396 346286
rect 333340 308196 333396 346220
rect 333340 308130 333396 308140
rect 333228 307906 333284 307916
rect 333452 304500 333508 354284
rect 334460 351652 334516 351662
rect 334012 342692 334068 342702
rect 333788 341796 333844 341806
rect 333452 304434 333508 304444
rect 333676 305620 333732 305630
rect 333452 292292 333508 292302
rect 333340 264740 333396 264750
rect 332220 156818 332276 156828
rect 332668 157220 332724 157230
rect 332668 156772 332724 157164
rect 332668 156706 332724 156716
rect 333116 156324 333172 157500
rect 333116 156258 333172 156268
rect 333228 243572 333284 243582
rect 333228 156100 333284 243516
rect 333340 239764 333396 264684
rect 333452 260932 333508 292236
rect 333564 273700 333620 273710
rect 333564 263844 333620 273644
rect 333564 263778 333620 263788
rect 333452 260866 333508 260876
rect 333676 258804 333732 305564
rect 333676 258738 333732 258748
rect 333564 250740 333620 250750
rect 333452 246820 333508 246830
rect 333452 243572 333508 246764
rect 333452 243506 333508 243516
rect 333340 239698 333396 239708
rect 333564 239652 333620 250684
rect 333564 239586 333620 239596
rect 333228 150948 333284 156044
rect 333228 150882 333284 150892
rect 333452 223972 333508 223982
rect 333452 183092 333508 223916
rect 332668 144340 332724 144350
rect 332668 139076 332724 144284
rect 332668 139010 332724 139020
rect 333452 136948 333508 183036
rect 333788 157108 333844 341740
rect 333900 340004 333956 340014
rect 333900 157220 333956 339948
rect 334012 157332 334068 342636
rect 334124 319172 334180 319182
rect 334124 305732 334180 319116
rect 334124 305676 334404 305732
rect 334236 303940 334292 303950
rect 334236 295652 334292 303884
rect 334348 296548 334404 305676
rect 334348 296482 334404 296492
rect 334236 295586 334292 295596
rect 334460 290668 334516 351596
rect 334572 307412 334628 360556
rect 334572 307346 334628 307356
rect 334684 336420 334740 336430
rect 334684 293972 334740 336364
rect 334796 334404 334852 334414
rect 334796 303940 334852 334348
rect 334796 303874 334852 303884
rect 334684 293906 334740 293916
rect 334796 295652 334852 295662
rect 334236 290612 334516 290668
rect 334124 283892 334180 283902
rect 334124 270452 334180 283836
rect 334236 276612 334292 290612
rect 334236 276546 334292 276556
rect 334348 283780 334404 283790
rect 334348 271012 334404 283724
rect 334796 281428 334852 295596
rect 334908 285796 334964 383068
rect 334908 285730 334964 285740
rect 335020 308980 335076 308990
rect 335020 283892 335076 308924
rect 335132 295428 335188 383180
rect 335244 308420 335300 390572
rect 335356 315812 335412 394268
rect 335468 390740 335524 390750
rect 335468 327684 335524 390684
rect 335580 384020 335636 384030
rect 335580 334404 335636 383964
rect 336588 383908 336644 407372
rect 336700 391748 336756 410088
rect 338604 410004 338660 410014
rect 338492 409668 338548 409678
rect 337484 409332 337540 409342
rect 336700 391524 336756 391692
rect 336700 391458 336756 391468
rect 336924 407876 336980 407886
rect 336588 383842 336644 383852
rect 336812 388276 336868 388286
rect 335580 334338 335636 334348
rect 336028 348964 336084 348974
rect 335468 327618 335524 327628
rect 335356 315746 335412 315756
rect 335244 308354 335300 308364
rect 335132 295362 335188 295372
rect 335244 304052 335300 304062
rect 335244 285572 335300 303996
rect 335244 285506 335300 285516
rect 335356 298564 335412 298574
rect 335020 283826 335076 283836
rect 335356 283892 335412 298508
rect 335916 297220 335972 297230
rect 335356 283826 335412 283836
rect 335468 293860 335524 293870
rect 334796 281362 334852 281372
rect 335356 282212 335412 282222
rect 334572 280868 334628 280878
rect 334572 275604 334628 280812
rect 334572 275538 334628 275548
rect 334348 270946 334404 270956
rect 334124 270386 334180 270396
rect 335132 270452 335188 270462
rect 334348 269220 334404 269230
rect 334348 258804 334404 269164
rect 334796 268996 334852 269006
rect 334236 258748 334404 258804
rect 334572 258916 334628 258926
rect 334236 250516 334292 258748
rect 334236 250450 334292 250460
rect 334012 157266 334068 157276
rect 334236 239876 334292 239886
rect 333900 157154 333956 157164
rect 333788 157042 333844 157052
rect 333900 156996 333956 157006
rect 333564 156436 333620 156446
rect 333564 155988 333620 156380
rect 333564 138964 333620 155932
rect 333676 156324 333732 156334
rect 333676 146020 333732 156268
rect 333900 147700 333956 156940
rect 334236 154420 334292 239820
rect 334572 230468 334628 258860
rect 334572 230244 334628 230412
rect 334572 230178 334628 230188
rect 334236 154354 334292 154364
rect 334796 152516 334852 268940
rect 335020 265524 335076 265534
rect 335020 259476 335076 265468
rect 335020 259410 335076 259420
rect 334908 258804 334964 258814
rect 334908 247044 334964 258748
rect 334908 246978 334964 246988
rect 335132 159572 335188 270396
rect 335356 264740 335412 282156
rect 335468 268884 335524 293804
rect 335804 289044 335860 289054
rect 335692 277508 335748 277518
rect 335468 268818 335524 268828
rect 335580 277284 335636 277294
rect 335356 264674 335412 264684
rect 335244 259588 335300 259598
rect 335244 160356 335300 259532
rect 335468 241220 335524 241230
rect 335468 238644 335524 241164
rect 335468 238578 335524 238588
rect 335244 160290 335300 160300
rect 335356 191604 335412 191614
rect 335132 159506 335188 159516
rect 335356 156436 335412 191548
rect 335580 159124 335636 277228
rect 335580 159058 335636 159068
rect 335356 156370 335412 156380
rect 335692 152628 335748 277452
rect 335804 156996 335860 288988
rect 335916 267652 335972 297164
rect 336028 292292 336084 348908
rect 336812 347396 336868 388220
rect 336924 383572 336980 407820
rect 337260 407540 337316 407550
rect 337036 406308 337092 406318
rect 337036 389284 337092 406252
rect 337036 389218 337092 389228
rect 337148 392868 337204 392878
rect 336924 379876 336980 383516
rect 336924 379810 336980 379820
rect 337036 386372 337092 386382
rect 336812 347330 336868 347340
rect 336812 341012 336868 341022
rect 336028 292226 336084 292236
rect 336700 297556 336756 297566
rect 336700 282436 336756 297500
rect 336700 282370 336756 282380
rect 335916 267586 335972 267596
rect 336028 277396 336084 277406
rect 336028 264180 336084 277340
rect 336588 275940 336644 275950
rect 336028 264114 336084 264124
rect 336140 266308 336196 266318
rect 335916 257124 335972 257134
rect 335916 250180 335972 257068
rect 335916 250114 335972 250124
rect 335916 248836 335972 248846
rect 335916 245364 335972 248780
rect 335916 245298 335972 245308
rect 336028 247044 336084 247054
rect 335916 244132 335972 244142
rect 335916 237300 335972 244076
rect 335916 237234 335972 237244
rect 336028 191604 336084 246988
rect 336140 238084 336196 266252
rect 336252 264068 336308 264078
rect 336252 253204 336308 264012
rect 336252 253138 336308 253148
rect 336140 238018 336196 238028
rect 336028 191538 336084 191548
rect 335804 156930 335860 156940
rect 335916 189812 335972 189822
rect 335692 152562 335748 152572
rect 334796 152450 334852 152460
rect 333900 147634 333956 147644
rect 333676 145954 333732 145964
rect 333564 138898 333620 138908
rect 333452 136882 333508 136892
rect 335916 22932 335972 189756
rect 336028 181412 336084 181422
rect 336028 180180 336084 181356
rect 336028 180114 336084 180124
rect 336028 178052 336084 178062
rect 336028 177044 336084 177996
rect 336028 176978 336084 176988
rect 336028 152964 336084 152974
rect 336028 144340 336084 152908
rect 336028 144274 336084 144284
rect 336588 151284 336644 275884
rect 336588 142436 336644 151228
rect 336588 142370 336644 142380
rect 336812 127652 336868 340956
rect 336924 334404 336980 334414
rect 336924 134372 336980 334348
rect 337036 214004 337092 386316
rect 337148 236404 337204 392812
rect 337260 269444 337316 407484
rect 337372 391524 337428 391534
rect 337372 373380 337428 391468
rect 337484 386372 337540 409276
rect 337484 386306 337540 386316
rect 337596 407764 337652 407774
rect 337372 373314 337428 373324
rect 337484 347396 337540 347406
rect 337260 250292 337316 269388
rect 337372 287476 337428 287486
rect 337372 265524 337428 287420
rect 337372 265458 337428 265468
rect 337260 250226 337316 250236
rect 337260 247156 337316 247166
rect 337260 237972 337316 247100
rect 337260 237906 337316 237916
rect 337148 236338 337204 236348
rect 337372 236740 337428 236750
rect 337260 224756 337316 224766
rect 337036 213938 337092 213948
rect 337148 217588 337204 217598
rect 337036 191492 337092 191502
rect 337036 168308 337092 191436
rect 337148 181412 337204 217532
rect 337260 210980 337316 224700
rect 337372 223972 337428 236684
rect 337372 223906 337428 223916
rect 337260 208348 337316 210924
rect 337260 208292 337428 208348
rect 337148 181346 337204 181356
rect 337372 178052 337428 208292
rect 337372 177986 337428 177996
rect 337036 168242 337092 168252
rect 336924 134306 336980 134316
rect 337036 144004 337092 144014
rect 337036 128660 337092 143948
rect 337484 144004 337540 347340
rect 337596 275940 337652 407708
rect 338044 406868 338100 406878
rect 338044 399588 338100 406812
rect 338044 399522 338100 399532
rect 338492 389172 338548 409612
rect 338604 399252 338660 409948
rect 338940 407652 338996 407662
rect 338604 399186 338660 399196
rect 338716 407092 338772 407102
rect 338492 389106 338548 389116
rect 338716 389060 338772 407036
rect 338716 388994 338772 389004
rect 338828 403844 338884 403854
rect 338828 382340 338884 403788
rect 338940 399140 338996 407596
rect 339164 406980 339220 406990
rect 338940 399074 338996 399084
rect 339052 403508 339108 403518
rect 339052 392532 339108 403452
rect 339164 399476 339220 406924
rect 339388 404180 339444 410284
rect 346332 410228 346388 410238
rect 340508 409220 340564 409230
rect 340284 408772 340340 408782
rect 339388 404114 339444 404124
rect 339836 405860 339892 405870
rect 339164 399410 339220 399420
rect 339276 403732 339332 403742
rect 339276 392756 339332 403676
rect 339836 396116 339892 405804
rect 340172 404964 340228 404974
rect 340060 404402 340116 404414
rect 340060 404350 340062 404402
rect 340114 404350 340116 404402
rect 340060 396228 340116 404350
rect 340060 396162 340116 396172
rect 339836 396050 339892 396060
rect 340172 393092 340228 404908
rect 340284 396452 340340 408716
rect 340284 396386 340340 396396
rect 340396 403284 340452 403294
rect 339948 393036 340228 393092
rect 339948 392980 340004 393036
rect 339948 392914 340004 392924
rect 339276 392690 339332 392700
rect 340396 392644 340452 403228
rect 340508 395892 340564 409164
rect 341852 407876 341908 410088
rect 341852 407810 341908 407820
rect 342748 407316 342804 407326
rect 340620 405188 340676 405198
rect 340620 397460 340676 405132
rect 342524 404852 342580 404862
rect 342748 404852 342804 407260
rect 342580 404796 342804 404852
rect 346332 404852 346388 410172
rect 347004 409332 347060 410088
rect 347004 409266 347060 409276
rect 352156 406756 352212 410088
rect 352828 409892 352884 410396
rect 478828 410452 478884 410462
rect 462364 410340 462420 410350
rect 352828 409826 352884 409836
rect 352940 410228 352996 410238
rect 352156 406690 352212 406700
rect 352828 409332 352884 409342
rect 352828 406644 352884 409276
rect 352940 408324 352996 410172
rect 358316 410228 358372 410238
rect 352940 408258 352996 408268
rect 352828 406578 352884 406588
rect 354732 406756 354788 406766
rect 354508 405300 354564 405310
rect 342524 404786 342580 404796
rect 346332 404786 346388 404796
rect 347564 405076 347620 405086
rect 347564 404852 347620 405020
rect 347564 404786 347620 404796
rect 343420 404404 343476 404414
rect 354508 404404 354564 405244
rect 343420 404402 344120 404404
rect 343420 404350 343422 404402
rect 343474 404350 344120 404402
rect 343420 404348 344120 404350
rect 343420 404338 343476 404348
rect 354508 404338 354564 404348
rect 354732 404404 354788 406700
rect 357308 405412 357364 410088
rect 357868 408548 357924 408558
rect 357868 406532 357924 408492
rect 358316 407652 358372 410172
rect 366156 410228 366212 410238
rect 361788 410060 362488 410116
rect 361788 410004 361844 410060
rect 361788 409938 361844 409948
rect 361452 408436 361508 408446
rect 358316 407586 358372 407596
rect 358876 407764 358932 407774
rect 357868 406466 357924 406476
rect 357308 405346 357364 405356
rect 358876 404936 358932 407708
rect 354732 404338 354788 404348
rect 361452 404404 361508 408380
rect 361452 404338 361508 404348
rect 364700 408324 364756 408334
rect 364700 404404 364756 408268
rect 366156 408100 366212 410172
rect 369628 410228 369684 410238
rect 366156 408034 366212 408044
rect 367276 407652 367332 407662
rect 367276 407316 367332 407596
rect 367276 407250 367332 407260
rect 366268 406756 366324 406766
rect 366268 404936 366324 406700
rect 367612 404964 367668 410088
rect 367612 404898 367668 404908
rect 367836 408436 367892 408446
rect 367836 404964 367892 408380
rect 369628 407764 369684 410172
rect 378812 410228 378868 410238
rect 372988 410116 373044 410126
rect 369628 407698 369684 407708
rect 372764 406644 372820 410088
rect 372988 408212 373044 410060
rect 372988 408146 373044 408156
rect 374668 408548 374724 408558
rect 372764 406578 372820 406588
rect 374668 406532 374724 408492
rect 374668 406466 374724 406476
rect 367836 404898 367892 404908
rect 377916 404516 377972 410088
rect 378812 409780 378868 410172
rect 378812 409714 378868 409724
rect 379708 410228 379764 410238
rect 379708 409108 379764 410172
rect 392252 410228 392308 410238
rect 389676 410116 389732 410126
rect 383096 410060 383236 410116
rect 379708 409042 379764 409052
rect 381052 408884 381108 408894
rect 381052 404936 381108 408828
rect 382172 408548 382228 408558
rect 382172 407540 382228 408492
rect 382172 407474 382228 407484
rect 383068 407540 383124 407550
rect 383068 406420 383124 407484
rect 383180 407428 383236 410060
rect 383180 407362 383236 407372
rect 383292 408772 383348 408782
rect 383292 406532 383348 408716
rect 384748 408324 384804 408334
rect 384748 407652 384804 408268
rect 388220 408100 388276 410088
rect 388220 408034 388276 408044
rect 384748 407586 384804 407596
rect 389676 407428 389732 410060
rect 389676 407362 389732 407372
rect 383292 406466 383348 406476
rect 388444 407092 388500 407102
rect 383068 406354 383124 406364
rect 388444 404936 388500 407036
rect 390572 407092 390628 407102
rect 377916 404450 377972 404460
rect 364700 404338 364756 404348
rect 390572 404404 390628 407036
rect 392252 406420 392308 410172
rect 460348 410228 460404 410238
rect 460348 410162 460404 410172
rect 393372 410116 393428 410126
rect 393372 410050 393428 410060
rect 398524 409780 398580 410088
rect 403704 410060 404068 410116
rect 398524 409714 398580 409724
rect 403228 409668 403284 409678
rect 403004 408548 403060 408558
rect 392252 406354 392308 406364
rect 398188 408436 398244 408446
rect 398188 405076 398244 408380
rect 398188 405010 398244 405020
rect 398412 408324 398468 408334
rect 390572 404338 390628 404348
rect 395836 404404 395892 404414
rect 395836 404338 395892 404348
rect 398412 404404 398468 408268
rect 403004 407540 403060 408492
rect 403004 407474 403060 407484
rect 403228 404936 403284 409612
rect 403900 408436 403956 408446
rect 403900 406308 403956 408380
rect 403900 406242 403956 406252
rect 403900 404964 403956 404974
rect 403900 404516 403956 404908
rect 403900 404450 403956 404460
rect 398412 404338 398468 404348
rect 404012 404404 404068 410060
rect 408828 409220 408884 410088
rect 408828 409154 408884 409164
rect 413980 408212 414036 410088
rect 419132 409332 419188 410088
rect 424312 410060 425012 410116
rect 419132 409266 419188 409276
rect 424956 409332 425012 410060
rect 424956 409266 425012 409276
rect 420028 409220 420084 409230
rect 413980 408146 414036 408156
rect 418012 408660 418068 408670
rect 410620 406980 410676 406990
rect 410620 404936 410676 406924
rect 418012 404936 418068 408604
rect 420028 408212 420084 409164
rect 420028 408146 420084 408156
rect 425404 408772 425460 408782
rect 425404 404936 425460 408716
rect 429436 404740 429492 410088
rect 432796 407092 432852 407102
rect 432796 404936 432852 407036
rect 434588 406644 434644 410088
rect 434588 406578 434644 406588
rect 439068 410060 439768 410116
rect 429436 404674 429492 404684
rect 439068 404740 439124 410060
rect 440188 406420 440244 406430
rect 440188 404936 440244 406364
rect 439068 404674 439124 404684
rect 444892 404628 444948 410088
rect 450044 409892 450100 410088
rect 450044 409826 450100 409836
rect 455196 405636 455252 410088
rect 455196 405570 455252 405580
rect 462364 404936 462420 410284
rect 465500 408100 465556 410088
rect 470652 408212 470708 410088
rect 470652 408146 470708 408156
rect 465500 408034 465556 408044
rect 469756 407428 469812 407438
rect 469756 404936 469812 407372
rect 475804 406196 475860 410088
rect 475804 406130 475860 406140
rect 477148 408548 477204 408558
rect 477148 404936 477204 408492
rect 478828 408212 478884 410396
rect 478828 408146 478884 408156
rect 484540 408436 484596 408446
rect 484540 404936 484596 408380
rect 486108 406084 486164 410088
rect 486108 406018 486164 406028
rect 491260 405748 491316 410088
rect 496412 409332 496468 410088
rect 496412 409266 496468 409276
rect 491260 405682 491316 405692
rect 491932 408324 491988 408334
rect 491932 404936 491988 408268
rect 499324 406644 499380 406654
rect 499324 404936 499380 406588
rect 501564 406644 501620 410088
rect 501564 406578 501620 406588
rect 506156 410060 506744 410116
rect 506156 405972 506212 410060
rect 506156 405906 506212 405916
rect 506716 406868 506772 406878
rect 506716 404936 506772 406812
rect 511868 406644 511924 410088
rect 511868 406578 511924 406588
rect 514108 406644 514164 406654
rect 514108 404936 514164 406588
rect 517020 406644 517076 410088
rect 517020 406578 517076 406588
rect 521500 407204 521556 407214
rect 521500 404936 521556 407148
rect 522172 406644 522228 410088
rect 522172 406578 522228 406588
rect 527324 405860 527380 410088
rect 591164 409108 591220 409118
rect 573244 406756 573300 406766
rect 527324 405794 527380 405804
rect 528892 406644 528948 406654
rect 528892 404936 528948 406588
rect 543676 406644 543732 406654
rect 543676 404936 543732 406588
rect 551068 406644 551124 406654
rect 551068 404936 551124 406588
rect 558236 406644 558292 406654
rect 558236 404964 558292 406588
rect 558236 404908 558488 404964
rect 573244 404936 573300 406700
rect 580636 406644 580692 406654
rect 580636 404936 580692 406588
rect 444892 404562 444948 404572
rect 590716 404516 590772 404526
rect 404012 404338 404068 404348
rect 536284 404404 536340 404414
rect 536284 404338 536340 404348
rect 351484 404292 351540 404302
rect 351484 404226 351540 404236
rect 373660 404292 373716 404302
rect 373660 404226 373716 404236
rect 447580 404292 447636 404302
rect 447580 404226 447636 404236
rect 454972 404292 455028 404302
rect 454972 404226 455028 404236
rect 565852 404292 565908 404302
rect 565852 404226 565908 404236
rect 590492 404068 590548 404078
rect 340620 397394 340676 397404
rect 585452 402388 585508 402398
rect 340508 395826 340564 395836
rect 585452 394884 585508 402332
rect 585452 394818 585508 394828
rect 340396 392578 340452 392588
rect 339052 392466 339108 392476
rect 338828 382274 338884 382284
rect 337820 374052 337876 374062
rect 337596 275874 337652 275884
rect 337708 369572 337764 369582
rect 337708 275716 337764 369516
rect 337820 296548 337876 373996
rect 340284 368676 340340 368686
rect 339612 367780 339668 367790
rect 338044 364196 338100 364206
rect 337820 296482 337876 296492
rect 337932 352548 337988 352558
rect 337932 277396 337988 352492
rect 338044 289044 338100 364140
rect 339500 358820 339556 358830
rect 338044 288978 338100 288988
rect 338492 357924 338548 357934
rect 337932 277330 337988 277340
rect 337708 275650 337764 275660
rect 337820 276612 337876 276622
rect 337820 268996 337876 276556
rect 337820 268930 337876 268940
rect 337932 270116 337988 270126
rect 337708 268884 337764 268894
rect 337708 260484 337764 268828
rect 337932 267148 337988 270060
rect 337708 260418 337764 260428
rect 337820 267092 337988 267148
rect 337596 256452 337652 256462
rect 337596 246932 337652 256396
rect 337820 255332 337876 267092
rect 338380 263732 338436 263742
rect 337596 246866 337652 246876
rect 337708 255276 337876 255332
rect 337932 257236 337988 257246
rect 337708 240548 337764 255276
rect 337932 255220 337988 257180
rect 338380 257124 338436 263676
rect 338380 257058 338436 257068
rect 337708 240482 337764 240492
rect 337820 255164 337988 255220
rect 337820 240546 337876 255164
rect 337932 254996 337988 255006
rect 337932 248724 337988 254940
rect 337932 248658 337988 248668
rect 338044 250180 338100 250190
rect 337820 240494 337822 240546
rect 337874 240494 337876 240546
rect 337820 240482 337876 240494
rect 337932 245476 337988 245486
rect 337932 240324 337988 245420
rect 337708 240268 337988 240324
rect 337708 236628 337764 240268
rect 337932 240098 337988 240110
rect 337932 240046 337934 240098
rect 337986 240046 337988 240098
rect 337932 237860 337988 240046
rect 337932 237794 337988 237804
rect 337708 236562 337764 236572
rect 338044 182308 338100 250124
rect 338044 182242 338100 182252
rect 338380 178052 338436 178062
rect 337484 143938 337540 143948
rect 337596 165508 337652 165518
rect 337036 128594 337092 128604
rect 336812 127586 336868 127596
rect 337596 57204 337652 165452
rect 338380 161028 338436 177996
rect 338380 160962 338436 160972
rect 338492 157780 338548 357868
rect 338492 157714 338548 157724
rect 338604 350756 338660 350766
rect 338604 155204 338660 350700
rect 338716 345380 338772 345390
rect 338716 157892 338772 345324
rect 338716 157826 338772 157836
rect 338828 304500 338884 304510
rect 338604 155138 338660 155148
rect 338828 149380 338884 304444
rect 338940 296548 338996 296558
rect 338940 287476 338996 296492
rect 338940 287410 338996 287420
rect 338940 277620 338996 277630
rect 338940 160244 338996 277564
rect 339052 253652 339108 253662
rect 339052 247044 339108 253596
rect 339500 247156 339556 358764
rect 339612 287812 339668 367724
rect 340172 357028 340228 357038
rect 339836 355236 339892 355246
rect 339724 337316 339780 337326
rect 339724 296548 339780 337260
rect 339724 296482 339780 296492
rect 339612 287746 339668 287756
rect 339500 247090 339556 247100
rect 339724 253540 339780 253550
rect 339052 246978 339108 246988
rect 339500 246932 339556 246942
rect 338940 160178 338996 160188
rect 339052 242004 339108 242014
rect 338828 149314 338884 149324
rect 339052 137508 339108 241948
rect 339500 241220 339556 246876
rect 339500 241154 339556 241164
rect 339724 229348 339780 253484
rect 339836 239876 339892 355180
rect 339836 239810 339892 239820
rect 339948 291060 340004 291070
rect 339948 236740 340004 291004
rect 339948 236674 340004 236684
rect 339724 229282 339780 229292
rect 339164 197764 339220 197774
rect 339164 172004 339220 197708
rect 339164 171938 339220 171948
rect 339276 181412 339332 181422
rect 339276 161140 339332 181356
rect 339276 161074 339332 161084
rect 339052 137442 339108 137452
rect 340172 135828 340228 356972
rect 340284 155988 340340 368620
rect 340284 155922 340340 155932
rect 340396 353108 340452 353118
rect 340396 152740 340452 353052
rect 590492 324548 590548 404012
rect 590604 394884 590660 394894
rect 590604 364196 590660 394828
rect 590604 364130 590660 364140
rect 590716 337652 590772 404460
rect 591164 403844 591220 409052
rect 591164 403778 591220 403788
rect 590716 337586 590772 337596
rect 590492 324482 590548 324492
rect 585452 284676 585508 284686
rect 340620 197204 340676 197214
rect 340620 196588 340676 197148
rect 340620 196532 341012 196588
rect 340396 152674 340452 152684
rect 340620 183764 340676 183774
rect 340172 135762 340228 135772
rect 337596 48692 337652 57148
rect 337596 48626 337652 48636
rect 335916 22866 335972 22876
rect 331884 21634 331940 21644
rect 340620 21364 340676 183708
rect 340620 21298 340676 21308
rect 340956 21252 341012 196532
rect 523292 160468 523348 160478
rect 491932 160356 491988 160366
rect 491932 160290 491988 160300
rect 506716 160244 506772 160254
rect 506716 160178 506772 160188
rect 344092 157892 344148 160104
rect 351148 160076 351512 160132
rect 351148 160020 351204 160076
rect 351148 159954 351204 159964
rect 358876 159572 358932 160104
rect 358876 159506 358932 159516
rect 344092 157826 344148 157836
rect 366268 156884 366324 160104
rect 373660 158564 373716 160104
rect 373660 158498 373716 158508
rect 381052 157668 381108 160104
rect 381052 157602 381108 157612
rect 366268 156818 366324 156828
rect 388444 155316 388500 160104
rect 388444 155250 388500 155260
rect 395836 152516 395892 160104
rect 403228 152628 403284 160104
rect 410620 152740 410676 160104
rect 410620 152674 410676 152684
rect 403228 152562 403284 152572
rect 395836 152450 395892 152460
rect 418012 149380 418068 160104
rect 422604 160020 422660 160030
rect 418012 149314 418068 149324
rect 420812 157556 420868 157566
rect 420812 144452 420868 157500
rect 420812 144386 420868 144396
rect 422380 145236 422436 145246
rect 422380 143892 422436 145180
rect 422268 143332 422324 143342
rect 421708 131012 421764 131022
rect 386204 128548 386260 128558
rect 379820 113540 379876 113550
rect 373548 106932 373604 106942
rect 373548 99988 373604 106876
rect 375116 106820 375172 106830
rect 375116 99988 375172 106764
rect 378028 104132 378084 104142
rect 376572 103236 376628 103246
rect 376572 99988 376628 103180
rect 378028 99988 378084 104076
rect 379820 99988 379876 113484
rect 384524 108724 384580 108734
rect 381388 104020 381444 104030
rect 381388 99988 381444 103964
rect 383180 103908 383236 103918
rect 383180 99988 383236 103852
rect 373548 99932 373688 99988
rect 375116 99932 375256 99988
rect 376572 99932 376824 99988
rect 378028 99932 378392 99988
rect 379820 99932 379960 99988
rect 381388 99932 381528 99988
rect 383096 99932 383236 99988
rect 384524 99988 384580 108668
rect 386204 102508 386260 128492
rect 387772 125188 387828 125198
rect 387772 102508 387828 125132
rect 411180 113428 411236 113438
rect 395500 110628 395556 110638
rect 386092 102452 386260 102508
rect 387660 102452 387828 102508
rect 388668 103796 388724 103806
rect 386092 99988 386148 102452
rect 387660 99988 387716 102452
rect 388668 99988 388724 103740
rect 390236 103684 390292 103694
rect 390236 99988 390292 103628
rect 393372 103572 393428 103582
rect 391804 103460 391860 103470
rect 391804 99988 391860 103404
rect 393372 99988 393428 103516
rect 395500 99988 395556 110572
rect 398636 110516 398692 110526
rect 396508 103348 396564 103358
rect 396508 99988 396564 103292
rect 398636 99988 398692 110460
rect 401772 110292 401828 110302
rect 400204 108388 400260 108398
rect 400204 99988 400260 108332
rect 401772 99988 401828 110236
rect 409612 110068 409668 110078
rect 404908 108500 404964 108510
rect 403228 103908 403284 103918
rect 403228 99988 403284 103852
rect 404908 99988 404964 108444
rect 407484 105364 407540 105374
rect 406700 104020 406756 104030
rect 406700 99988 406756 103964
rect 384524 99932 384664 99988
rect 386092 99932 386232 99988
rect 387660 99932 387800 99988
rect 388668 99932 389368 99988
rect 390236 99932 390936 99988
rect 391804 99932 392504 99988
rect 393372 99932 394072 99988
rect 395500 99932 395640 99988
rect 396508 99932 397208 99988
rect 398636 99932 398776 99988
rect 400204 99932 400344 99988
rect 401772 99932 401912 99988
rect 403228 99932 403480 99988
rect 404908 99932 405048 99988
rect 406616 99932 406756 99988
rect 407484 99988 407540 105308
rect 409612 99988 409668 110012
rect 411180 99988 411236 113372
rect 412188 105028 412244 105038
rect 412188 99988 412244 104972
rect 414092 104132 414148 104142
rect 414092 99988 414148 104076
rect 415660 104132 415716 104142
rect 415660 99988 415716 104076
rect 407484 99932 408184 99988
rect 409612 99932 409752 99988
rect 411180 99932 411320 99988
rect 412188 99932 412888 99988
rect 414092 99932 414456 99988
rect 415660 99932 416024 99988
rect 367052 84868 367108 84878
rect 367052 75012 367108 84812
rect 420140 77364 420196 77374
rect 367052 74946 367108 74956
rect 420028 77308 420140 77364
rect 367836 58324 367892 58334
rect 367836 57204 367892 58268
rect 367836 24612 367892 57148
rect 419244 52164 419300 52174
rect 419244 51716 419300 52108
rect 420028 52052 420084 77308
rect 420140 77298 420196 77308
rect 420028 51986 420084 51996
rect 420140 72436 420196 72446
rect 419244 51650 419300 51660
rect 420140 50372 420196 72380
rect 420252 62580 420308 62590
rect 420252 51940 420308 62524
rect 420252 51874 420308 51884
rect 421708 57652 421764 130956
rect 422268 131012 422324 143276
rect 422380 137788 422436 143836
rect 422604 143780 422660 159964
rect 422828 160020 422884 160030
rect 422604 143714 422660 143724
rect 422716 147812 422772 147822
rect 422716 144116 422772 147756
rect 422380 137732 422548 137788
rect 422380 136948 422436 136958
rect 422380 135716 422436 136892
rect 422380 135650 422436 135660
rect 422268 130946 422324 130956
rect 421820 122612 421876 122622
rect 421820 87220 421876 122556
rect 421820 87154 421876 87164
rect 421708 51828 421764 57596
rect 421708 51762 421764 51772
rect 421820 68852 421876 68862
rect 421820 67508 421876 68796
rect 420140 50306 420196 50316
rect 421820 50260 421876 67452
rect 422492 52724 422548 137732
rect 422604 135716 422660 135726
rect 422604 77364 422660 135660
rect 422604 77298 422660 77308
rect 422716 62580 422772 144060
rect 422828 143556 422884 159964
rect 425404 154420 425460 160104
rect 425404 154354 425460 154364
rect 432796 151172 432852 160104
rect 432796 151106 432852 151116
rect 423276 144116 423332 144126
rect 422828 137788 422884 143500
rect 423164 143780 423220 143790
rect 423276 143780 423332 144060
rect 423388 143780 423444 143790
rect 423276 143724 423388 143780
rect 423164 143220 423220 143724
rect 423388 143714 423444 143724
rect 422828 137732 422996 137788
rect 422940 68852 422996 137732
rect 423164 72436 423220 143164
rect 425852 141540 425908 141550
rect 425068 117572 425124 117582
rect 425068 116788 425124 117516
rect 425852 117572 425908 141484
rect 440188 135828 440244 160104
rect 447580 157780 447636 160104
rect 447580 157714 447636 157724
rect 454972 157556 455028 160104
rect 454972 157490 455028 157500
rect 457772 157556 457828 157566
rect 457772 135940 457828 157500
rect 457996 156324 458052 156334
rect 457772 135874 457828 135884
rect 457884 152628 457940 152638
rect 440188 135762 440244 135772
rect 457884 134148 457940 152572
rect 457996 137620 458052 156268
rect 462364 156324 462420 160104
rect 462364 156258 462420 156268
rect 467852 160020 467908 160030
rect 457996 137554 458052 137564
rect 458220 153076 458276 153086
rect 458220 137508 458276 153020
rect 466508 152516 466564 152526
rect 465388 148036 465444 148046
rect 458444 144564 458500 144574
rect 458220 137442 458276 137452
rect 458332 142884 458388 142894
rect 458332 135716 458388 142828
rect 458444 137732 458500 144508
rect 465388 140980 465444 147980
rect 465388 140914 465444 140924
rect 466508 143892 466564 152460
rect 466508 139944 466564 143836
rect 467852 143332 467908 159964
rect 469532 155316 469588 155326
rect 469532 143780 469588 155260
rect 469756 149492 469812 160104
rect 477148 157556 477204 160104
rect 477148 157490 477204 157500
rect 484540 155876 484596 160104
rect 499324 156996 499380 160104
rect 514108 157556 514164 160104
rect 521500 159012 521556 160104
rect 521500 158946 521556 158956
rect 514108 157490 514164 157500
rect 499324 156930 499380 156940
rect 484540 155810 484596 155820
rect 514892 155764 514948 155774
rect 469756 149426 469812 149436
rect 479052 152964 479108 152974
rect 469588 143724 469700 143780
rect 469532 143714 469588 143724
rect 467852 139972 467908 143276
rect 468524 141764 468580 141774
rect 468524 141316 468580 141708
rect 468524 141250 468580 141260
rect 467852 139916 468104 139972
rect 469644 139944 469700 143724
rect 471212 143556 471268 143566
rect 471212 139944 471268 143500
rect 472108 143220 472164 143230
rect 472108 139972 472164 143164
rect 474348 142884 474404 142894
rect 472108 139916 472808 139972
rect 474348 139944 474404 142828
rect 475916 141652 475972 141662
rect 475916 139944 475972 141596
rect 479052 139944 479108 152908
rect 510636 152404 510692 152414
rect 486892 151284 486948 151294
rect 483756 149604 483812 149614
rect 483756 139944 483812 149548
rect 485324 141204 485380 141214
rect 485324 139944 485380 141148
rect 486892 139944 486948 151228
rect 499436 149716 499492 149726
rect 494732 147924 494788 147934
rect 488460 146356 488516 146366
rect 488460 139944 488516 146300
rect 493164 146244 493220 146254
rect 490028 142884 490084 142894
rect 490028 139944 490084 142828
rect 491596 141428 491652 141438
rect 491596 139944 491652 141372
rect 493164 139944 493220 146188
rect 494732 139944 494788 147868
rect 497868 142884 497924 142894
rect 497868 139944 497924 142828
rect 499436 139944 499492 149660
rect 505596 146132 505652 146142
rect 504140 144004 504196 144014
rect 501676 142996 501732 143006
rect 480620 139748 480676 139758
rect 480620 139682 480676 139692
rect 477484 139636 477540 139646
rect 477484 139570 477540 139580
rect 482188 139636 482244 139646
rect 482188 139570 482244 139580
rect 501004 139524 501060 139534
rect 501004 139458 501060 139468
rect 501676 139524 501732 142940
rect 502572 141316 502628 141326
rect 502572 139944 502628 141260
rect 504140 139944 504196 143948
rect 505596 144004 505652 146076
rect 505596 143938 505652 143948
rect 510636 143668 510692 152348
rect 512428 149044 512484 149054
rect 512428 144116 512484 148988
rect 512428 144050 512484 144060
rect 514892 143892 514948 155708
rect 516908 154084 516964 154094
rect 514892 143826 514948 143836
rect 516684 144004 516740 144014
rect 510636 143602 510692 143612
rect 515116 143780 515172 143790
rect 507500 143556 507556 143566
rect 505708 142884 505764 142894
rect 505708 139944 505764 142828
rect 507276 142884 507332 142894
rect 507276 139944 507332 142828
rect 507500 141092 507556 143500
rect 510412 143444 510468 143454
rect 507500 141026 507556 141036
rect 508844 142884 508900 142894
rect 508844 139944 508900 142828
rect 510412 139944 510468 143388
rect 510748 143332 510804 143342
rect 510748 142772 510804 143276
rect 510748 142706 510804 142716
rect 511980 142884 512036 142894
rect 511980 139944 512036 142828
rect 513548 142884 513604 142894
rect 513548 139944 513604 142828
rect 515116 139944 515172 143724
rect 516684 139944 516740 143948
rect 516908 144004 516964 154028
rect 516908 143938 516964 143948
rect 519820 145124 519876 145134
rect 518252 142212 518308 142222
rect 518252 139944 518308 142156
rect 519820 139944 519876 145068
rect 521388 144564 521444 144574
rect 521388 139944 521444 144508
rect 522956 144116 523012 144126
rect 522956 139944 523012 144060
rect 523292 144004 523348 160412
rect 543676 160132 543732 160142
rect 528892 159124 528948 160104
rect 528892 159058 528948 159068
rect 536284 155988 536340 160104
rect 543676 160066 543732 160076
rect 551068 156100 551124 160104
rect 558460 157668 558516 160104
rect 558460 157602 558516 157612
rect 551068 156034 551124 156044
rect 536284 155922 536340 155932
rect 548044 155540 548100 155550
rect 535052 153972 535108 153982
rect 527660 150724 527716 150734
rect 523292 143938 523348 143948
rect 524524 148932 524580 148942
rect 524524 139944 524580 148876
rect 526092 147588 526148 147598
rect 526092 139944 526148 147532
rect 527660 139944 527716 150668
rect 532364 150612 532420 150622
rect 530796 150500 530852 150510
rect 529228 150388 529284 150398
rect 529228 139944 529284 150332
rect 530796 139944 530852 150444
rect 532364 139944 532420 150556
rect 533932 143892 533988 143902
rect 533932 139944 533988 143836
rect 535052 143892 535108 153916
rect 538636 145796 538692 145806
rect 535052 143826 535108 143836
rect 537068 144004 537124 144014
rect 535500 143332 535556 143342
rect 535500 139944 535556 143276
rect 537068 139944 537124 143948
rect 538636 139944 538692 145740
rect 540204 145684 540260 145694
rect 540204 139944 540260 145628
rect 541772 145572 541828 145582
rect 541772 139944 541828 145516
rect 543340 145460 543396 145470
rect 543340 139944 543396 145404
rect 544908 143780 544964 143790
rect 544908 139944 544964 143724
rect 546476 143668 546532 143678
rect 546476 139944 546532 143612
rect 548044 139944 548100 155484
rect 565852 152628 565908 160104
rect 573244 156212 573300 160104
rect 575372 158900 575428 158910
rect 574812 157444 574868 157454
rect 573244 156146 573300 156156
rect 574588 157332 574644 157342
rect 565852 152562 565908 152572
rect 562156 152292 562212 152302
rect 552748 147476 552804 147486
rect 551180 147140 551236 147150
rect 549612 141988 549668 141998
rect 549612 139944 549668 141932
rect 551180 139944 551236 147084
rect 552748 139944 552804 147420
rect 559020 147364 559076 147374
rect 555884 147252 555940 147262
rect 554316 142996 554372 143006
rect 554316 139944 554372 142940
rect 555884 139944 555940 147196
rect 557452 147028 557508 147038
rect 557452 139944 557508 146972
rect 559020 139944 559076 147308
rect 560588 143892 560644 143902
rect 560588 139944 560644 143836
rect 562156 139944 562212 152236
rect 565292 151060 565348 151070
rect 563724 143556 563780 143566
rect 563724 139944 563780 143500
rect 565292 139944 565348 151004
rect 568428 148708 568484 148718
rect 566860 145348 566916 145358
rect 566860 139944 566916 145292
rect 568428 139944 568484 148652
rect 501676 139458 501732 139468
rect 496300 139300 496356 139310
rect 496300 139234 496356 139244
rect 458444 137666 458500 137676
rect 458332 135650 458388 135660
rect 457884 134082 457940 134092
rect 574588 134036 574644 157276
rect 574588 133970 574644 133980
rect 574700 153860 574756 153870
rect 425852 117506 425908 117516
rect 425068 82292 425124 116732
rect 574700 107492 574756 153804
rect 574812 130004 574868 157388
rect 574812 129938 574868 129948
rect 574924 152068 574980 152078
rect 574924 111860 574980 152012
rect 575148 148820 575204 148830
rect 574924 111794 574980 111804
rect 575036 131908 575092 131918
rect 574700 107426 574756 107436
rect 575036 101780 575092 131852
rect 575148 117348 575204 148764
rect 575260 147700 575316 147710
rect 575260 119364 575316 147644
rect 575260 119298 575316 119308
rect 575148 117282 575204 117292
rect 575036 101714 575092 101724
rect 575372 99204 575428 158844
rect 578172 158788 578228 158798
rect 576492 157220 576548 157230
rect 576268 157108 576324 157118
rect 575596 140756 575652 140766
rect 575372 99138 575428 99148
rect 575484 138740 575540 138750
rect 458556 99092 458612 99102
rect 457772 98868 457828 98878
rect 457436 98756 457492 98766
rect 457436 91812 457492 98700
rect 457660 98420 457716 98430
rect 457660 95172 457716 98364
rect 457660 95106 457716 95116
rect 457436 91746 457492 91756
rect 425068 82226 425124 82236
rect 423164 72370 423220 72380
rect 457772 71652 457828 98812
rect 458444 97636 458500 97646
rect 458444 81732 458500 97580
rect 458444 81666 458500 81676
rect 458556 78372 458612 99036
rect 575484 93156 575540 138684
rect 575596 131908 575652 140700
rect 575596 131842 575652 131852
rect 576268 131460 576324 157052
rect 576268 131394 576324 131404
rect 576380 138964 576436 138974
rect 576380 123396 576436 138908
rect 576492 127428 576548 157164
rect 576492 127362 576548 127372
rect 576604 150948 576660 150958
rect 576380 123330 576436 123340
rect 576604 121380 576660 150892
rect 576828 140868 576884 140878
rect 576604 121314 576660 121324
rect 576716 140532 576772 140542
rect 576716 115332 576772 140476
rect 576716 115266 576772 115276
rect 576828 103236 576884 140812
rect 577948 140644 578004 140654
rect 576828 103170 576884 103180
rect 576940 140420 576996 140430
rect 576940 95172 576996 140364
rect 577948 135492 578004 140588
rect 577948 135426 578004 135436
rect 578060 138852 578116 138862
rect 576940 95106 576996 95116
rect 575484 93090 575540 93100
rect 458556 78306 458612 78316
rect 457772 71586 457828 71596
rect 578060 68964 578116 138796
rect 578172 105252 578228 158732
rect 580636 152852 580692 160104
rect 585452 155316 585508 284620
rect 587132 245028 587188 245038
rect 585452 155250 585508 155260
rect 585564 205380 585620 205390
rect 580636 152786 580692 152796
rect 585564 152516 585620 205324
rect 587132 160916 587188 244972
rect 587132 160850 587188 160860
rect 590380 178948 590436 178958
rect 590380 159236 590436 178892
rect 591276 159684 591332 430108
rect 591276 159618 591332 159628
rect 590380 159170 590436 159180
rect 585564 152450 585620 152460
rect 578396 148036 578452 148046
rect 578284 142100 578340 142110
rect 578284 109284 578340 142044
rect 578284 109218 578340 109228
rect 578172 105186 578228 105196
rect 578060 68898 578116 68908
rect 422940 68786 422996 68796
rect 578396 62916 578452 147980
rect 579628 146020 579684 146030
rect 579628 125412 579684 145964
rect 579628 125346 579684 125356
rect 581308 140308 581364 140318
rect 581308 97188 581364 140252
rect 581308 97122 581364 97132
rect 578396 62850 578452 62860
rect 422716 62514 422772 62524
rect 422492 52658 422548 52668
rect 421820 50194 421876 50204
rect 578620 48804 578676 48814
rect 578508 46788 578564 46798
rect 578172 42756 578228 42766
rect 367836 24546 367892 24556
rect 577948 30660 578004 30670
rect 574588 24052 574644 24062
rect 574588 21364 574644 23996
rect 574588 21298 574644 21308
rect 340956 21186 341012 21196
rect 577948 21252 578004 30604
rect 577948 21186 578004 21196
rect 578172 20132 578228 42700
rect 578284 38724 578340 38734
rect 578284 23044 578340 38668
rect 578284 22978 578340 22988
rect 578396 34692 578452 34702
rect 578396 21476 578452 34636
rect 578508 21812 578564 46732
rect 578508 21746 578564 21756
rect 578620 21700 578676 48748
rect 578620 21634 578676 21644
rect 578396 21410 578452 21420
rect 578172 20066 578228 20076
rect 582540 7700 582596 7710
rect 273980 4274 274036 4284
rect 580636 7588 580692 7598
rect 270508 4162 270564 4172
rect 580636 480 580692 7532
rect 582540 480 582596 7644
rect 584444 5908 584500 5918
rect 584444 480 584500 5852
rect 165564 392 165816 480
rect 167468 392 167720 480
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 392 169652 480
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 176988 392 177240 480
rect 178892 392 179144 480
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 184604 392 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 190316 392 190568 480
rect 192220 392 192472 480
rect 194124 392 194376 480
rect 196028 392 196280 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 392 198212 480
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 205548 392 205800 480
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 4956 587132 5012 587188
rect 4956 583772 5012 583828
rect 4172 390348 4228 390404
rect 4172 333340 4228 333396
rect 33292 590492 33348 590548
rect 52892 573020 52948 573076
rect 99484 590604 99540 590660
rect 77420 588812 77476 588868
rect 143388 583884 143444 583940
rect 152012 590604 152068 590660
rect 121324 582092 121380 582148
rect 94892 446012 94948 446068
rect 68572 417452 68628 417508
rect 66332 417004 66388 417060
rect 55132 414092 55188 414148
rect 64092 416892 64148 416948
rect 85260 417452 85316 417508
rect 73052 417340 73108 417396
rect 70812 417228 70868 417284
rect 75292 417116 75348 417172
rect 85036 417116 85092 417172
rect 77532 416780 77588 416836
rect 79772 416668 79828 416724
rect 62076 413420 62132 413476
rect 82236 413420 82292 413476
rect 84812 413420 84868 413476
rect 52892 390572 52948 390628
rect 59612 403676 59668 403732
rect 37996 390012 38052 390068
rect 11004 296492 11060 296548
rect 20860 388108 20916 388164
rect 4172 290780 4228 290836
rect 4172 239932 4228 239988
rect 13244 227724 13300 227780
rect 11340 47852 11396 47908
rect 15372 4172 15428 4228
rect 17276 4172 17332 4228
rect 19180 4172 19236 4228
rect 24332 384076 24388 384132
rect 34412 383964 34468 384020
rect 34412 276668 34468 276724
rect 53116 389788 53172 389844
rect 38444 384860 38500 384916
rect 37996 238476 38052 238532
rect 38220 380156 38276 380212
rect 38220 238364 38276 238420
rect 38332 379932 38388 379988
rect 40236 384748 40292 384804
rect 40124 380044 40180 380100
rect 40124 238252 40180 238308
rect 38332 238140 38388 238196
rect 44492 379596 44548 379652
rect 50652 364476 50708 364532
rect 83356 391804 83412 391860
rect 59612 383852 59668 383908
rect 69692 388220 69748 388276
rect 53116 364476 53172 364532
rect 58268 379708 58324 379764
rect 54460 362908 54516 362964
rect 65884 363804 65940 363860
rect 62076 363692 62132 363748
rect 73500 386428 73556 386484
rect 81116 379820 81172 379876
rect 77308 363916 77364 363972
rect 90076 417228 90132 417284
rect 86828 417004 86884 417060
rect 85260 397292 85316 397348
rect 86492 416668 86548 416724
rect 85036 393932 85092 393988
rect 88284 416892 88340 416948
rect 87276 409052 87332 409108
rect 87276 407484 87332 407540
rect 86828 392252 86884 392308
rect 88172 400316 88228 400372
rect 86492 385644 86548 385700
rect 86604 391580 86660 391636
rect 84812 385532 84868 385588
rect 83356 363916 83412 363972
rect 84924 379372 84980 379428
rect 88284 394044 88340 394100
rect 93324 403228 93380 403284
rect 90076 392364 90132 392420
rect 93212 397404 93268 397460
rect 89852 391580 89908 391636
rect 88172 374556 88228 374612
rect 88956 374556 89012 374612
rect 88956 373772 89012 373828
rect 86492 365372 86548 365428
rect 86492 362908 86548 362964
rect 88732 363916 88788 363972
rect 44492 319004 44548 319060
rect 86492 360332 86548 360388
rect 88956 359884 89012 359940
rect 72156 293916 72212 293972
rect 46844 292348 46900 292404
rect 59052 293132 59108 293188
rect 84588 293916 84644 293972
rect 91532 388444 91588 388500
rect 89964 360332 90020 360388
rect 89964 330876 90020 330932
rect 48300 240604 48356 240660
rect 60844 240492 60900 240548
rect 44716 240380 44772 240436
rect 53676 240268 53732 240324
rect 50092 240156 50148 240212
rect 42924 238476 42980 238532
rect 46508 238364 46564 238420
rect 51884 238252 51940 238308
rect 57260 239820 57316 239876
rect 55468 238140 55524 238196
rect 40236 237916 40292 237972
rect 59052 237916 59108 237972
rect 38220 236124 38276 236180
rect 24332 234332 24388 234388
rect 36876 236012 36932 236068
rect 35196 232764 35252 232820
rect 22764 232652 22820 232708
rect 30380 222796 30436 222852
rect 26572 219212 26628 219268
rect 24668 212492 24724 212548
rect 34412 222684 34468 222740
rect 33516 214172 33572 214228
rect 33516 4844 33572 4900
rect 32508 4284 32564 4340
rect 36092 213388 36148 213444
rect 36092 121436 36148 121492
rect 36876 49532 36932 49588
rect 37996 229404 38052 229460
rect 35196 4620 35252 4676
rect 34300 4284 34356 4340
rect 34412 4172 34468 4228
rect 41356 234556 41412 234612
rect 40012 234444 40068 234500
rect 39788 227836 39844 227892
rect 39676 222908 39732 222964
rect 38556 219436 38612 219492
rect 38444 217644 38500 217700
rect 38220 49644 38276 49700
rect 38332 214284 38388 214340
rect 38332 4956 38388 5012
rect 38444 4732 38500 4788
rect 39676 50764 39732 50820
rect 39788 50092 39844 50148
rect 39900 227612 39956 227668
rect 41244 234332 41300 234388
rect 41020 231084 41076 231140
rect 40908 219548 40964 219604
rect 40236 214396 40292 214452
rect 40012 51212 40068 51268
rect 40124 212604 40180 212660
rect 39900 49980 39956 50036
rect 40124 4508 40180 4564
rect 40908 50428 40964 50484
rect 41020 49868 41076 49924
rect 41132 230972 41188 231028
rect 41244 50652 41300 50708
rect 66220 240044 66276 240100
rect 64428 238364 64484 238420
rect 69804 237804 69860 237860
rect 68012 237692 68068 237748
rect 75180 238140 75236 238196
rect 73388 237916 73444 237972
rect 71596 237580 71652 237636
rect 77308 239372 77364 239428
rect 77308 238364 77364 238420
rect 80556 238364 80612 238420
rect 78764 238028 78820 238084
rect 85932 239708 85988 239764
rect 87724 238476 87780 238532
rect 84140 238252 84196 238308
rect 82348 237692 82404 237748
rect 76972 237580 77028 237636
rect 93212 367052 93268 367108
rect 92428 359884 92484 359940
rect 92428 250572 92484 250628
rect 92540 330876 92596 330932
rect 94892 397404 94948 397460
rect 160412 590492 160468 590548
rect 153692 583772 153748 583828
rect 155372 582092 155428 582148
rect 155372 407372 155428 407428
rect 153692 407036 153748 407092
rect 152012 395724 152068 395780
rect 186172 590940 186228 590996
rect 165676 590492 165732 590548
rect 177212 590492 177268 590548
rect 165452 588812 165508 588868
rect 163660 407484 163716 407540
rect 163100 406588 163156 406644
rect 160412 394268 160468 394324
rect 162988 405020 163044 405076
rect 99932 390124 99988 390180
rect 95116 388668 95172 388724
rect 93324 320796 93380 320852
rect 94892 388556 94948 388612
rect 93436 284732 93492 284788
rect 93436 263340 93492 263396
rect 93324 254828 93380 254884
rect 93212 246316 93268 246372
rect 93324 250572 93380 250628
rect 92540 241948 92596 242004
rect 93212 241948 93268 242004
rect 91532 237580 91588 237636
rect 62636 233324 62692 233380
rect 41356 50540 41412 50596
rect 41468 219324 41524 219380
rect 41132 49756 41188 49812
rect 40236 4284 40292 4340
rect 38556 4172 38612 4228
rect 39900 4172 39956 4228
rect 93324 224252 93380 224308
rect 93436 246316 93492 246372
rect 96572 386988 96628 387044
rect 95116 238364 95172 238420
rect 95340 386652 95396 386708
rect 94892 238252 94948 238308
rect 95340 238140 95396 238196
rect 96796 380268 96852 380324
rect 99932 238476 99988 238532
rect 103292 385084 103348 385140
rect 96796 238028 96852 238084
rect 96572 237804 96628 237860
rect 113484 383516 113540 383572
rect 111692 382060 111748 382116
rect 104972 381500 105028 381556
rect 106652 321692 106708 321748
rect 106652 267596 106708 267652
rect 104972 239820 105028 239876
rect 113372 381612 113428 381668
rect 160412 381948 160468 382004
rect 118412 381836 118468 381892
rect 113484 361340 113540 361396
rect 116732 381724 116788 381780
rect 113372 240380 113428 240436
rect 147756 320012 147812 320068
rect 139244 288988 139300 289044
rect 156268 294812 156324 294868
rect 118412 240604 118468 240660
rect 116732 240268 116788 240324
rect 162092 380380 162148 380436
rect 161308 346220 161364 346276
rect 160412 240156 160468 240212
rect 160524 318220 160580 318276
rect 111692 239708 111748 239764
rect 103292 237692 103348 237748
rect 93436 222572 93492 222628
rect 93212 217532 93268 217588
rect 154924 216748 154980 216804
rect 161308 284732 161364 284788
rect 163660 406588 163716 406644
rect 163660 406140 163716 406196
rect 163660 405020 163716 405076
rect 163100 346220 163156 346276
rect 163772 386764 163828 386820
rect 162988 342860 163044 342916
rect 163100 340956 163156 341012
rect 163100 339388 163156 339444
rect 163100 320796 163156 320852
rect 163772 340956 163828 341012
rect 170492 583884 170548 583940
rect 168812 404124 168868 404180
rect 167132 397516 167188 397572
rect 165564 395836 165620 395892
rect 166348 366156 166404 366212
rect 167132 366156 167188 366212
rect 168028 367052 168084 367108
rect 166348 365372 166404 365428
rect 165564 323372 165620 323428
rect 165676 357420 165732 357476
rect 166236 355180 166292 355236
rect 166124 328300 166180 328356
rect 165676 294812 165732 294868
rect 166012 324940 166068 324996
rect 165452 275660 165508 275716
rect 163212 259084 163268 259140
rect 162092 237916 162148 237972
rect 166124 231308 166180 231364
rect 166012 229740 166068 229796
rect 167804 354060 167860 354116
rect 166348 329420 166404 329476
rect 167692 345100 167748 345156
rect 167580 327180 167636 327236
rect 167580 233100 167636 233156
rect 166236 224476 166292 224532
rect 167804 227948 167860 228004
rect 167916 347340 167972 347396
rect 167692 223020 167748 223076
rect 168812 367052 168868 367108
rect 169596 346220 169652 346276
rect 168028 332780 168084 332836
rect 169372 342860 169428 342916
rect 169260 323820 169316 323876
rect 168812 296492 168868 296548
rect 168812 276780 168868 276836
rect 169260 234780 169316 234836
rect 167916 220892 167972 220948
rect 169372 217756 169428 217812
rect 169484 341740 169540 341796
rect 160524 216748 160580 216804
rect 169484 215964 169540 216020
rect 172956 578732 173012 578788
rect 172844 577052 172900 577108
rect 172172 407596 172228 407652
rect 171388 374556 171444 374612
rect 172172 374556 172228 374612
rect 171388 373772 171444 373828
rect 171276 352940 171332 352996
rect 171164 343980 171220 344036
rect 170940 339500 170996 339556
rect 170492 274540 170548 274596
rect 170828 330540 170884 330596
rect 170940 228060 170996 228116
rect 171052 337260 171108 337316
rect 170828 226156 170884 226212
rect 172732 348460 172788 348516
rect 171388 336140 171444 336196
rect 172396 340620 172452 340676
rect 172284 335020 172340 335076
rect 172620 333900 172676 333956
rect 172396 234668 172452 234724
rect 172508 329420 172564 329476
rect 172284 232988 172340 233044
rect 171276 231196 171332 231252
rect 171164 224588 171220 224644
rect 180012 588812 180068 588868
rect 179676 583772 179732 583828
rect 177212 397180 177268 397236
rect 179564 570444 179620 570500
rect 178892 387100 178948 387156
rect 177212 386876 177268 386932
rect 176988 383404 177044 383460
rect 177212 363916 177268 363972
rect 177436 383292 177492 383348
rect 177884 368620 177940 368676
rect 177772 367500 177828 367556
rect 177436 363804 177492 363860
rect 177660 365260 177716 365316
rect 176988 363692 177044 363748
rect 177212 356300 177268 356356
rect 176316 350700 176372 350756
rect 176204 338380 176260 338436
rect 174524 336140 174580 336196
rect 174412 326060 174468 326116
rect 172956 268940 173012 268996
rect 174300 322700 174356 322756
rect 172844 267820 172900 267876
rect 172732 232876 172788 232932
rect 172620 224812 172676 224868
rect 172508 223244 172564 223300
rect 171052 223132 171108 223188
rect 174524 229628 174580 229684
rect 174636 332780 174692 332836
rect 174412 221116 174468 221172
rect 174300 219772 174356 219828
rect 176092 321580 176148 321636
rect 176204 231420 176260 231476
rect 176092 228284 176148 228340
rect 177212 320012 177268 320068
rect 176316 219660 176372 219716
rect 177548 251020 177604 251076
rect 174636 217980 174692 218036
rect 169596 215852 169652 215908
rect 177660 239484 177716 239540
rect 177884 216076 177940 216132
rect 177996 366380 178052 366436
rect 177772 214508 177828 214564
rect 177548 213276 177604 213332
rect 178892 240044 178948 240100
rect 179116 383628 179172 383684
rect 179452 349580 179508 349636
rect 179116 239372 179172 239428
rect 179340 331660 179396 331716
rect 179340 228172 179396 228228
rect 179676 273420 179732 273476
rect 179564 272300 179620 272356
rect 184716 572908 184772 572964
rect 183036 536396 183092 536452
rect 182252 417340 182308 417396
rect 180572 416780 180628 416836
rect 182364 414092 182420 414148
rect 182364 408044 182420 408100
rect 184604 529228 184660 529284
rect 184492 514892 184548 514948
rect 183036 390796 183092 390852
rect 183932 411964 183988 412020
rect 182252 388892 182308 388948
rect 186396 590716 186452 590772
rect 186172 404460 186228 404516
rect 186284 590492 186340 590548
rect 184716 402780 184772 402836
rect 184604 395948 184660 396004
rect 186284 394604 186340 394660
rect 187740 590156 187796 590212
rect 189532 591276 189588 591332
rect 189308 576492 189364 576548
rect 188972 575036 189028 575092
rect 187964 573020 188020 573076
rect 187740 567308 187796 567364
rect 187628 557900 187684 557956
rect 187740 402444 187796 402500
rect 187852 565068 187908 565124
rect 187964 402892 188020 402948
rect 188076 569548 188132 569604
rect 187852 400652 187908 400708
rect 187628 399084 187684 399140
rect 188860 566076 188916 566132
rect 189196 569660 189252 569716
rect 188972 409948 189028 410004
rect 189084 567084 189140 567140
rect 188860 409388 188916 409444
rect 189084 401100 189140 401156
rect 189308 402668 189364 402724
rect 189420 574924 189476 574980
rect 189196 400876 189252 400932
rect 189532 410508 189588 410564
rect 189644 591052 189700 591108
rect 189644 405692 189700 405748
rect 189756 590380 189812 590436
rect 231644 590380 231700 590436
rect 253708 590156 253764 590212
rect 209580 583772 209636 583828
rect 200620 573804 200676 573860
rect 198268 573692 198324 573748
rect 193788 570332 193844 570388
rect 297836 591276 297892 591332
rect 319900 591164 319956 591220
rect 364028 591052 364084 591108
rect 341964 590156 342020 590212
rect 430220 590940 430276 590996
rect 452284 590828 452340 590884
rect 408268 588812 408324 588868
rect 386092 587244 386148 587300
rect 496412 590716 496468 590772
rect 518476 590604 518532 590660
rect 474348 578732 474404 578788
rect 562604 590492 562660 590548
rect 584668 587132 584724 587188
rect 540540 577052 540596 577108
rect 590828 576268 590884 576324
rect 530124 574924 530180 574980
rect 529676 573020 529732 573076
rect 275772 570444 275828 570500
rect 529340 572908 529396 572964
rect 200620 570332 200676 570388
rect 252028 570332 252084 570388
rect 198268 569884 198324 569940
rect 252028 568652 252084 568708
rect 193788 567084 193844 567140
rect 194012 567308 194068 567364
rect 194012 567084 194068 567140
rect 189868 566972 189924 567028
rect 189868 566076 189924 566132
rect 529564 569772 529620 569828
rect 529340 448028 529396 448084
rect 529452 567084 529508 567140
rect 530012 569660 530068 569716
rect 529900 568316 529956 568372
rect 529788 568204 529844 568260
rect 590604 574588 590660 574644
rect 532924 573580 532980 573636
rect 532812 573132 532868 573188
rect 532700 571676 532756 571732
rect 531132 571452 531188 571508
rect 530908 569548 530964 569604
rect 530124 485100 530180 485156
rect 530236 567196 530292 567252
rect 530124 480396 530180 480452
rect 529900 476252 529956 476308
rect 529788 461916 529844 461972
rect 529676 456988 529732 457044
rect 529564 452732 529620 452788
rect 529452 443324 529508 443380
rect 530236 433356 530292 433412
rect 531020 566972 531076 567028
rect 532588 569884 532644 569940
rect 532588 536844 532644 536900
rect 533372 573468 533428 573524
rect 533260 573356 533316 573412
rect 533036 571564 533092 571620
rect 533148 569996 533204 570052
rect 533372 527436 533428 527492
rect 533484 571900 533540 571956
rect 533260 522732 533316 522788
rect 533148 518028 533204 518084
rect 533036 513324 533092 513380
rect 532924 503916 532980 503972
rect 532812 499212 532868 499268
rect 532700 470988 532756 471044
rect 531132 438060 531188 438116
rect 531020 423948 531076 424004
rect 530908 419244 530964 419300
rect 590492 567980 590548 568036
rect 590716 571340 590772 571396
rect 591164 574700 591220 574756
rect 590828 522732 590884 522788
rect 590940 571228 590996 571284
rect 591052 567868 591108 567924
rect 591164 562380 591220 562436
rect 591052 535836 591108 535892
rect 590940 483084 590996 483140
rect 590716 456652 590772 456708
rect 590604 443436 590660 443492
rect 590492 417004 590548 417060
rect 591276 430108 591332 430164
rect 533484 414540 533540 414596
rect 203756 410508 203812 410564
rect 189756 403788 189812 403844
rect 192332 409948 192388 410004
rect 189420 399420 189476 399476
rect 188076 397964 188132 398020
rect 186396 394380 186452 394436
rect 197484 407148 197540 407204
rect 200732 409724 200788 409780
rect 200732 409052 200788 409108
rect 202524 409388 202580 409444
rect 197596 404124 197652 404180
rect 199052 406700 199108 406756
rect 197484 398076 197540 398132
rect 202412 404460 202468 404516
rect 199052 397740 199108 397796
rect 200508 398076 200564 398132
rect 192444 397516 192500 397572
rect 192332 392588 192388 392644
rect 196364 395612 196420 395668
rect 184492 392476 184548 392532
rect 183932 385868 183988 385924
rect 180572 385756 180628 385812
rect 200508 389004 200564 389060
rect 201068 394604 201124 394660
rect 199724 382844 199780 382900
rect 198380 382284 198436 382340
rect 197036 382172 197092 382228
rect 198156 382172 198212 382228
rect 199052 382172 199108 382228
rect 199948 382172 200004 382228
rect 201740 394380 201796 394436
rect 202748 407596 202804 407652
rect 203084 405692 203140 405748
rect 202524 394380 202580 394436
rect 202636 397740 202692 397796
rect 202636 387212 202692 387268
rect 480508 410508 480564 410564
rect 352828 410396 352884 410452
rect 339388 410284 339444 410340
rect 206556 409724 206612 409780
rect 204988 409052 205044 409108
rect 204428 403788 204484 403844
rect 204988 398076 205044 398132
rect 206556 407932 206612 407988
rect 205212 397180 205268 397236
rect 205772 395724 205828 395780
rect 206444 394268 206500 394324
rect 206556 382172 206612 382228
rect 207116 390572 207172 390628
rect 207900 409724 207956 409780
rect 213052 406140 213108 406196
rect 213052 405804 213108 405860
rect 216636 406588 216692 406644
rect 207452 387996 207508 388052
rect 209132 397404 209188 397460
rect 208236 384188 208292 384244
rect 207788 382956 207844 383012
rect 208908 383068 208964 383124
rect 208908 380492 208964 380548
rect 212492 384076 212548 384132
rect 211820 383964 211876 384020
rect 209804 383852 209860 383908
rect 210476 383516 210532 383572
rect 214508 381388 214564 381444
rect 216524 381388 216580 381444
rect 215852 379932 215908 379988
rect 218204 406588 218260 406644
rect 233660 407260 233716 407316
rect 238028 410060 238084 410116
rect 228508 398076 228564 398132
rect 223356 396396 223412 396452
rect 223356 395724 223412 395780
rect 229404 394380 229460 394436
rect 227612 392588 227668 392644
rect 219884 390012 219940 390068
rect 217532 389004 217588 389060
rect 217532 384636 217588 384692
rect 218204 387212 218260 387268
rect 216636 380604 216692 380660
rect 217868 382620 217924 382676
rect 218204 382508 218260 382564
rect 219212 384860 219268 384916
rect 225932 384748 225988 384804
rect 225148 384636 225204 384692
rect 225148 382620 225204 382676
rect 222572 381948 222628 382004
rect 221900 381836 221956 381892
rect 220556 381612 220612 381668
rect 221228 380156 221284 380212
rect 223916 381724 223972 381780
rect 223244 380492 223300 380548
rect 225260 381500 225316 381556
rect 224140 380044 224196 380100
rect 227612 383964 227668 384020
rect 228620 387100 228676 387156
rect 227276 383740 227332 383796
rect 226604 383180 226660 383236
rect 227948 383628 228004 383684
rect 229292 384972 229348 385028
rect 229628 392476 229684 392532
rect 237356 391580 237412 391636
rect 229852 390684 229908 390740
rect 236684 390124 236740 390180
rect 233996 388668 234052 388724
rect 232652 388444 232708 388500
rect 229852 382956 229908 383012
rect 229964 386988 230020 387044
rect 229628 382844 229684 382900
rect 229404 382732 229460 382788
rect 231980 386652 232036 386708
rect 230636 386540 230692 386596
rect 231308 380380 231364 380436
rect 233324 380268 233380 380324
rect 235340 388556 235396 388612
rect 234668 385084 234724 385140
rect 236012 382060 236068 382116
rect 238812 409276 238868 409332
rect 238700 409164 238756 409220
rect 249116 409388 249172 409444
rect 249788 409388 249844 409444
rect 249788 407596 249844 407652
rect 253484 407484 253540 407540
rect 243964 406476 244020 406532
rect 252812 406700 252868 406756
rect 252140 404684 252196 404740
rect 242060 404460 242116 404516
rect 240716 402332 240772 402388
rect 240044 397964 240100 398020
rect 239372 382284 239428 382340
rect 241388 401100 241444 401156
rect 244076 403900 244132 403956
rect 243404 383852 243460 383908
rect 242732 381948 242788 382004
rect 250796 402892 250852 402948
rect 248108 402780 248164 402836
rect 246764 402444 246820 402500
rect 244748 399084 244804 399140
rect 245420 397852 245476 397908
rect 246092 382060 246148 382116
rect 247436 402444 247492 402500
rect 249452 400988 249508 401044
rect 248780 392476 248836 392532
rect 250124 395836 250180 395892
rect 251468 382844 251524 382900
rect 253708 407484 253764 407540
rect 259420 409500 259476 409556
rect 259420 409276 259476 409332
rect 261996 409276 262052 409332
rect 261548 407820 261604 407876
rect 254268 407484 254324 407540
rect 254828 407708 254884 407764
rect 253708 407148 253764 407204
rect 254156 382732 254212 382788
rect 255500 404684 255556 404740
rect 256172 404572 256228 404628
rect 259532 404572 259588 404628
rect 257516 400876 257572 400932
rect 256844 392588 256900 392644
rect 258860 399420 258916 399476
rect 258188 392700 258244 392756
rect 260204 402668 260260 402724
rect 260876 381612 260932 381668
rect 264572 407932 264628 407988
rect 264908 409052 264964 409108
rect 261996 407708 262052 407764
rect 264236 404796 264292 404852
rect 262892 404012 262948 404068
rect 262220 381948 262276 382004
rect 263564 382508 263620 382564
rect 273756 409948 273812 410004
rect 273756 407932 273812 407988
rect 274652 409612 274708 409668
rect 268716 404908 268772 404964
rect 271628 405692 271684 405748
rect 267596 404012 267652 404068
rect 265580 400764 265636 400820
rect 266924 395948 266980 396004
rect 266252 383964 266308 384020
rect 268716 385980 268772 386036
rect 269612 404348 269668 404404
rect 268940 382620 268996 382676
rect 268268 382396 268324 382452
rect 270956 399308 271012 399364
rect 270284 382396 270340 382452
rect 272972 405244 273028 405300
rect 272300 397740 272356 397796
rect 273644 404124 273700 404180
rect 274316 397404 274372 397460
rect 274876 409612 274932 409668
rect 277228 407372 277284 407428
rect 274652 383180 274708 383236
rect 274652 380604 274708 380660
rect 274988 404236 275044 404292
rect 276332 397628 276388 397684
rect 275660 395948 275716 396004
rect 280028 407372 280084 407428
rect 284732 408044 284788 408100
rect 284396 402668 284452 402724
rect 281708 402556 281764 402612
rect 277676 400652 277732 400708
rect 277228 394492 277284 394548
rect 277340 390796 277396 390852
rect 277340 390460 277396 390516
rect 277228 387212 277284 387268
rect 277004 382508 277060 382564
rect 280364 399196 280420 399252
rect 279020 397516 279076 397572
rect 278012 390796 278068 390852
rect 278012 380604 278068 380660
rect 278796 381948 278852 382004
rect 279692 397516 279748 397572
rect 281036 396060 281092 396116
rect 283724 402556 283780 402612
rect 283052 396172 283108 396228
rect 286412 408828 286468 408884
rect 284732 390572 284788 390628
rect 285068 404348 285124 404404
rect 285740 399196 285796 399252
rect 289772 408380 289828 408436
rect 289100 399420 289156 399476
rect 287756 396284 287812 396340
rect 287084 389004 287140 389060
rect 288428 389116 288484 389172
rect 289884 407036 289940 407092
rect 291788 409052 291844 409108
rect 291116 402892 291172 402948
rect 289884 394268 289940 394324
rect 290444 396396 290500 396452
rect 294812 407932 294868 407988
rect 293804 404124 293860 404180
rect 292460 392924 292516 392980
rect 293132 381388 293188 381444
rect 299964 407820 300020 407876
rect 299180 407148 299236 407204
rect 296492 405020 296548 405076
rect 294812 386092 294868 386148
rect 295148 392812 295204 392868
rect 294476 381612 294532 381668
rect 295820 389228 295876 389284
rect 297836 399532 297892 399588
rect 297164 381948 297220 382004
rect 298956 381948 299012 382004
rect 299852 399644 299908 399700
rect 299964 390684 300020 390740
rect 302540 408604 302596 408660
rect 301196 382060 301252 382116
rect 300524 381948 300580 382004
rect 302204 381948 302260 382004
rect 310940 409836 310996 409892
rect 305788 408044 305844 408100
rect 305788 406588 305844 406644
rect 306796 406588 306852 406644
rect 305228 389788 305284 389844
rect 303212 382060 303268 382116
rect 303884 381948 303940 382004
rect 304556 381612 304612 381668
rect 309260 391804 309316 391860
rect 306796 383964 306852 384020
rect 307916 388220 307972 388276
rect 306572 383404 306628 383460
rect 307244 383292 307300 383348
rect 308588 386428 308644 386484
rect 311276 386876 311332 386932
rect 315308 397292 315364 397348
rect 313964 394044 314020 394100
rect 311612 380716 311668 380772
rect 311948 387212 312004 387268
rect 312620 385868 312676 385924
rect 313292 381948 313348 382004
rect 314636 392252 314692 392308
rect 315980 392364 316036 392420
rect 317324 393932 317380 393988
rect 316092 388220 316148 388276
rect 316652 388892 316708 388948
rect 321692 390348 321748 390404
rect 317996 385756 318052 385812
rect 318668 385644 318724 385700
rect 319340 385532 319396 385588
rect 326396 385196 326452 385252
rect 329644 399868 329700 399924
rect 321692 380828 321748 380884
rect 309932 379820 309988 379876
rect 305900 379708 305956 379764
rect 211148 379596 211204 379652
rect 218540 379596 218596 379652
rect 190764 379484 190820 379540
rect 191324 379484 191380 379540
rect 192108 379484 192164 379540
rect 192668 379484 192724 379540
rect 193340 379484 193396 379540
rect 194684 379484 194740 379540
rect 195244 379484 195300 379540
rect 282380 379484 282436 379540
rect 310604 379372 310660 379428
rect 193004 379260 193060 379316
rect 195020 379260 195076 379316
rect 213164 379260 213220 379316
rect 213836 379260 213892 379316
rect 215180 379260 215236 379316
rect 217196 379260 217252 379316
rect 329532 366268 329588 366324
rect 329420 362908 329476 362964
rect 180012 270396 180068 270452
rect 180124 351260 180180 351316
rect 180124 229516 180180 229572
rect 180236 293020 180292 293076
rect 179452 217868 179508 217924
rect 329532 308364 329588 308420
rect 330988 398188 331044 398244
rect 330316 395724 330372 395780
rect 330092 385980 330148 386036
rect 329756 346556 329812 346612
rect 329980 308924 330036 308980
rect 329980 307916 330036 307972
rect 329644 295596 329700 295652
rect 329756 307356 329812 307412
rect 329420 259532 329476 259588
rect 329532 270508 329588 270564
rect 329420 241948 329476 242004
rect 327964 240492 328020 240548
rect 184940 240044 184996 240100
rect 184940 238476 184996 238532
rect 186396 238476 186452 238532
rect 186732 232652 186788 232708
rect 186396 229292 186452 229348
rect 185836 227724 185892 227780
rect 188524 229404 188580 229460
rect 189420 222908 189476 222964
rect 187628 222796 187684 222852
rect 191212 232764 191268 232820
rect 190316 219548 190372 219604
rect 180236 212940 180292 212996
rect 177996 212828 178052 212884
rect 196588 234556 196644 234612
rect 195692 234444 195748 234500
rect 198380 236124 198436 236180
rect 199276 236012 199332 236068
rect 200172 234444 200228 234500
rect 197484 234332 197540 234388
rect 194796 231084 194852 231140
rect 193900 227836 193956 227892
rect 202860 233436 202916 233492
rect 201964 233324 202020 233380
rect 203756 229964 203812 230020
rect 201068 225036 201124 225092
rect 208236 232540 208292 232596
rect 209132 231756 209188 231812
rect 207340 230076 207396 230132
rect 210924 228396 210980 228452
rect 210028 227836 210084 227892
rect 213612 234556 213668 234612
rect 214508 230860 214564 230916
rect 212716 229180 212772 229236
rect 211820 227724 211876 227780
rect 206444 224140 206500 224196
rect 205548 221564 205604 221620
rect 204652 217420 204708 217476
rect 193004 214396 193060 214452
rect 192108 212604 192164 212660
rect 216300 222684 216356 222740
rect 217196 219436 217252 219492
rect 218092 214284 218148 214340
rect 220780 224364 220836 224420
rect 226716 236908 226772 236964
rect 225260 235116 225316 235172
rect 224364 235004 224420 235060
rect 223468 230972 223524 231028
rect 227052 230972 227108 231028
rect 222572 227612 222628 227668
rect 228844 227612 228900 227668
rect 227948 227500 228004 227556
rect 231756 236908 231812 236964
rect 230636 234220 230692 234276
rect 236012 238028 236068 238084
rect 235116 237132 235172 237188
rect 234220 237020 234276 237076
rect 233324 236908 233380 236964
rect 232428 224364 232484 224420
rect 229740 221676 229796 221732
rect 221676 219324 221732 219380
rect 219884 217644 219940 217700
rect 218988 214172 219044 214228
rect 237804 238140 237860 238196
rect 239596 238364 239652 238420
rect 240492 237804 240548 237860
rect 238700 237692 238756 237748
rect 236908 213052 236964 213108
rect 215404 212492 215460 212548
rect 243180 238252 243236 238308
rect 242284 237916 242340 237972
rect 244972 217644 245028 217700
rect 244076 216636 244132 216692
rect 247660 222684 247716 222740
rect 248556 214284 248612 214340
rect 246764 214172 246820 214228
rect 245868 212492 245924 212548
rect 251244 238476 251300 238532
rect 252140 237580 252196 237636
rect 250348 222460 250404 222516
rect 253932 213164 253988 213220
rect 256620 215740 256676 215796
rect 255724 213276 255780 213332
rect 258412 219324 258468 219380
rect 257516 211596 257572 211652
rect 254828 211372 254884 211428
rect 253036 211260 253092 211316
rect 249452 211148 249508 211204
rect 260204 219436 260260 219492
rect 261996 219100 262052 219156
rect 261100 212380 261156 212436
rect 264460 237020 264516 237076
rect 265356 236908 265412 236964
rect 266252 236908 266308 236964
rect 268044 237020 268100 237076
rect 267036 236908 267092 236964
rect 269836 237020 269892 237076
rect 270172 239820 270228 239876
rect 268604 236908 268660 236964
rect 270284 236908 270340 236964
rect 270620 238140 270676 238196
rect 270172 235004 270228 235060
rect 268940 228396 268996 228452
rect 268828 227836 268884 227892
rect 262892 211484 262948 211540
rect 267932 211596 267988 211652
rect 267932 211372 267988 211428
rect 259308 210700 259364 210756
rect 241388 210028 241444 210084
rect 98924 50652 98980 50708
rect 87500 50540 87556 50596
rect 53228 50428 53284 50484
rect 45612 50316 45668 50372
rect 41468 4172 41524 4228
rect 41804 4956 41860 5012
rect 49420 41132 49476 41188
rect 47516 4956 47572 5012
rect 76076 50092 76132 50148
rect 74172 48076 74228 48132
rect 68460 41468 68516 41524
rect 62748 41356 62804 41412
rect 57148 41244 57204 41300
rect 55132 4844 55188 4900
rect 60844 4732 60900 4788
rect 58940 4620 58996 4676
rect 64652 4508 64708 4564
rect 66556 4396 66612 4452
rect 70364 4284 70420 4340
rect 72268 4172 72324 4228
rect 77980 49980 78036 50036
rect 81788 49868 81844 49924
rect 79884 41580 79940 41636
rect 83692 49756 83748 49812
rect 85708 41692 85764 41748
rect 89404 50540 89460 50596
rect 93212 50428 93268 50484
rect 91308 47964 91364 48020
rect 97356 48636 97412 48692
rect 97020 48188 97076 48244
rect 95116 42812 95172 42868
rect 97356 47852 97412 47908
rect 137004 50652 137060 50708
rect 104636 49644 104692 49700
rect 102732 47852 102788 47908
rect 100828 46172 100884 46228
rect 110348 49532 110404 49588
rect 108444 44492 108500 44548
rect 106540 42924 106596 42980
rect 114268 49532 114324 49588
rect 112252 43148 112308 43204
rect 125580 44828 125636 44884
rect 119868 44604 119924 44660
rect 116060 43036 116116 43092
rect 117964 39452 118020 39508
rect 123676 39564 123732 39620
rect 121772 32732 121828 32788
rect 131292 44716 131348 44772
rect 129388 36092 129444 36148
rect 127484 32844 127540 32900
rect 135100 39676 135156 39732
rect 133196 32956 133252 33012
rect 173180 50540 173236 50596
rect 167468 49868 167524 49924
rect 152236 49756 152292 49812
rect 150332 46284 150388 46340
rect 148428 44940 148484 44996
rect 144620 43260 144676 43316
rect 140812 36204 140868 36260
rect 138908 33068 138964 33124
rect 142828 29372 142884 29428
rect 146524 36316 146580 36372
rect 156044 49644 156100 49700
rect 154140 45052 154196 45108
rect 159852 48300 159908 48356
rect 158172 7532 158228 7588
rect 161756 46396 161812 46452
rect 165564 26012 165620 26068
rect 163884 9212 163940 9268
rect 171388 45164 171444 45220
rect 169596 4172 169652 4228
rect 178892 50540 178948 50596
rect 175084 41804 175140 41860
rect 176988 37772 177044 37828
rect 268828 50540 268884 50596
rect 184604 50428 184660 50484
rect 182700 26124 182756 26180
rect 180796 19292 180852 19348
rect 269836 222684 269892 222740
rect 269612 222460 269668 222516
rect 268940 50428 268996 50484
rect 269052 212940 269108 212996
rect 190316 50316 190372 50372
rect 188412 47628 188468 47684
rect 186508 34412 186564 34468
rect 196028 50316 196084 50372
rect 194124 45276 194180 45332
rect 192220 15932 192276 15988
rect 201740 50316 201796 50372
rect 199948 41916 200004 41972
rect 198156 4284 198212 4340
rect 209356 50316 209412 50372
rect 207452 48524 207508 48580
rect 205548 44380 205604 44436
rect 203644 43372 203700 43428
rect 212268 47740 212324 47796
rect 269500 209804 269556 209860
rect 269500 207564 269556 207620
rect 270508 213052 270564 213108
rect 269948 113484 270004 113540
rect 269612 108668 269668 108724
rect 269052 47740 269108 47796
rect 211260 37884 211316 37940
rect 270844 229180 270900 229236
rect 270620 41804 270676 41860
rect 270732 221676 270788 221732
rect 272076 236908 272132 236964
rect 272188 238364 272244 238420
rect 271516 234556 271572 234612
rect 271404 230860 271460 230916
rect 270956 137676 271012 137732
rect 271068 227724 271124 227780
rect 270844 51548 270900 51604
rect 271292 210588 271348 210644
rect 271516 197372 271572 197428
rect 271404 190652 271460 190708
rect 271292 108332 271348 108388
rect 271068 51436 271124 51492
rect 270732 39564 270788 39620
rect 272636 237692 272692 237748
rect 272300 232764 272356 232820
rect 272300 199164 272356 199220
rect 272524 210476 272580 210532
rect 272300 197372 272356 197428
rect 272300 51660 272356 51716
rect 272412 190652 272468 190708
rect 273644 211596 273700 211652
rect 273868 237804 273924 237860
rect 272748 211260 272804 211316
rect 273196 209804 273252 209860
rect 272636 186396 272692 186452
rect 272748 209468 272804 209524
rect 272860 209356 272916 209412
rect 273084 209132 273140 209188
rect 272972 206332 273028 206388
rect 272972 190652 273028 190708
rect 272860 166236 272916 166292
rect 272972 185948 273028 186004
rect 272748 163324 272804 163380
rect 272524 148764 272580 148820
rect 272860 121772 272916 121828
rect 272860 119644 272916 119700
rect 272860 58492 272916 58548
rect 272860 51884 272916 51940
rect 273196 174972 273252 175028
rect 273420 176316 273476 176372
rect 273084 169148 273140 169204
rect 273196 143388 273252 143444
rect 273084 139020 273140 139076
rect 273420 143388 273476 143444
rect 273196 134204 273252 134260
rect 273084 75964 273140 76020
rect 273196 91532 273252 91588
rect 273196 73052 273252 73108
rect 273308 86492 273364 86548
rect 273420 83132 273476 83188
rect 273420 78876 273476 78932
rect 273308 70140 273364 70196
rect 273084 67228 273140 67284
rect 273084 51996 273140 52052
rect 273196 64316 273252 64372
rect 273196 50316 273252 50372
rect 272972 49868 273028 49924
rect 272412 48524 272468 48580
rect 272188 34412 272244 34468
rect 274764 237580 274820 237636
rect 274092 233436 274148 233492
rect 273868 15932 273924 15988
rect 273980 208908 274036 208964
rect 274092 32956 274148 33012
rect 274204 225036 274260 225092
rect 274316 224364 274372 224420
rect 274428 221564 274484 221620
rect 274652 211372 274708 211428
rect 275212 237020 275268 237076
rect 275884 238252 275940 238308
rect 275436 236908 275492 236964
rect 275660 237916 275716 237972
rect 275548 233324 275604 233380
rect 274876 211596 274932 211652
rect 274876 147532 274932 147588
rect 274764 125132 274820 125188
rect 274652 103292 274708 103348
rect 274652 99036 274708 99092
rect 274652 81788 274708 81844
rect 274428 46284 274484 46340
rect 274316 36204 274372 36260
rect 275660 43372 275716 43428
rect 275772 234444 275828 234500
rect 277900 237020 277956 237076
rect 277004 236908 277060 236964
rect 278684 236908 278740 236964
rect 277452 232540 277508 232596
rect 275996 231644 276052 231700
rect 277228 229292 277284 229348
rect 276332 224252 276388 224308
rect 276332 204092 276388 204148
rect 276444 217644 276500 217700
rect 275996 178444 276052 178500
rect 276332 197708 276388 197764
rect 275884 51772 275940 51828
rect 275772 43036 275828 43092
rect 276780 211148 276836 211204
rect 276444 106764 276500 106820
rect 276556 210924 276612 210980
rect 276780 103852 276836 103908
rect 276556 103404 276612 103460
rect 276444 61404 276500 61460
rect 276444 50204 276500 50260
rect 277228 48636 277284 48692
rect 277340 217420 277396 217476
rect 278908 229964 278964 230020
rect 278124 219436 278180 219492
rect 277452 185948 277508 186004
rect 278012 214284 278068 214340
rect 278348 219324 278404 219380
rect 278124 110236 278180 110292
rect 278236 213164 278292 213220
rect 278012 103964 278068 104020
rect 278684 211260 278740 211316
rect 278348 110460 278404 110516
rect 278460 210700 278516 210756
rect 278684 148876 278740 148932
rect 278460 103740 278516 103796
rect 278236 103628 278292 103684
rect 277340 43260 277396 43316
rect 276332 41916 276388 41972
rect 279020 142716 279076 142772
rect 279132 224140 279188 224196
rect 279692 219100 279748 219156
rect 279692 108444 279748 108500
rect 279804 213276 279860 213332
rect 280364 237916 280420 237972
rect 279916 160300 279972 160356
rect 280028 215740 280084 215796
rect 280476 237132 280532 237188
rect 280476 147084 280532 147140
rect 280588 235900 280644 235956
rect 280364 146972 280420 147028
rect 280028 110572 280084 110628
rect 279804 103516 279860 103572
rect 280812 145740 280868 145796
rect 281372 239484 281428 239540
rect 280588 93436 280644 93492
rect 279132 49644 279188 49700
rect 278908 33068 278964 33124
rect 275548 32844 275604 32900
rect 274204 32732 274260 32788
rect 281596 233212 281652 233268
rect 281484 231532 281540 231588
rect 281484 45276 281540 45332
rect 281372 26124 281428 26180
rect 281708 145628 281764 145684
rect 281820 238476 281876 238532
rect 282044 238140 282100 238196
rect 282044 148652 282100 148708
rect 282156 237020 282212 237076
rect 282156 141932 282212 141988
rect 282268 230076 282324 230132
rect 281820 128492 281876 128548
rect 282156 93996 282212 94052
rect 282156 93436 282212 93492
rect 282268 46396 282324 46452
rect 282380 221452 282436 221508
rect 282604 145516 282660 145572
rect 283052 214172 283108 214228
rect 283388 199388 283444 199444
rect 283388 157500 283444 157556
rect 283836 236908 283892 236964
rect 283612 199612 283668 199668
rect 283612 157724 283668 157780
rect 283724 199500 283780 199556
rect 283724 157276 283780 157332
rect 284732 239708 284788 239764
rect 284620 199724 284676 199780
rect 284620 157836 284676 157892
rect 284396 152348 284452 152404
rect 283836 147420 283892 147476
rect 283500 145404 283556 145460
rect 283052 104076 283108 104132
rect 285068 234220 285124 234276
rect 284956 210924 285012 210980
rect 284956 160524 285012 160580
rect 285180 234108 285236 234164
rect 285404 155484 285460 155540
rect 285516 237356 285572 237412
rect 285292 154028 285348 154084
rect 287308 238700 287364 238756
rect 287308 237804 287364 237860
rect 287980 237132 288036 237188
rect 287084 237020 287140 237076
rect 288876 236908 288932 236964
rect 291564 237916 291620 237972
rect 292460 237692 292516 237748
rect 290668 237356 290724 237412
rect 290444 236908 290500 236964
rect 294252 238028 294308 238084
rect 293804 236908 293860 236964
rect 296044 237916 296100 237972
rect 297836 238140 297892 238196
rect 296940 237020 296996 237076
rect 295372 236908 295428 236964
rect 298956 236908 299012 236964
rect 285964 235004 286020 235060
rect 285516 147196 285572 147252
rect 285852 216636 285908 216692
rect 285852 106876 285908 106932
rect 284732 45052 284788 45108
rect 282380 44380 282436 44436
rect 290444 234780 290500 234836
rect 288204 228284 288260 228340
rect 289324 219772 289380 219828
rect 293804 233100 293860 233156
rect 291564 229740 291620 229796
rect 292684 221116 292740 221172
rect 294924 231308 294980 231364
rect 298284 228172 298340 228228
rect 297164 226156 297220 226212
rect 296044 223244 296100 223300
rect 299404 217980 299460 218036
rect 300300 200060 300356 200116
rect 300412 224812 300468 224868
rect 299628 199948 299684 200004
rect 301196 199948 301252 200004
rect 301644 232988 301700 233044
rect 301420 199948 301476 200004
rect 302764 229628 302820 229684
rect 304108 238140 304164 238196
rect 305900 238252 305956 238308
rect 305676 236908 305732 236964
rect 305004 231420 305060 231476
rect 303884 223132 303940 223188
rect 306124 228060 306180 228116
rect 307692 238364 307748 238420
rect 306796 202636 306852 202692
rect 307244 234668 307300 234724
rect 308364 215964 308420 216020
rect 303212 199388 303268 199444
rect 309372 217756 309428 217812
rect 309484 202748 309540 202804
rect 308588 199388 308644 199444
rect 310604 224588 310660 224644
rect 311724 223020 311780 223076
rect 310380 199388 310436 199444
rect 313964 234220 314020 234276
rect 313068 234108 313124 234164
rect 313964 220892 314020 220948
rect 312172 210924 312228 210980
rect 312844 215852 312900 215908
rect 315084 232876 315140 232932
rect 314860 199724 314916 199780
rect 316204 217868 316260 217924
rect 315756 199612 315812 199668
rect 317324 219660 317380 219716
rect 316652 199500 316708 199556
rect 311836 199388 311892 199444
rect 318444 238028 318500 238084
rect 318444 229516 318500 229572
rect 319564 231196 319620 231252
rect 321132 237580 321188 237636
rect 320236 199948 320292 200004
rect 320684 227948 320740 228004
rect 321804 224476 321860 224532
rect 322924 237468 322980 237524
rect 322028 199948 322084 200004
rect 325388 238364 325444 238420
rect 325164 238140 325220 238196
rect 323820 199612 323876 199668
rect 324492 238028 324548 238084
rect 319340 199500 319396 199556
rect 317548 199388 317604 199444
rect 324380 236460 324436 236516
rect 324940 237916 324996 237972
rect 324156 198268 324212 198324
rect 324268 199724 324324 199780
rect 286188 160524 286244 160580
rect 298060 160300 298116 160356
rect 307692 160188 307748 160244
rect 291564 157836 291620 157892
rect 293356 157724 293412 157780
rect 296940 157500 296996 157556
rect 295148 157276 295204 157332
rect 304108 160076 304164 160132
rect 302316 157724 302372 157780
rect 311276 159180 311332 159236
rect 309484 157836 309540 157892
rect 305900 157612 305956 157668
rect 300524 157164 300580 157220
rect 313068 156044 313124 156100
rect 316652 157500 316708 157556
rect 320236 157388 320292 157444
rect 324380 198268 324436 198324
rect 324380 195132 324436 195188
rect 324268 157724 324324 157780
rect 324492 159180 324548 159236
rect 323820 157276 323876 157332
rect 322028 157052 322084 157108
rect 324604 199836 324660 199892
rect 324716 192220 324772 192276
rect 324604 157612 324660 157668
rect 324492 156940 324548 156996
rect 318444 156716 318500 156772
rect 314860 155932 314916 155988
rect 324940 151004 324996 151060
rect 325052 212492 325108 212548
rect 324156 144060 324212 144116
rect 318556 142604 318612 142660
rect 318332 142380 318388 142436
rect 309932 142268 309988 142324
rect 308252 138796 308308 138852
rect 287756 128604 287812 128660
rect 287756 122556 287812 122612
rect 308252 107996 308308 108052
rect 309932 87612 309988 87668
rect 311612 139132 311668 139188
rect 323372 142492 323428 142548
rect 323372 105084 323428 105140
rect 323484 122668 323540 122724
rect 318556 96348 318612 96404
rect 324156 122668 324212 122724
rect 325836 237916 325892 237972
rect 326732 237804 326788 237860
rect 326060 237580 326116 237636
rect 325948 237468 326004 237524
rect 325948 160188 326004 160244
rect 326060 160076 326116 160132
rect 326284 199612 326340 199668
rect 326284 157836 326340 157892
rect 326508 199500 326564 199556
rect 326508 157164 326564 157220
rect 327516 237804 327572 237860
rect 327404 237692 327460 237748
rect 326844 236348 326900 236404
rect 327516 234892 327572 234948
rect 327852 237580 327908 237636
rect 326844 217532 326900 217588
rect 326956 222572 327012 222628
rect 326732 152236 326788 152292
rect 326844 198828 326900 198884
rect 326956 198044 327012 198100
rect 326844 148764 326900 148820
rect 327404 186396 327460 186452
rect 327404 185276 327460 185332
rect 325836 144396 325892 144452
rect 325388 142044 325444 142100
rect 325164 140588 325220 140644
rect 325052 103180 325108 103236
rect 326732 117516 326788 117572
rect 327516 158508 327572 158564
rect 327628 188860 327684 188916
rect 329196 240268 329252 240324
rect 329084 238700 329140 238756
rect 328972 237580 329028 237636
rect 327964 233436 328020 233492
rect 328860 237244 328916 237300
rect 328636 230188 328692 230244
rect 327852 188860 327908 188916
rect 328524 191548 328580 191604
rect 327628 144060 327684 144116
rect 328412 188076 328468 188132
rect 327404 117516 327460 117572
rect 326732 116732 326788 116788
rect 323484 91532 323540 91588
rect 318332 90524 318388 90580
rect 326732 86492 326788 86548
rect 311612 84700 311668 84756
rect 288092 55580 288148 55636
rect 288092 51772 288148 51828
rect 288988 52668 289044 52724
rect 288988 51660 289044 51716
rect 293580 48636 293636 48692
rect 307916 48412 307972 48468
rect 322252 48524 322308 48580
rect 315084 48300 315140 48356
rect 300748 47740 300804 47796
rect 285964 41580 286020 41636
rect 281596 26012 281652 26068
rect 328636 186396 328692 186452
rect 328524 143612 328580 143668
rect 328972 236908 329028 236964
rect 328860 142268 328916 142324
rect 328972 235900 329028 235956
rect 328972 138908 329028 138964
rect 329084 134316 329140 134372
rect 329420 239820 329476 239876
rect 329532 231532 329588 231588
rect 329756 149436 329812 149492
rect 330204 380604 330260 380660
rect 330652 380828 330708 380884
rect 330428 380716 330484 380772
rect 330652 353836 330708 353892
rect 330428 340956 330484 341012
rect 330316 319116 330372 319172
rect 330540 309148 330596 309204
rect 330204 301868 330260 301924
rect 330428 308252 330484 308308
rect 330092 288988 330148 289044
rect 330428 287308 330484 287364
rect 330316 285628 330372 285684
rect 330092 260876 330148 260932
rect 330092 237692 330148 237748
rect 330204 256060 330260 256116
rect 330092 236572 330148 236628
rect 329980 197820 330036 197876
rect 329980 140812 330036 140868
rect 329868 137564 329924 137620
rect 330540 277564 330596 277620
rect 330652 308140 330708 308196
rect 330540 267148 330596 267204
rect 330540 263788 330596 263844
rect 330316 246876 330372 246932
rect 330428 252028 330484 252084
rect 330204 232764 330260 232820
rect 330428 160076 330484 160132
rect 330540 250348 330596 250404
rect 331100 388108 331156 388164
rect 336588 407372 336644 407428
rect 335356 394268 335412 394324
rect 335244 390572 335300 390628
rect 331548 387996 331604 388052
rect 332556 387996 332612 388052
rect 332108 386092 332164 386148
rect 331884 382172 331940 382228
rect 331212 365036 331268 365092
rect 331212 309148 331268 309204
rect 331772 361452 331828 361508
rect 331100 308252 331156 308308
rect 330988 294252 331044 294308
rect 331548 299180 331604 299236
rect 330876 289100 330932 289156
rect 330988 287308 331044 287364
rect 330988 274540 331044 274596
rect 330876 273308 330932 273364
rect 331548 268716 331604 268772
rect 330764 263788 330820 263844
rect 330876 258636 330932 258692
rect 331212 256956 331268 257012
rect 330764 250684 330820 250740
rect 331212 248668 331268 248724
rect 331660 250460 331716 250516
rect 331548 245196 331604 245252
rect 330988 242060 331044 242116
rect 331212 240268 331268 240324
rect 331660 239484 331716 239540
rect 331548 238588 331604 238644
rect 330988 232876 331044 232932
rect 330652 159964 330708 160020
rect 330988 231084 331044 231140
rect 330988 142604 331044 142660
rect 330540 138796 330596 138852
rect 331884 297500 331940 297556
rect 331996 349804 332052 349860
rect 331884 265468 331940 265524
rect 331884 256396 331940 256452
rect 331772 135884 331828 135940
rect 331884 246876 331940 246932
rect 330092 47964 330148 48020
rect 329196 22988 329252 23044
rect 328412 21756 328468 21812
rect 335132 383180 335188 383236
rect 332556 366828 332612 366884
rect 334908 383068 334964 383124
rect 334572 360556 334628 360612
rect 333228 359660 333284 359716
rect 332108 321356 332164 321412
rect 332220 348012 332276 348068
rect 332108 308364 332164 308420
rect 332108 158956 332164 159012
rect 331996 157612 332052 157668
rect 333004 340844 333060 340900
rect 332332 338156 332388 338212
rect 332332 305564 332388 305620
rect 332556 316988 332612 317044
rect 332556 298508 332612 298564
rect 332668 308252 332724 308308
rect 332444 297388 332500 297444
rect 332444 283724 332500 283780
rect 332556 296492 332612 296548
rect 332444 270956 332500 271012
rect 332332 264124 332388 264180
rect 332780 308028 332836 308084
rect 332780 290668 332836 290724
rect 332668 288876 332724 288932
rect 332780 268268 332836 268324
rect 332780 264012 332836 264068
rect 332668 261996 332724 262052
rect 332332 261436 332388 261492
rect 332556 261324 332612 261380
rect 332332 259420 332388 259476
rect 332444 254604 332500 254660
rect 332780 258860 332836 258916
rect 332668 256956 332724 257012
rect 332780 258412 332836 258468
rect 332668 249900 332724 249956
rect 332780 249452 332836 249508
rect 332332 243628 332388 243684
rect 332780 248556 332836 248612
rect 332780 243404 332836 243460
rect 332444 240268 332500 240324
rect 332668 238700 332724 238756
rect 332668 238476 332724 238532
rect 332668 236460 332724 236516
rect 332444 235900 332500 235956
rect 333004 157388 333060 157444
rect 333116 339052 333172 339108
rect 333452 354284 333508 354340
rect 333340 346220 333396 346276
rect 333340 308140 333396 308196
rect 333228 307916 333284 307972
rect 334460 351596 334516 351652
rect 334012 342636 334068 342692
rect 333788 341740 333844 341796
rect 333452 304444 333508 304500
rect 333676 305564 333732 305620
rect 333452 292236 333508 292292
rect 333340 264684 333396 264740
rect 333116 157500 333172 157556
rect 332220 156828 332276 156884
rect 332668 157164 332724 157220
rect 332668 156716 332724 156772
rect 333116 156268 333172 156324
rect 333228 243516 333284 243572
rect 333564 273644 333620 273700
rect 333564 263788 333620 263844
rect 333452 260876 333508 260932
rect 333676 258748 333732 258804
rect 333564 250684 333620 250740
rect 333452 246764 333508 246820
rect 333452 243516 333508 243572
rect 333340 239708 333396 239764
rect 333564 239596 333620 239652
rect 333228 156044 333284 156100
rect 333228 150892 333284 150948
rect 333452 223916 333508 223972
rect 333452 183036 333508 183092
rect 332668 144284 332724 144340
rect 332668 139020 332724 139076
rect 333900 339948 333956 340004
rect 334124 319116 334180 319172
rect 334236 303884 334292 303940
rect 334348 296492 334404 296548
rect 334236 295596 334292 295652
rect 334572 307356 334628 307412
rect 334684 336364 334740 336420
rect 334796 334348 334852 334404
rect 334796 303884 334852 303940
rect 334684 293916 334740 293972
rect 334796 295596 334852 295652
rect 334124 283836 334180 283892
rect 334236 276556 334292 276612
rect 334348 283724 334404 283780
rect 334908 285740 334964 285796
rect 335020 308924 335076 308980
rect 335468 390684 335524 390740
rect 335580 383964 335636 384020
rect 338604 409948 338660 410004
rect 338492 409612 338548 409668
rect 337484 409276 337540 409332
rect 336700 391692 336756 391748
rect 336700 391468 336756 391524
rect 336924 407820 336980 407876
rect 336588 383852 336644 383908
rect 336812 388220 336868 388276
rect 335580 334348 335636 334404
rect 336028 348908 336084 348964
rect 335468 327628 335524 327684
rect 335356 315756 335412 315812
rect 335244 308364 335300 308420
rect 335132 295372 335188 295428
rect 335244 303996 335300 304052
rect 335244 285516 335300 285572
rect 335356 298508 335412 298564
rect 335020 283836 335076 283892
rect 335916 297164 335972 297220
rect 335356 283836 335412 283892
rect 335468 293804 335524 293860
rect 334796 281372 334852 281428
rect 335356 282156 335412 282212
rect 334572 280812 334628 280868
rect 334572 275548 334628 275604
rect 334348 270956 334404 271012
rect 334124 270396 334180 270452
rect 335132 270396 335188 270452
rect 334348 269164 334404 269220
rect 334796 268940 334852 268996
rect 334572 258860 334628 258916
rect 334236 250460 334292 250516
rect 334012 157276 334068 157332
rect 334236 239820 334292 239876
rect 333900 157164 333956 157220
rect 333788 157052 333844 157108
rect 333900 156940 333956 156996
rect 333564 156380 333620 156436
rect 333564 155932 333620 155988
rect 333676 156268 333732 156324
rect 334572 230412 334628 230468
rect 334572 230188 334628 230244
rect 334236 154364 334292 154420
rect 335020 265468 335076 265524
rect 335020 259420 335076 259476
rect 334908 258748 334964 258804
rect 334908 246988 334964 247044
rect 335804 288988 335860 289044
rect 335692 277452 335748 277508
rect 335468 268828 335524 268884
rect 335580 277228 335636 277284
rect 335356 264684 335412 264740
rect 335244 259532 335300 259588
rect 335468 241164 335524 241220
rect 335468 238588 335524 238644
rect 335244 160300 335300 160356
rect 335356 191548 335412 191604
rect 335132 159516 335188 159572
rect 335580 159068 335636 159124
rect 335356 156380 335412 156436
rect 337260 407484 337316 407540
rect 337036 406252 337092 406308
rect 337036 389228 337092 389284
rect 337148 392812 337204 392868
rect 336924 383516 336980 383572
rect 336924 379820 336980 379876
rect 337036 386316 337092 386372
rect 336812 347340 336868 347396
rect 336812 340956 336868 341012
rect 336028 292236 336084 292292
rect 336700 297500 336756 297556
rect 336700 282380 336756 282436
rect 335916 267596 335972 267652
rect 336028 277340 336084 277396
rect 336588 275884 336644 275940
rect 336028 264124 336084 264180
rect 336140 266252 336196 266308
rect 335916 257068 335972 257124
rect 335916 250124 335972 250180
rect 335916 248780 335972 248836
rect 335916 245308 335972 245364
rect 336028 246988 336084 247044
rect 335916 244076 335972 244132
rect 335916 237244 335972 237300
rect 336252 264012 336308 264068
rect 336252 253148 336308 253204
rect 336140 238028 336196 238084
rect 336028 191548 336084 191604
rect 335804 156940 335860 156996
rect 335916 189756 335972 189812
rect 335692 152572 335748 152628
rect 334796 152460 334852 152516
rect 333900 147644 333956 147700
rect 333676 145964 333732 146020
rect 333564 138908 333620 138964
rect 333452 136892 333508 136948
rect 336028 181356 336084 181412
rect 336028 180124 336084 180180
rect 336028 177996 336084 178052
rect 336028 176988 336084 177044
rect 336028 152908 336084 152964
rect 336028 144284 336084 144340
rect 336588 151228 336644 151284
rect 336588 142380 336644 142436
rect 336924 334348 336980 334404
rect 337372 391468 337428 391524
rect 337484 386316 337540 386372
rect 337596 407708 337652 407764
rect 337372 373324 337428 373380
rect 337484 347340 337540 347396
rect 337260 269388 337316 269444
rect 337372 287420 337428 287476
rect 337372 265468 337428 265524
rect 337260 250236 337316 250292
rect 337260 247100 337316 247156
rect 337260 237916 337316 237972
rect 337148 236348 337204 236404
rect 337372 236684 337428 236740
rect 337260 224700 337316 224756
rect 337036 213948 337092 214004
rect 337148 217532 337204 217588
rect 337036 191436 337092 191492
rect 337372 223916 337428 223972
rect 337260 210924 337316 210980
rect 337148 181356 337204 181412
rect 337372 177996 337428 178052
rect 337036 168252 337092 168308
rect 336924 134316 336980 134372
rect 337036 143948 337092 144004
rect 338044 406812 338100 406868
rect 338044 399532 338100 399588
rect 338940 407596 338996 407652
rect 338604 399196 338660 399252
rect 338716 407036 338772 407092
rect 338492 389116 338548 389172
rect 338716 389004 338772 389060
rect 338828 403788 338884 403844
rect 339164 406924 339220 406980
rect 338940 399084 338996 399140
rect 339052 403452 339108 403508
rect 346332 410172 346388 410228
rect 340508 409164 340564 409220
rect 340284 408716 340340 408772
rect 339388 404124 339444 404180
rect 339836 405804 339892 405860
rect 339164 399420 339220 399476
rect 339276 403676 339332 403732
rect 340172 404908 340228 404964
rect 340060 396172 340116 396228
rect 339836 396060 339892 396116
rect 340284 396396 340340 396452
rect 340396 403228 340452 403284
rect 339948 392924 340004 392980
rect 339276 392700 339332 392756
rect 341852 407820 341908 407876
rect 342748 407260 342804 407316
rect 340620 405132 340676 405188
rect 342524 404796 342580 404852
rect 347004 409276 347060 409332
rect 478828 410396 478884 410452
rect 462364 410284 462420 410340
rect 352828 409836 352884 409892
rect 352940 410172 352996 410228
rect 352156 406700 352212 406756
rect 352828 409276 352884 409332
rect 358316 410172 358372 410228
rect 352940 408268 352996 408324
rect 352828 406588 352884 406644
rect 354732 406700 354788 406756
rect 354508 405244 354564 405300
rect 346332 404796 346388 404852
rect 347564 405020 347620 405076
rect 347564 404796 347620 404852
rect 354508 404348 354564 404404
rect 357868 408492 357924 408548
rect 366156 410172 366212 410228
rect 361788 409948 361844 410004
rect 361452 408380 361508 408436
rect 358316 407596 358372 407652
rect 358876 407708 358932 407764
rect 357868 406476 357924 406532
rect 357308 405356 357364 405412
rect 354732 404348 354788 404404
rect 361452 404348 361508 404404
rect 364700 408268 364756 408324
rect 369628 410172 369684 410228
rect 366156 408044 366212 408100
rect 367276 407596 367332 407652
rect 367276 407260 367332 407316
rect 366268 406700 366324 406756
rect 367612 404908 367668 404964
rect 367836 408380 367892 408436
rect 378812 410172 378868 410228
rect 369628 407708 369684 407764
rect 372988 410060 373044 410116
rect 372988 408156 373044 408212
rect 374668 408492 374724 408548
rect 372764 406588 372820 406644
rect 374668 406476 374724 406532
rect 367836 404908 367892 404964
rect 378812 409724 378868 409780
rect 379708 410172 379764 410228
rect 392252 410172 392308 410228
rect 379708 409052 379764 409108
rect 381052 408828 381108 408884
rect 382172 408492 382228 408548
rect 382172 407484 382228 407540
rect 383068 407484 383124 407540
rect 383180 407372 383236 407428
rect 383292 408716 383348 408772
rect 384748 408268 384804 408324
rect 388220 408044 388276 408100
rect 389676 410060 389732 410116
rect 384748 407596 384804 407652
rect 389676 407372 389732 407428
rect 383292 406476 383348 406532
rect 388444 407036 388500 407092
rect 383068 406364 383124 406420
rect 390572 407036 390628 407092
rect 377916 404460 377972 404516
rect 364700 404348 364756 404404
rect 460348 410172 460404 410228
rect 393372 410060 393428 410116
rect 398524 409724 398580 409780
rect 403228 409612 403284 409668
rect 403004 408492 403060 408548
rect 392252 406364 392308 406420
rect 398188 408380 398244 408436
rect 398188 405020 398244 405076
rect 398412 408268 398468 408324
rect 390572 404348 390628 404404
rect 395836 404348 395892 404404
rect 403004 407484 403060 407540
rect 403900 408380 403956 408436
rect 403900 406252 403956 406308
rect 403900 404908 403956 404964
rect 403900 404460 403956 404516
rect 398412 404348 398468 404404
rect 408828 409164 408884 409220
rect 419132 409276 419188 409332
rect 424956 409276 425012 409332
rect 420028 409164 420084 409220
rect 413980 408156 414036 408212
rect 418012 408604 418068 408660
rect 410620 406924 410676 406980
rect 420028 408156 420084 408212
rect 425404 408716 425460 408772
rect 432796 407036 432852 407092
rect 434588 406588 434644 406644
rect 429436 404684 429492 404740
rect 440188 406364 440244 406420
rect 439068 404684 439124 404740
rect 450044 409836 450100 409892
rect 455196 405580 455252 405636
rect 470652 408156 470708 408212
rect 465500 408044 465556 408100
rect 469756 407372 469812 407428
rect 475804 406140 475860 406196
rect 477148 408492 477204 408548
rect 478828 408156 478884 408212
rect 484540 408380 484596 408436
rect 486108 406028 486164 406084
rect 496412 409276 496468 409332
rect 491260 405692 491316 405748
rect 491932 408268 491988 408324
rect 499324 406588 499380 406644
rect 501564 406588 501620 406644
rect 506156 405916 506212 405972
rect 506716 406812 506772 406868
rect 511868 406588 511924 406644
rect 514108 406588 514164 406644
rect 517020 406588 517076 406644
rect 521500 407148 521556 407204
rect 522172 406588 522228 406644
rect 591164 409052 591220 409108
rect 573244 406700 573300 406756
rect 527324 405804 527380 405860
rect 528892 406588 528948 406644
rect 543676 406588 543732 406644
rect 551068 406588 551124 406644
rect 558236 406588 558292 406644
rect 580636 406588 580692 406644
rect 444892 404572 444948 404628
rect 590716 404460 590772 404516
rect 404012 404348 404068 404404
rect 536284 404348 536340 404404
rect 351484 404236 351540 404292
rect 373660 404236 373716 404292
rect 447580 404236 447636 404292
rect 454972 404236 455028 404292
rect 565852 404236 565908 404292
rect 590492 404012 590548 404068
rect 340620 397404 340676 397460
rect 585452 402332 585508 402388
rect 340508 395836 340564 395892
rect 585452 394828 585508 394884
rect 340396 392588 340452 392644
rect 339052 392476 339108 392532
rect 338828 382284 338884 382340
rect 337820 373996 337876 374052
rect 337596 275884 337652 275940
rect 337708 369516 337764 369572
rect 340284 368620 340340 368676
rect 339612 367724 339668 367780
rect 338044 364140 338100 364196
rect 337820 296492 337876 296548
rect 337932 352492 337988 352548
rect 339500 358764 339556 358820
rect 338044 288988 338100 289044
rect 338492 357868 338548 357924
rect 337932 277340 337988 277396
rect 337708 275660 337764 275716
rect 337820 276556 337876 276612
rect 337820 268940 337876 268996
rect 337932 270060 337988 270116
rect 337708 268828 337764 268884
rect 337708 260428 337764 260484
rect 337596 256396 337652 256452
rect 338380 263676 338436 263732
rect 337596 246876 337652 246932
rect 337932 257180 337988 257236
rect 338380 257068 338436 257124
rect 337708 240492 337764 240548
rect 337932 254940 337988 254996
rect 337932 248668 337988 248724
rect 338044 250124 338100 250180
rect 337932 245420 337988 245476
rect 337932 237804 337988 237860
rect 337708 236572 337764 236628
rect 338044 182252 338100 182308
rect 338380 177996 338436 178052
rect 337484 143948 337540 144004
rect 337596 165452 337652 165508
rect 337036 128604 337092 128660
rect 336812 127596 336868 127652
rect 338380 160972 338436 161028
rect 338492 157724 338548 157780
rect 338604 350700 338660 350756
rect 338716 345324 338772 345380
rect 338716 157836 338772 157892
rect 338828 304444 338884 304500
rect 338604 155148 338660 155204
rect 338940 296492 338996 296548
rect 338940 287420 338996 287476
rect 338940 277564 338996 277620
rect 339052 253596 339108 253652
rect 340172 356972 340228 357028
rect 339836 355180 339892 355236
rect 339724 337260 339780 337316
rect 339724 296492 339780 296548
rect 339612 287756 339668 287812
rect 339500 247100 339556 247156
rect 339724 253484 339780 253540
rect 339052 246988 339108 247044
rect 339500 246876 339556 246932
rect 338940 160188 338996 160244
rect 339052 241948 339108 242004
rect 338828 149324 338884 149380
rect 339500 241164 339556 241220
rect 339836 239820 339892 239876
rect 339948 291004 340004 291060
rect 339948 236684 340004 236740
rect 339724 229292 339780 229348
rect 339164 197708 339220 197764
rect 339164 171948 339220 172004
rect 339276 181356 339332 181412
rect 339276 161084 339332 161140
rect 339052 137452 339108 137508
rect 340284 155932 340340 155988
rect 340396 353052 340452 353108
rect 590604 394828 590660 394884
rect 590604 364140 590660 364196
rect 591164 403788 591220 403844
rect 590716 337596 590772 337652
rect 590492 324492 590548 324548
rect 585452 284620 585508 284676
rect 340620 197148 340676 197204
rect 340396 152684 340452 152740
rect 340620 183708 340676 183764
rect 340172 135772 340228 135828
rect 337596 57148 337652 57204
rect 337596 48636 337652 48692
rect 335916 22876 335972 22932
rect 331884 21644 331940 21700
rect 340620 21308 340676 21364
rect 523292 160412 523348 160468
rect 491932 160300 491988 160356
rect 506716 160188 506772 160244
rect 351148 159964 351204 160020
rect 358876 159516 358932 159572
rect 344092 157836 344148 157892
rect 373660 158508 373716 158564
rect 381052 157612 381108 157668
rect 366268 156828 366324 156884
rect 388444 155260 388500 155316
rect 410620 152684 410676 152740
rect 403228 152572 403284 152628
rect 395836 152460 395892 152516
rect 422604 159964 422660 160020
rect 418012 149324 418068 149380
rect 420812 157500 420868 157556
rect 420812 144396 420868 144452
rect 422380 145180 422436 145236
rect 422380 143836 422436 143892
rect 422268 143276 422324 143332
rect 421708 130956 421764 131012
rect 386204 128492 386260 128548
rect 379820 113484 379876 113540
rect 373548 106876 373604 106932
rect 375116 106764 375172 106820
rect 378028 104076 378084 104132
rect 376572 103180 376628 103236
rect 384524 108668 384580 108724
rect 381388 103964 381444 104020
rect 383180 103852 383236 103908
rect 387772 125132 387828 125188
rect 411180 113372 411236 113428
rect 395500 110572 395556 110628
rect 388668 103740 388724 103796
rect 390236 103628 390292 103684
rect 393372 103516 393428 103572
rect 391804 103404 391860 103460
rect 398636 110460 398692 110516
rect 396508 103292 396564 103348
rect 401772 110236 401828 110292
rect 400204 108332 400260 108388
rect 409612 110012 409668 110068
rect 404908 108444 404964 108500
rect 403228 103852 403284 103908
rect 407484 105308 407540 105364
rect 406700 103964 406756 104020
rect 412188 104972 412244 105028
rect 414092 104076 414148 104132
rect 415660 104076 415716 104132
rect 367052 84812 367108 84868
rect 367052 74956 367108 75012
rect 420140 77308 420196 77364
rect 367836 58268 367892 58324
rect 367836 57148 367892 57204
rect 419244 52108 419300 52164
rect 420028 51996 420084 52052
rect 420140 72380 420196 72436
rect 419244 51660 419300 51716
rect 420252 62524 420308 62580
rect 420252 51884 420308 51940
rect 422828 159964 422884 160020
rect 422604 143724 422660 143780
rect 422716 147756 422772 147812
rect 422716 144060 422772 144116
rect 422380 136892 422436 136948
rect 422380 135660 422436 135716
rect 422268 130956 422324 131012
rect 421820 122556 421876 122612
rect 421820 87164 421876 87220
rect 421708 57596 421764 57652
rect 421708 51772 421764 51828
rect 421820 68796 421876 68852
rect 421820 67452 421876 67508
rect 420140 50316 420196 50372
rect 422604 135660 422660 135716
rect 422604 77308 422660 77364
rect 425404 154364 425460 154420
rect 432796 151116 432852 151172
rect 423276 144060 423332 144116
rect 422828 143500 422884 143556
rect 423164 143724 423220 143780
rect 423388 143724 423444 143780
rect 423164 143164 423220 143220
rect 425852 141484 425908 141540
rect 425068 117516 425124 117572
rect 447580 157724 447636 157780
rect 454972 157500 455028 157556
rect 457772 157500 457828 157556
rect 457996 156268 458052 156324
rect 457772 135884 457828 135940
rect 457884 152572 457940 152628
rect 440188 135772 440244 135828
rect 462364 156268 462420 156324
rect 467852 159964 467908 160020
rect 457996 137564 458052 137620
rect 458220 153020 458276 153076
rect 466508 152460 466564 152516
rect 465388 147980 465444 148036
rect 458444 144508 458500 144564
rect 458220 137452 458276 137508
rect 458332 142828 458388 142884
rect 465388 140924 465444 140980
rect 466508 143836 466564 143892
rect 469532 155260 469588 155316
rect 477148 157500 477204 157556
rect 521500 158956 521556 159012
rect 514108 157500 514164 157556
rect 499324 156940 499380 156996
rect 484540 155820 484596 155876
rect 514892 155708 514948 155764
rect 469756 149436 469812 149492
rect 479052 152908 479108 152964
rect 469532 143724 469588 143780
rect 467852 143276 467908 143332
rect 468524 141708 468580 141764
rect 468524 141260 468580 141316
rect 471212 143500 471268 143556
rect 472108 143164 472164 143220
rect 474348 142828 474404 142884
rect 475916 141596 475972 141652
rect 510636 152348 510692 152404
rect 486892 151228 486948 151284
rect 483756 149548 483812 149604
rect 485324 141148 485380 141204
rect 499436 149660 499492 149716
rect 494732 147868 494788 147924
rect 488460 146300 488516 146356
rect 493164 146188 493220 146244
rect 490028 142828 490084 142884
rect 491596 141372 491652 141428
rect 497868 142828 497924 142884
rect 505596 146076 505652 146132
rect 504140 143948 504196 144004
rect 501676 142940 501732 142996
rect 480620 139692 480676 139748
rect 477484 139580 477540 139636
rect 482188 139580 482244 139636
rect 501004 139468 501060 139524
rect 502572 141260 502628 141316
rect 505596 143948 505652 144004
rect 512428 148988 512484 149044
rect 512428 144060 512484 144116
rect 516908 154028 516964 154084
rect 514892 143836 514948 143892
rect 516684 143948 516740 144004
rect 510636 143612 510692 143668
rect 515116 143724 515172 143780
rect 507500 143500 507556 143556
rect 505708 142828 505764 142884
rect 507276 142828 507332 142884
rect 510412 143388 510468 143444
rect 507500 141036 507556 141092
rect 508844 142828 508900 142884
rect 510748 143276 510804 143332
rect 510748 142716 510804 142772
rect 511980 142828 512036 142884
rect 513548 142828 513604 142884
rect 516908 143948 516964 144004
rect 519820 145068 519876 145124
rect 518252 142156 518308 142212
rect 521388 144508 521444 144564
rect 522956 144060 523012 144116
rect 528892 159068 528948 159124
rect 543676 160076 543732 160132
rect 558460 157612 558516 157668
rect 551068 156044 551124 156100
rect 536284 155932 536340 155988
rect 548044 155484 548100 155540
rect 535052 153916 535108 153972
rect 527660 150668 527716 150724
rect 523292 143948 523348 144004
rect 524524 148876 524580 148932
rect 526092 147532 526148 147588
rect 532364 150556 532420 150612
rect 530796 150444 530852 150500
rect 529228 150332 529284 150388
rect 533932 143836 533988 143892
rect 538636 145740 538692 145796
rect 535052 143836 535108 143892
rect 537068 143948 537124 144004
rect 535500 143276 535556 143332
rect 540204 145628 540260 145684
rect 541772 145516 541828 145572
rect 543340 145404 543396 145460
rect 544908 143724 544964 143780
rect 546476 143612 546532 143668
rect 575372 158844 575428 158900
rect 574812 157388 574868 157444
rect 573244 156156 573300 156212
rect 574588 157276 574644 157332
rect 565852 152572 565908 152628
rect 562156 152236 562212 152292
rect 552748 147420 552804 147476
rect 551180 147084 551236 147140
rect 549612 141932 549668 141988
rect 559020 147308 559076 147364
rect 555884 147196 555940 147252
rect 554316 142940 554372 142996
rect 557452 146972 557508 147028
rect 560588 143836 560644 143892
rect 565292 151004 565348 151060
rect 563724 143500 563780 143556
rect 568428 148652 568484 148708
rect 566860 145292 566916 145348
rect 501676 139468 501732 139524
rect 496300 139244 496356 139300
rect 458444 137676 458500 137732
rect 458332 135660 458388 135716
rect 457884 134092 457940 134148
rect 574588 133980 574644 134036
rect 574700 153804 574756 153860
rect 425852 117516 425908 117572
rect 425068 116732 425124 116788
rect 574812 129948 574868 130004
rect 574924 152012 574980 152068
rect 575148 148764 575204 148820
rect 574924 111804 574980 111860
rect 575036 131852 575092 131908
rect 574700 107436 574756 107492
rect 575260 147644 575316 147700
rect 575260 119308 575316 119364
rect 575148 117292 575204 117348
rect 575036 101724 575092 101780
rect 578172 158732 578228 158788
rect 576492 157164 576548 157220
rect 576268 157052 576324 157108
rect 575596 140700 575652 140756
rect 575372 99148 575428 99204
rect 575484 138684 575540 138740
rect 458556 99036 458612 99092
rect 457772 98812 457828 98868
rect 457436 98700 457492 98756
rect 457660 98364 457716 98420
rect 457660 95116 457716 95172
rect 457436 91756 457492 91812
rect 425068 82236 425124 82292
rect 423164 72380 423220 72436
rect 458444 97580 458500 97636
rect 458444 81676 458500 81732
rect 575596 131852 575652 131908
rect 576268 131404 576324 131460
rect 576380 138908 576436 138964
rect 576492 127372 576548 127428
rect 576604 150892 576660 150948
rect 576380 123340 576436 123396
rect 576828 140812 576884 140868
rect 576604 121324 576660 121380
rect 576716 140476 576772 140532
rect 576716 115276 576772 115332
rect 577948 140588 578004 140644
rect 576828 103180 576884 103236
rect 576940 140364 576996 140420
rect 577948 135436 578004 135492
rect 578060 138796 578116 138852
rect 576940 95116 576996 95172
rect 575484 93100 575540 93156
rect 458556 78316 458612 78372
rect 457772 71596 457828 71652
rect 587132 244972 587188 245028
rect 585452 155260 585508 155316
rect 585564 205324 585620 205380
rect 580636 152796 580692 152852
rect 587132 160860 587188 160916
rect 590380 178892 590436 178948
rect 591276 159628 591332 159684
rect 590380 159180 590436 159236
rect 585564 152460 585620 152516
rect 578396 147980 578452 148036
rect 578284 142044 578340 142100
rect 578284 109228 578340 109284
rect 578172 105196 578228 105252
rect 578060 68908 578116 68964
rect 422940 68796 422996 68852
rect 579628 145964 579684 146020
rect 579628 125356 579684 125412
rect 581308 140252 581364 140308
rect 581308 97132 581364 97188
rect 578396 62860 578452 62916
rect 422716 62524 422772 62580
rect 422492 52668 422548 52724
rect 421820 50204 421876 50260
rect 578620 48748 578676 48804
rect 578508 46732 578564 46788
rect 578172 42700 578228 42756
rect 367836 24556 367892 24612
rect 577948 30604 578004 30660
rect 574588 23996 574644 24052
rect 574588 21308 574644 21364
rect 340956 21196 341012 21252
rect 577948 21196 578004 21252
rect 578284 38668 578340 38724
rect 578284 22988 578340 23044
rect 578396 34636 578452 34692
rect 578508 21756 578564 21812
rect 578620 21644 578676 21700
rect 578396 21420 578452 21476
rect 578172 20076 578228 20132
rect 582540 7644 582596 7700
rect 273980 4284 274036 4340
rect 580636 7532 580692 7588
rect 270508 4172 270564 4228
rect 584444 5852 584500 5908
<< metal3 >>
rect 189522 591276 189532 591332
rect 189588 591276 297836 591332
rect 297892 591276 297902 591332
rect 202962 591164 202972 591220
rect 203028 591164 319900 591220
rect 319956 591164 319966 591220
rect 189634 591052 189644 591108
rect 189700 591052 364028 591108
rect 364084 591052 364094 591108
rect 186162 590940 186172 590996
rect 186228 590940 430220 590996
rect 430276 590940 430286 590996
rect 203186 590828 203196 590884
rect 203252 590828 452284 590884
rect 452340 590828 452350 590884
rect 186386 590716 186396 590772
rect 186452 590716 496412 590772
rect 496468 590716 496478 590772
rect 99474 590604 99484 590660
rect 99540 590604 152012 590660
rect 152068 590604 152078 590660
rect 203074 590604 203084 590660
rect 203140 590604 518476 590660
rect 518532 590604 518542 590660
rect 33282 590492 33292 590548
rect 33348 590492 160412 590548
rect 160468 590492 160478 590548
rect 165666 590492 165676 590548
rect 165732 590492 177212 590548
rect 177268 590492 177278 590548
rect 186274 590492 186284 590548
rect 186340 590492 562604 590548
rect 562660 590492 562670 590548
rect 189746 590380 189756 590436
rect 189812 590380 231644 590436
rect 231700 590380 231710 590436
rect 187730 590156 187740 590212
rect 187796 590156 188972 590212
rect 189028 590156 189038 590212
rect 253670 590156 253708 590212
rect 253764 590156 253774 590212
rect 341058 590156 341068 590212
rect 341124 590156 341964 590212
rect 342020 590156 342030 590212
rect 77410 588812 77420 588868
rect 77476 588812 165452 588868
rect 165508 588812 165518 588868
rect 180002 588812 180012 588868
rect 180068 588812 408268 588868
rect 408324 588812 408334 588868
rect 595560 588644 597000 588840
rect 590482 588588 590492 588644
rect 590548 588616 597000 588644
rect 590548 588588 595672 588616
rect -960 587188 480 587384
rect 202850 587244 202860 587300
rect 202916 587244 386092 587300
rect 386148 587244 386158 587300
rect -960 587160 4956 587188
rect 392 587132 4956 587160
rect 5012 587132 5022 587188
rect 196466 587132 196476 587188
rect 196532 587132 584668 587188
rect 584724 587132 584734 587188
rect 143378 583884 143388 583940
rect 143444 583884 170492 583940
rect 170548 583884 170558 583940
rect 4946 583772 4956 583828
rect 5012 583772 153692 583828
rect 153748 583772 153758 583828
rect 179666 583772 179676 583828
rect 179732 583772 209580 583828
rect 209636 583772 209646 583828
rect 121314 582092 121324 582148
rect 121380 582092 155372 582148
rect 155428 582092 155438 582148
rect 172946 578732 172956 578788
rect 173012 578732 474348 578788
rect 474404 578732 474414 578788
rect 172834 577052 172844 577108
rect 172900 577052 540540 577108
rect 540596 577052 540606 577108
rect 189298 576492 189308 576548
rect 189364 576492 529676 576548
rect 529732 576492 529742 576548
rect 189410 576380 189420 576436
rect 189476 576380 532588 576436
rect 532644 576380 532654 576436
rect 202738 576268 202748 576324
rect 202804 576268 590828 576324
rect 590884 576268 590894 576324
rect 595560 575428 597000 575624
rect 189186 575372 189196 575428
rect 189252 575400 597000 575428
rect 189252 575372 595672 575400
rect 190418 575148 190428 575204
rect 190484 575148 478828 575204
rect 478884 575148 478894 575204
rect 188962 575036 188972 575092
rect 189028 575036 480620 575092
rect 480676 575036 480686 575092
rect 189410 574924 189420 574980
rect 189476 574924 530124 574980
rect 530180 574924 530190 574980
rect 189298 574812 189308 574868
rect 189364 574812 532812 574868
rect 532868 574812 532878 574868
rect 201170 574700 201180 574756
rect 201236 574700 591164 574756
rect 591220 574700 591230 574756
rect 198034 574588 198044 574644
rect 198100 574588 590604 574644
rect 590660 574588 590670 574644
rect 200610 573804 200620 573860
rect 200676 573804 478940 573860
rect 478996 573804 479006 573860
rect 198258 573692 198268 573748
rect 198324 573692 480508 573748
rect 480564 573692 480574 573748
rect 199602 573580 199612 573636
rect 199668 573580 532924 573636
rect 532980 573580 532990 573636
rect 197810 573468 197820 573524
rect 197876 573468 533372 573524
rect 533428 573468 533438 573524
rect 197698 573356 197708 573412
rect 197764 573356 533260 573412
rect 533316 573356 533326 573412
rect -960 573076 480 573272
rect 192882 573244 192892 573300
rect 192948 573244 529452 573300
rect 529508 573244 529518 573300
rect 196242 573132 196252 573188
rect 196308 573132 532812 573188
rect 532868 573132 532878 573188
rect -960 573048 52892 573076
rect 392 573020 52892 573048
rect 52948 573020 52958 573076
rect 187954 573020 187964 573076
rect 188020 573020 529676 573076
rect 529732 573020 529742 573076
rect 184706 572908 184716 572964
rect 184772 572908 529340 572964
rect 529396 572908 529406 572964
rect 193106 572124 193116 572180
rect 193172 572124 479052 572180
rect 479108 572124 479118 572180
rect 200946 572012 200956 572068
rect 201012 572012 529564 572068
rect 529620 572012 529630 572068
rect 201058 571900 201068 571956
rect 201124 571900 533484 571956
rect 533540 571900 533550 571956
rect 201282 571788 201292 571844
rect 201348 571788 533260 571844
rect 533316 571788 533326 571844
rect 199378 571676 199388 571732
rect 199444 571676 532700 571732
rect 532756 571676 532766 571732
rect 197922 571564 197932 571620
rect 197988 571564 533036 571620
rect 533092 571564 533102 571620
rect 192994 571452 193004 571508
rect 193060 571452 531132 571508
rect 531188 571452 531198 571508
rect 199826 571340 199836 571396
rect 199892 571340 590716 571396
rect 590772 571340 590782 571396
rect 192658 571228 192668 571284
rect 192724 571228 590940 571284
rect 590996 571228 591006 571284
rect 179554 570444 179564 570500
rect 179620 570444 275772 570500
rect 275828 570444 275838 570500
rect 193778 570332 193788 570388
rect 193844 570332 200620 570388
rect 200676 570332 200686 570388
rect 252018 570332 252028 570388
rect 252084 570332 479164 570388
rect 479220 570332 479230 570388
rect 203522 570220 203532 570276
rect 203588 570220 533036 570276
rect 533092 570220 533102 570276
rect 202514 570108 202524 570164
rect 202580 570108 532700 570164
rect 532756 570108 532766 570164
rect 201506 569996 201516 570052
rect 201572 569996 533148 570052
rect 533204 569996 533214 570052
rect 192546 569884 192556 569940
rect 192612 569884 198268 569940
rect 198324 569884 198334 569940
rect 199490 569884 199500 569940
rect 199556 569884 532588 569940
rect 532644 569884 532654 569940
rect 196354 569772 196364 569828
rect 196420 569772 529564 569828
rect 529620 569772 529630 569828
rect 189186 569660 189196 569716
rect 189252 569660 530012 569716
rect 530068 569660 530078 569716
rect 188066 569548 188076 569604
rect 188132 569548 530908 569604
rect 530964 569548 530974 569604
rect 196018 568652 196028 568708
rect 196084 568652 252028 568708
rect 252084 568652 252094 568708
rect 202626 568540 202636 568596
rect 202692 568540 532924 568596
rect 532980 568540 532990 568596
rect 195906 568428 195916 568484
rect 195972 568428 529340 568484
rect 529396 568428 529406 568484
rect 196130 568316 196140 568372
rect 196196 568316 529900 568372
rect 529956 568316 529966 568372
rect 192770 568204 192780 568260
rect 192836 568204 529788 568260
rect 529844 568204 529854 568260
rect 200722 568092 200732 568148
rect 200788 568092 590716 568148
rect 590772 568092 590782 568148
rect 198146 567980 198156 568036
rect 198212 567980 590492 568036
rect 590548 567980 590558 568036
rect 189522 567868 189532 567924
rect 189588 567868 591052 567924
rect 591108 567868 591118 567924
rect 187730 567308 187740 567364
rect 187796 567308 194012 567364
rect 194068 567308 194078 567364
rect 199266 567308 199276 567364
rect 199332 567308 479276 567364
rect 479332 567308 479342 567364
rect 191314 567196 191324 567252
rect 191380 567196 530236 567252
rect 530292 567196 530302 567252
rect 189074 567084 189084 567140
rect 189140 567084 190932 567140
rect 191426 567084 191436 567140
rect 191492 567084 193788 567140
rect 193844 567084 193854 567140
rect 194002 567084 194012 567140
rect 194068 567084 529452 567140
rect 529508 567084 529518 567140
rect 190876 567028 190932 567084
rect 189858 566972 189868 567028
rect 189924 566972 190428 567028
rect 190484 566972 190494 567028
rect 190876 566972 531020 567028
rect 531076 566972 531086 567028
rect 188850 566076 188860 566132
rect 188916 566076 189868 566132
rect 189924 566076 189934 566132
rect 187842 565068 187852 565124
rect 187908 565068 190120 565124
rect 529928 565068 532812 565124
rect 532868 565068 532878 565124
rect 532802 564844 532812 564900
rect 532868 564844 533260 564900
rect 533316 564844 533326 564900
rect 591154 562380 591164 562436
rect 591220 562408 595672 562436
rect 591220 562380 597000 562408
rect 595560 562184 597000 562380
rect 529928 560364 532588 560420
rect 532644 560364 532654 560420
rect -960 558964 480 559160
rect -960 558936 4396 558964
rect 392 558908 4396 558936
rect 4452 558908 4462 558964
rect 187618 557900 187628 557956
rect 187684 557900 190120 557956
rect 529928 555660 533036 555716
rect 533092 555660 533102 555716
rect 529928 550956 532924 551012
rect 532980 550956 532990 551012
rect 184706 550732 184716 550788
rect 184772 550732 190120 550788
rect 590818 549164 590828 549220
rect 590884 549192 595672 549220
rect 590884 549164 597000 549192
rect 595560 548968 597000 549164
rect 529928 546252 532812 546308
rect 532868 546252 532878 546308
rect -960 544852 480 545048
rect -960 544824 4172 544852
rect 392 544796 4172 544824
rect 4228 544796 4238 544852
rect 184594 543564 184604 543620
rect 184660 543564 190120 543620
rect 529928 541548 532700 541604
rect 532756 541548 532766 541604
rect 529928 536844 532588 536900
rect 532644 536844 532654 536900
rect 183026 536396 183036 536452
rect 183092 536396 190120 536452
rect 595560 535892 597000 535976
rect 591042 535836 591052 535892
rect 591108 535836 597000 535892
rect 595560 535752 597000 535836
rect 529554 532140 529564 532196
rect 529620 532140 529630 532196
rect -960 530740 480 530936
rect -960 530712 57932 530740
rect 392 530684 57932 530712
rect 57988 530684 57998 530740
rect 184594 529228 184604 529284
rect 184660 529228 190120 529284
rect 529928 527436 533372 527492
rect 533428 527436 533438 527492
rect 529928 522732 533260 522788
rect 533316 522732 533326 522788
rect 590818 522732 590828 522788
rect 590884 522760 595672 522788
rect 590884 522732 597000 522760
rect 595560 522536 597000 522732
rect 186386 522060 186396 522116
rect 186452 522060 190120 522116
rect 529928 518028 533148 518084
rect 533204 518028 533214 518084
rect -960 516628 480 516824
rect -960 516600 4508 516628
rect 392 516572 4508 516600
rect 4564 516572 4574 516628
rect 184482 514892 184492 514948
rect 184548 514892 190120 514948
rect 529928 513324 533036 513380
rect 533092 513324 533102 513380
rect 590706 509516 590716 509572
rect 590772 509544 595672 509572
rect 590772 509516 597000 509544
rect 595560 509320 597000 509516
rect 529442 508620 529452 508676
rect 529508 508620 529518 508676
rect 180450 507724 180460 507780
rect 180516 507724 190120 507780
rect 529928 503916 532924 503972
rect 532980 503916 532990 503972
rect -960 502516 480 502712
rect -960 502488 4284 502516
rect 392 502460 4284 502488
rect 4340 502460 4350 502516
rect 180562 500556 180572 500612
rect 180628 500556 190120 500612
rect 529928 499212 532812 499268
rect 532868 499212 532878 499268
rect 590594 496300 590604 496356
rect 590660 496328 595672 496356
rect 590660 496300 597000 496328
rect 595560 496104 597000 496300
rect 529330 494508 529340 494564
rect 529396 494508 529406 494564
rect 187282 493388 187292 493444
rect 187348 493388 190120 493444
rect 529666 489804 529676 489860
rect 529732 489804 529742 489860
rect -960 488404 480 488600
rect -960 488376 12572 488404
rect 392 488348 12572 488376
rect 12628 488348 12638 488404
rect 188066 486220 188076 486276
rect 188132 486220 190120 486276
rect 529928 485100 530124 485156
rect 530180 485100 530190 485156
rect 590930 483084 590940 483140
rect 590996 483112 595672 483140
rect 590996 483084 597000 483112
rect 595560 482888 597000 483084
rect 529928 480396 530124 480452
rect 530180 480396 530190 480452
rect 187170 479052 187180 479108
rect 187236 479052 190120 479108
rect 529890 476252 529900 476308
rect 529956 476252 529966 476308
rect 529900 475720 529956 476252
rect -960 474292 480 474488
rect -960 474264 4620 474292
rect 392 474236 4620 474264
rect 4676 474236 4686 474292
rect 187954 471884 187964 471940
rect 188020 471884 190120 471940
rect 529928 470988 532700 471044
rect 532756 470988 532766 471044
rect 590482 469868 590492 469924
rect 590548 469896 595672 469924
rect 590548 469868 597000 469896
rect 595560 469672 597000 469868
rect 4386 469532 4396 469588
rect 4452 469532 167132 469588
rect 167188 469532 167198 469588
rect 4498 467852 4508 467908
rect 4564 467852 168812 467908
rect 168868 467852 168878 467908
rect 529928 466284 533148 466340
rect 533204 466284 533214 466340
rect 4610 466172 4620 466228
rect 4676 466172 170492 466228
rect 170548 466172 170558 466228
rect 187842 464716 187852 464772
rect 187908 464716 190120 464772
rect 529778 461916 529788 461972
rect 529844 461916 529854 461972
rect 529788 461608 529844 461916
rect -960 460180 480 460376
rect -960 460152 4508 460180
rect 392 460124 4508 460152
rect 4564 460124 4574 460180
rect 187730 457548 187740 457604
rect 187796 457548 190120 457604
rect 529666 456988 529676 457044
rect 529732 456988 529742 457044
rect 529676 456904 529732 456988
rect 590706 456652 590716 456708
rect 590772 456680 595672 456708
rect 590772 456652 597000 456680
rect 595560 456456 597000 456652
rect 529554 452732 529564 452788
rect 529620 452732 529630 452788
rect 529564 452200 529620 452732
rect 187394 450380 187404 450436
rect 187460 450380 190120 450436
rect 529330 448028 529340 448084
rect 529396 448028 529406 448084
rect 529340 447496 529396 448028
rect -960 446068 480 446264
rect -960 446040 94892 446068
rect 392 446012 94892 446040
rect 94948 446012 94958 446068
rect 590594 443436 590604 443492
rect 590660 443464 595672 443492
rect 590660 443436 597000 443464
rect 529442 443324 529452 443380
rect 529508 443324 529518 443380
rect 187506 443212 187516 443268
rect 187572 443212 190120 443268
rect 529452 442792 529508 443324
rect 595560 443240 597000 443436
rect 529928 438060 531132 438116
rect 531188 438060 531198 438116
rect 187618 436044 187628 436100
rect 187684 436044 190120 436100
rect 529928 433356 530236 433412
rect 530292 433356 530302 433412
rect -960 431956 480 432152
rect -960 431928 162092 431956
rect 392 431900 162092 431928
rect 162148 431900 162158 431956
rect 595560 430164 597000 430248
rect 591266 430108 591276 430164
rect 591332 430108 597000 430164
rect 595560 430024 597000 430108
rect 189074 428876 189084 428932
rect 189140 428876 190120 428932
rect 529928 428652 532588 428708
rect 532644 428652 532654 428708
rect 529928 423948 531020 424004
rect 531076 423948 531086 424004
rect 186274 421708 186284 421764
rect 186340 421708 190120 421764
rect 529928 419244 530908 419300
rect 530964 419244 530974 419300
rect -960 417844 480 418040
rect -960 417816 4172 417844
rect 392 417788 4172 417816
rect 4228 417788 4238 417844
rect 68562 417452 68572 417508
rect 68628 417452 85260 417508
rect 85316 417452 85326 417508
rect 73042 417340 73052 417396
rect 73108 417340 182252 417396
rect 182308 417340 182318 417396
rect 70802 417228 70812 417284
rect 70868 417228 90076 417284
rect 90132 417228 90142 417284
rect 75282 417116 75292 417172
rect 75348 417116 85036 417172
rect 85092 417116 85102 417172
rect 66322 417004 66332 417060
rect 66388 417004 86828 417060
rect 86884 417004 86894 417060
rect 590482 417004 590492 417060
rect 590548 417032 595672 417060
rect 590548 417004 597000 417032
rect 64082 416892 64092 416948
rect 64148 416892 88284 416948
rect 88340 416892 88350 416948
rect 77522 416780 77532 416836
rect 77588 416780 180572 416836
rect 180628 416780 180638 416836
rect 595560 416808 597000 417004
rect 79762 416668 79772 416724
rect 79828 416668 86492 416724
rect 86548 416668 86558 416724
rect 185602 414540 185612 414596
rect 185668 414540 190120 414596
rect 529928 414540 533484 414596
rect 533540 414540 533550 414596
rect 55122 414092 55132 414148
rect 55188 414092 182364 414148
rect 182420 414092 182430 414148
rect 62038 413420 62076 413476
rect 62132 413420 62142 413476
rect 82226 413420 82236 413476
rect 82292 413420 84812 413476
rect 84868 413420 84878 413476
rect 83944 411964 183932 412020
rect 183988 411964 183998 412020
rect 189522 410508 189532 410564
rect 189588 410508 203756 410564
rect 203812 410508 203822 410564
rect 480470 410508 480508 410564
rect 480564 410508 480574 410564
rect 352818 410396 352828 410452
rect 352884 410396 359884 410452
rect 359940 410396 359950 410452
rect 478818 410396 478828 410452
rect 478884 410396 480620 410452
rect 480676 410396 480686 410452
rect 339378 410284 339388 410340
rect 339444 410284 462364 410340
rect 462420 410284 462430 410340
rect 346322 410172 346332 410228
rect 346388 410172 352940 410228
rect 352996 410172 353006 410228
rect 358306 410172 358316 410228
rect 358372 410172 366156 410228
rect 366212 410172 366222 410228
rect 369618 410172 369628 410228
rect 369684 410172 378812 410228
rect 378868 410172 378878 410228
rect 379698 410172 379708 410228
rect 379764 410172 392252 410228
rect 392308 410172 392318 410228
rect 460338 410172 460348 410228
rect 460404 410172 479164 410228
rect 479220 410172 479230 410228
rect 238018 410060 238028 410116
rect 238084 410060 351316 410116
rect 359538 410060 359548 410116
rect 359604 410060 366212 410116
rect 372978 410060 372988 410116
rect 373044 410060 389676 410116
rect 389732 410060 389742 410116
rect 393362 410060 393372 410116
rect 393428 410060 478940 410116
rect 478996 410060 479006 410116
rect 351260 410004 351316 410060
rect 188962 409948 188972 410004
rect 189028 409948 192332 410004
rect 192388 409948 192398 410004
rect 202290 409948 202300 410004
rect 202356 409948 273756 410004
rect 273812 409948 273822 410004
rect 338594 409948 338604 410004
rect 338660 409948 347732 410004
rect 351260 409948 361788 410004
rect 361844 409948 361854 410004
rect 347676 409892 347732 409948
rect 366156 409892 366212 410060
rect 83906 409836 83916 409892
rect 83972 409836 310940 409892
rect 310996 409836 311006 409892
rect 347676 409836 352828 409892
rect 352884 409836 352894 409892
rect 366156 409836 386204 409892
rect 386260 409836 386270 409892
rect 404898 409836 404908 409892
rect 404964 409836 450044 409892
rect 450100 409836 450110 409892
rect 192658 409724 192668 409780
rect 192724 409724 200732 409780
rect 200788 409724 200798 409780
rect 202962 409724 202972 409780
rect 203028 409724 206556 409780
rect 206612 409724 206622 409780
rect 207890 409724 207900 409780
rect 207956 409724 352828 409780
rect 352884 409724 352894 409780
rect 359650 409724 359660 409780
rect 359716 409724 366268 409780
rect 366324 409724 366334 409780
rect 378802 409724 378812 409780
rect 378868 409724 398524 409780
rect 398580 409724 398590 409780
rect 188962 409612 188972 409668
rect 189028 409612 274652 409668
rect 274708 409612 274876 409668
rect 274932 409612 274942 409668
rect 338482 409612 338492 409668
rect 338548 409612 403228 409668
rect 403284 409612 403294 409668
rect 202850 409500 202860 409556
rect 202916 409500 259420 409556
rect 259476 409500 259486 409556
rect 188850 409388 188860 409444
rect 188916 409388 202524 409444
rect 202580 409388 202590 409444
rect 203074 409388 203084 409444
rect 203140 409388 249116 409444
rect 249172 409388 249788 409444
rect 249844 409388 249854 409444
rect 201170 409276 201180 409332
rect 201236 409276 238812 409332
rect 238868 409276 240268 409332
rect 240324 409276 240334 409332
rect 259410 409276 259420 409332
rect 259476 409276 261996 409332
rect 262052 409276 262062 409332
rect 337474 409276 337484 409332
rect 337540 409276 347004 409332
rect 347060 409276 347070 409332
rect 352818 409276 352828 409332
rect 352884 409276 419132 409332
rect 419188 409276 419198 409332
rect 424946 409276 424956 409332
rect 425012 409276 478828 409332
rect 478884 409276 478894 409332
rect 496374 409276 496412 409332
rect 496468 409276 496478 409332
rect 201058 409164 201068 409220
rect 201124 409164 238700 409220
rect 238756 409164 238766 409220
rect 340498 409164 340508 409220
rect 340564 409164 408828 409220
rect 408884 409164 408894 409220
rect 420018 409164 420028 409220
rect 420084 409164 479052 409220
rect 479108 409164 479118 409220
rect 83944 409052 87276 409108
rect 87332 409052 87342 409108
rect 200722 409052 200732 409108
rect 200788 409052 204988 409108
rect 205044 409052 205054 409108
rect 208292 409052 264908 409108
rect 264964 409052 264974 409108
rect 291778 409052 291788 409108
rect 291844 409052 379708 409108
rect 379764 409052 379774 409108
rect 386082 409052 386092 409108
rect 386148 409052 591164 409108
rect 591220 409052 591230 409108
rect 208292 408996 208348 409052
rect 199266 408940 199276 408996
rect 199332 408940 208348 408996
rect 366034 408940 366044 408996
rect 366100 408940 369628 408996
rect 369684 408940 369694 408996
rect 286402 408828 286412 408884
rect 286468 408828 381052 408884
rect 381108 408828 381118 408884
rect 340274 408716 340284 408772
rect 340340 408716 361228 408772
rect 383282 408716 383292 408772
rect 383348 408716 425404 408772
rect 425460 408716 425470 408772
rect 302530 408604 302540 408660
rect 302596 408604 354508 408660
rect 354564 408604 354574 408660
rect 361172 408548 361228 408716
rect 374658 408604 374668 408660
rect 374724 408604 418012 408660
rect 418068 408604 418078 408660
rect 356178 408492 356188 408548
rect 356244 408492 357868 408548
rect 357924 408492 357934 408548
rect 361172 408492 374668 408548
rect 374724 408492 374734 408548
rect 382162 408492 382172 408548
rect 382228 408492 384860 408548
rect 384916 408492 384926 408548
rect 402994 408492 403004 408548
rect 403060 408492 477148 408548
rect 477204 408492 477214 408548
rect 289762 408380 289772 408436
rect 289828 408380 361452 408436
rect 361508 408380 361518 408436
rect 367826 408380 367836 408436
rect 367892 408380 398188 408436
rect 398244 408380 398254 408436
rect 403890 408380 403900 408436
rect 403956 408380 484540 408436
rect 484596 408380 484606 408436
rect 352930 408268 352940 408324
rect 352996 408268 364700 408324
rect 364756 408268 364766 408324
rect 384738 408268 384748 408324
rect 384804 408268 393484 408324
rect 393540 408268 393550 408324
rect 398402 408268 398412 408324
rect 398468 408268 491932 408324
rect 491988 408268 491998 408324
rect 366146 408156 366156 408212
rect 366212 408156 372988 408212
rect 373044 408156 373054 408212
rect 413970 408156 413980 408212
rect 414036 408156 420028 408212
rect 420084 408156 420094 408212
rect 470642 408156 470652 408212
rect 470708 408156 478828 408212
rect 478884 408156 478894 408212
rect 182354 408044 182364 408100
rect 182420 408044 284732 408100
rect 284788 408044 284798 408100
rect 288082 408044 288092 408100
rect 288148 408044 305788 408100
rect 305844 408044 305854 408100
rect 366146 408044 366156 408100
rect 366212 408044 388220 408100
rect 388276 408044 388286 408100
rect 465490 408044 465500 408100
rect 465556 408044 479276 408100
rect 479332 408044 479342 408100
rect 206546 407932 206556 407988
rect 206612 407932 264572 407988
rect 264628 407932 264638 407988
rect 273746 407932 273756 407988
rect 273812 407932 294812 407988
rect 294868 407932 294878 407988
rect 195906 407820 195916 407876
rect 195972 407820 261548 407876
rect 261604 407820 261614 407876
rect 278898 407820 278908 407876
rect 278964 407820 299964 407876
rect 300020 407820 300030 407876
rect 336914 407820 336924 407876
rect 336980 407820 341852 407876
rect 341908 407820 341918 407876
rect 199378 407708 199388 407764
rect 199444 407708 254828 407764
rect 254884 407708 254894 407764
rect 261986 407708 261996 407764
rect 262052 407708 337596 407764
rect 337652 407708 337662 407764
rect 342626 407708 342636 407764
rect 342692 407708 358876 407764
rect 358932 407708 358942 407764
rect 362786 407708 362796 407764
rect 362852 407708 369628 407764
rect 369684 407708 369694 407764
rect 172162 407596 172172 407652
rect 172228 407596 202748 407652
rect 202804 407596 202814 407652
rect 249778 407596 249788 407652
rect 249844 407596 328524 407652
rect 328580 407596 328590 407652
rect 338930 407596 338940 407652
rect 338996 407596 358316 407652
rect 358372 407596 358382 407652
rect 358530 407596 358540 407652
rect 358596 407596 367108 407652
rect 367266 407596 367276 407652
rect 367332 407596 384748 407652
rect 384804 407596 384814 407652
rect 367052 407540 367108 407596
rect 87266 407484 87276 407540
rect 87332 407484 163660 407540
rect 163716 407484 163726 407540
rect 197586 407484 197596 407540
rect 197652 407484 253484 407540
rect 253540 407484 253550 407540
rect 253698 407484 253708 407540
rect 253764 407484 254268 407540
rect 254324 407484 337260 407540
rect 337316 407484 337326 407540
rect 350466 407484 350476 407540
rect 350532 407484 362796 407540
rect 362852 407484 362862 407540
rect 367052 407484 382172 407540
rect 382228 407484 382238 407540
rect 383058 407484 383068 407540
rect 383124 407484 403004 407540
rect 403060 407484 403070 407540
rect 155362 407372 155372 407428
rect 155428 407372 277228 407428
rect 277284 407372 280028 407428
rect 280084 407372 280094 407428
rect 336578 407372 336588 407428
rect 336644 407372 383180 407428
rect 383236 407372 383246 407428
rect 389666 407372 389676 407428
rect 389732 407372 469756 407428
rect 469812 407372 469822 407428
rect 232306 407260 232316 407316
rect 232372 407260 233660 407316
rect 233716 407260 233726 407316
rect 342738 407260 342748 407316
rect 342804 407260 367276 407316
rect 367332 407260 367342 407316
rect 192546 407148 192556 407204
rect 192612 407148 197484 407204
rect 197540 407148 197550 407204
rect 203186 407148 203196 407204
rect 203252 407148 253708 407204
rect 253764 407148 253774 407204
rect 299170 407148 299180 407204
rect 299236 407148 521500 407204
rect 521556 407148 521566 407204
rect 153682 407036 153692 407092
rect 153748 407036 289884 407092
rect 289940 407036 289950 407092
rect 338706 407036 338716 407092
rect 338772 407036 388444 407092
rect 388500 407036 388510 407092
rect 390562 407036 390572 407092
rect 390628 407036 432796 407092
rect 432852 407036 432862 407092
rect 339154 406924 339164 406980
rect 339220 406924 410620 406980
rect 410676 406924 410686 406980
rect 338034 406812 338044 406868
rect 338100 406812 506716 406868
rect 506772 406812 506782 406868
rect 196018 406700 196028 406756
rect 196084 406700 199052 406756
rect 199108 406700 199118 406756
rect 252802 406700 252812 406756
rect 252868 406700 337708 406756
rect 352118 406700 352156 406756
rect 352212 406700 352222 406756
rect 354722 406700 354732 406756
rect 354788 406700 366268 406756
rect 366324 406700 366334 406756
rect 383058 406700 383068 406756
rect 383124 406700 573244 406756
rect 573300 406700 573310 406756
rect 337652 406644 337708 406700
rect 163090 406588 163100 406644
rect 163156 406588 163660 406644
rect 163716 406588 216636 406644
rect 216692 406588 218204 406644
rect 218260 406588 218270 406644
rect 305778 406588 305788 406644
rect 305844 406588 306796 406644
rect 306852 406588 306862 406644
rect 337652 406588 352828 406644
rect 352884 406588 352894 406644
rect 372726 406588 372764 406644
rect 372820 406588 372830 406644
rect 434550 406588 434588 406644
rect 434644 406588 434654 406644
rect 499286 406588 499324 406644
rect 499380 406588 499390 406644
rect 501526 406588 501564 406644
rect 501620 406588 501630 406644
rect 511830 406588 511868 406644
rect 511924 406588 511934 406644
rect 514098 406588 514108 406644
rect 514164 406588 514202 406644
rect 516982 406588 517020 406644
rect 517076 406588 517086 406644
rect 522134 406588 522172 406644
rect 522228 406588 522238 406644
rect 528854 406588 528892 406644
rect 528948 406588 528958 406644
rect 543638 406588 543676 406644
rect 543732 406588 543742 406644
rect 551030 406588 551068 406644
rect 551124 406588 551134 406644
rect 558198 406588 558236 406644
rect 558292 406588 558302 406644
rect 580598 406588 580636 406644
rect 580692 406588 580702 406644
rect 196466 406476 196476 406532
rect 196532 406476 243964 406532
rect 244020 406476 246876 406532
rect 246932 406476 246942 406532
rect 357858 406476 357868 406532
rect 357924 406476 362796 406532
rect 362852 406476 362862 406532
rect 374658 406476 374668 406532
rect 374724 406476 383292 406532
rect 383348 406476 383358 406532
rect 354610 406364 354620 406420
rect 354676 406364 383068 406420
rect 383124 406364 383134 406420
rect 392242 406364 392252 406420
rect 392308 406364 440188 406420
rect 440244 406364 440254 406420
rect 337026 406252 337036 406308
rect 337092 406252 403900 406308
rect 403956 406252 403966 406308
rect 83944 406140 163660 406196
rect 163716 406140 163726 406196
rect 213042 406140 213052 406196
rect 213108 406140 340956 406196
rect 341012 406140 341022 406196
rect 403218 406140 403228 406196
rect 403284 406140 475804 406196
rect 475860 406140 475870 406196
rect 338594 406028 338604 406084
rect 338660 406028 486108 406084
rect 486164 406028 486174 406084
rect 338818 405916 338828 405972
rect 338884 405916 506156 405972
rect 506212 405916 506222 405972
rect 202738 405804 202748 405860
rect 202804 405804 213052 405860
rect 213108 405804 213118 405860
rect 339826 405804 339836 405860
rect 339892 405804 527324 405860
rect 527380 405804 527390 405860
rect 189634 405692 189644 405748
rect 189700 405692 203084 405748
rect 203140 405692 203150 405748
rect 271618 405692 271628 405748
rect 271684 405692 491260 405748
rect 491316 405692 491326 405748
rect 371298 405580 371308 405636
rect 371364 405580 455196 405636
rect 455252 405580 455262 405636
rect 347890 405356 347900 405412
rect 347956 405356 354732 405412
rect 354788 405356 354798 405412
rect 357270 405356 357308 405412
rect 357364 405356 357374 405412
rect 272962 405244 272972 405300
rect 273028 405244 347788 405300
rect 347844 405244 347854 405300
rect 354498 405244 354508 405300
rect 354564 405244 393148 405300
rect 393204 405244 393214 405300
rect 340610 405132 340620 405188
rect 340676 405132 350308 405188
rect 354498 405132 354508 405188
rect 354564 405132 367948 405188
rect 368004 405132 368014 405188
rect 350252 405076 350308 405132
rect 162978 405020 162988 405076
rect 163044 405020 163660 405076
rect 163716 405020 202748 405076
rect 202804 405020 202814 405076
rect 296482 405020 296492 405076
rect 296548 405020 347564 405076
rect 347620 405020 347630 405076
rect 350252 405020 356188 405076
rect 356244 405020 356254 405076
rect 398150 405020 398188 405076
rect 398244 405020 398254 405076
rect 202402 404908 202412 404964
rect 202468 404908 268716 404964
rect 268772 404908 268782 404964
rect 340162 404908 340172 404964
rect 340228 404908 350588 404964
rect 350644 404908 350654 404964
rect 350914 404908 350924 404964
rect 350980 404908 356188 404964
rect 356132 404852 356188 404908
rect 361172 404908 365092 404964
rect 367574 404908 367612 404964
rect 367668 404908 367678 404964
rect 367798 404908 367836 404964
rect 367892 404908 367902 404964
rect 391458 404908 391468 404964
rect 391524 404908 403900 404964
rect 403956 404908 403966 404964
rect 361172 404852 361228 404908
rect 365036 404852 365092 404908
rect 199602 404796 199612 404852
rect 199668 404796 264236 404852
rect 264292 404796 264302 404852
rect 342486 404796 342524 404852
rect 342580 404796 342590 404852
rect 342738 404796 342748 404852
rect 342804 404796 346332 404852
rect 346388 404796 346398 404852
rect 347554 404796 347564 404852
rect 347620 404796 350700 404852
rect 350756 404796 350766 404852
rect 356132 404796 361228 404852
rect 362898 404796 362908 404852
rect 362964 404796 364812 404852
rect 364868 404796 364878 404852
rect 365036 404796 527436 404852
rect 527492 404796 527502 404852
rect 192770 404684 192780 404740
rect 192836 404684 252140 404740
rect 252196 404684 252206 404740
rect 255490 404684 255500 404740
rect 255556 404684 429436 404740
rect 429492 404684 429502 404740
rect 439030 404684 439068 404740
rect 439124 404684 439134 404740
rect 196130 404572 196140 404628
rect 196196 404572 256172 404628
rect 256228 404572 256238 404628
rect 259522 404572 259532 404628
rect 259588 404572 444892 404628
rect 444948 404572 444958 404628
rect 186162 404460 186172 404516
rect 186228 404460 202412 404516
rect 202468 404460 202478 404516
rect 242050 404460 242060 404516
rect 242116 404460 377916 404516
rect 377972 404460 377982 404516
rect 383170 404460 383180 404516
rect 383236 404460 389676 404516
rect 389732 404460 389742 404516
rect 389890 404460 389900 404516
rect 389956 404460 398300 404516
rect 398356 404460 398366 404516
rect 403890 404460 403900 404516
rect 403956 404460 590716 404516
rect 590772 404460 590782 404516
rect 197698 404348 197708 404404
rect 197764 404348 269612 404404
rect 269668 404348 269678 404404
rect 285058 404348 285068 404404
rect 285124 404348 344428 404404
rect 350802 404348 350812 404404
rect 350868 404348 354508 404404
rect 354564 404348 354574 404404
rect 354722 404348 354732 404404
rect 354788 404348 354798 404404
rect 361442 404348 361452 404404
rect 361508 404348 363020 404404
rect 363076 404348 363086 404404
rect 364662 404348 364700 404404
rect 364756 404348 364766 404404
rect 366146 404348 366156 404404
rect 366212 404348 384748 404404
rect 390534 404348 390572 404404
rect 390628 404348 390638 404404
rect 395798 404348 395836 404404
rect 395892 404348 395902 404404
rect 398402 404348 398412 404404
rect 398468 404348 398506 404404
rect 398626 404348 398636 404404
rect 398692 404348 404012 404404
rect 404068 404348 404078 404404
rect 408212 404348 536284 404404
rect 536340 404348 536350 404404
rect 202514 404236 202524 404292
rect 202580 404236 274988 404292
rect 275044 404236 275054 404292
rect 344372 404180 344428 404348
rect 351446 404236 351484 404292
rect 351540 404236 351550 404292
rect 354732 404180 354788 404348
rect 384692 404292 384748 404348
rect 408212 404292 408268 404348
rect 357858 404236 357868 404292
rect 357924 404236 367836 404292
rect 367892 404236 367902 404292
rect 373622 404236 373660 404292
rect 373716 404236 373726 404292
rect 384692 404236 408268 404292
rect 447542 404236 447580 404292
rect 447636 404236 447646 404292
rect 454934 404236 454972 404292
rect 455028 404236 455038 404292
rect 565814 404236 565852 404292
rect 565908 404236 565918 404292
rect 168802 404124 168812 404180
rect 168868 404124 197596 404180
rect 197652 404124 197662 404180
rect 199490 404124 199500 404180
rect 199556 404124 273644 404180
rect 273700 404124 273710 404180
rect 293794 404124 293804 404180
rect 293860 404124 339388 404180
rect 339444 404124 339454 404180
rect 344372 404124 354788 404180
rect 389442 404124 389452 404180
rect 389508 404124 398412 404180
rect 398468 404124 398478 404180
rect 196242 404012 196252 404068
rect 196308 404012 262892 404068
rect 262948 404012 262958 404068
rect 267586 404012 267596 404068
rect 267652 404012 342524 404068
rect 342580 404012 342590 404068
rect 374546 404012 374556 404068
rect 374612 404012 590492 404068
rect 590548 404012 590558 404068
rect -960 403732 480 403928
rect 191314 403900 191324 403956
rect 191380 403900 244076 403956
rect 244132 403900 244142 403956
rect 346882 403900 346892 403956
rect 346948 403900 439068 403956
rect 439124 403900 439134 403956
rect 189746 403788 189756 403844
rect 189812 403788 204428 403844
rect 204484 403788 204494 403844
rect 338818 403788 338828 403844
rect 338884 403788 347172 403844
rect 347116 403732 347172 403788
rect 352772 403788 367612 403844
rect 367668 403788 367678 403844
rect 591154 403788 591164 403844
rect 591220 403816 595672 403844
rect 591220 403788 597000 403816
rect 352772 403732 352828 403788
rect -960 403704 59612 403732
rect 392 403676 59612 403704
rect 59668 403676 59678 403732
rect 339266 403676 339276 403732
rect 339332 403676 346892 403732
rect 346948 403676 346958 403732
rect 347116 403676 352828 403732
rect 364690 403676 364700 403732
rect 364756 403676 390572 403732
rect 390628 403676 390638 403732
rect 398178 403676 398188 403732
rect 398244 403676 447580 403732
rect 447636 403676 447646 403732
rect 356178 403564 356188 403620
rect 356244 403564 389788 403620
rect 389844 403564 389854 403620
rect 595560 403592 597000 403788
rect 339042 403452 339052 403508
rect 339108 403452 352716 403508
rect 352772 403452 352782 403508
rect 359762 403452 359772 403508
rect 359828 403452 374556 403508
rect 374612 403452 374622 403508
rect 350466 403340 350476 403396
rect 350532 403340 359996 403396
rect 360052 403340 360062 403396
rect 83944 403228 93324 403284
rect 93380 403228 93390 403284
rect 340386 403228 340396 403284
rect 340452 403228 361228 403284
rect 351026 403116 351036 403172
rect 351092 403116 357868 403172
rect 357924 403116 357934 403172
rect 361172 403116 361228 403228
rect 361284 403116 361294 403172
rect 384850 403116 384860 403172
rect 384916 403116 389900 403172
rect 389956 403116 389966 403172
rect 393474 403116 393484 403172
rect 393540 403116 403228 403172
rect 403284 403116 403294 403172
rect 347778 403004 347788 403060
rect 347844 403004 356636 403060
rect 356692 403004 356702 403060
rect 363010 403004 363020 403060
rect 363076 403004 374668 403060
rect 374724 403004 374734 403060
rect 383058 403004 383068 403060
rect 383124 403004 391468 403060
rect 391524 403004 391534 403060
rect 393138 403004 393148 403060
rect 393204 403004 454972 403060
rect 455028 403004 455038 403060
rect 187954 402892 187964 402948
rect 188020 402892 250796 402948
rect 250852 402892 250862 402948
rect 291106 402892 291116 402948
rect 291172 402892 342748 402948
rect 342804 402892 342814 402948
rect 359874 402892 359884 402948
rect 359940 402892 373660 402948
rect 373716 402892 373726 402948
rect 389666 402892 389676 402948
rect 389732 402892 434588 402948
rect 434644 402892 434654 402948
rect 184706 402780 184716 402836
rect 184772 402780 248108 402836
rect 248164 402780 248174 402836
rect 341170 402780 341180 402836
rect 341236 402780 395836 402836
rect 395892 402780 395902 402836
rect 189298 402668 189308 402724
rect 189364 402668 260204 402724
rect 260260 402668 260270 402724
rect 284386 402668 284396 402724
rect 284452 402668 342636 402724
rect 342692 402668 342702 402724
rect 367826 402668 367836 402724
rect 367892 402668 383180 402724
rect 383236 402668 383246 402724
rect 389778 402668 389788 402724
rect 389844 402668 501564 402724
rect 501620 402668 501630 402724
rect 189298 402556 189308 402612
rect 189364 402556 281708 402612
rect 281764 402556 281774 402612
rect 283714 402556 283724 402612
rect 283780 402556 351484 402612
rect 351540 402556 351550 402612
rect 366146 402556 366156 402612
rect 366212 402556 389452 402612
rect 389508 402556 389518 402612
rect 187730 402444 187740 402500
rect 187796 402444 246764 402500
rect 246820 402444 246830 402500
rect 247426 402444 247436 402500
rect 247492 402444 350588 402500
rect 350644 402444 350654 402500
rect 240706 402332 240716 402388
rect 240772 402332 372764 402388
rect 372820 402332 372830 402388
rect 527426 402332 527436 402388
rect 527492 402332 585452 402388
rect 585508 402332 585518 402388
rect 337652 402220 340172 402276
rect 340228 402220 340238 402276
rect 336130 402108 336140 402164
rect 336196 402108 337596 402164
rect 337652 402108 337708 402220
rect 197586 401548 197596 401604
rect 197652 401548 336140 401604
rect 336196 401548 336206 401604
rect 189074 401100 189084 401156
rect 189140 401100 241388 401156
rect 241444 401100 241454 401156
rect 196354 400988 196364 401044
rect 196420 400988 249452 401044
rect 249508 400988 249518 401044
rect 189186 400876 189196 400932
rect 189252 400876 257516 400932
rect 257572 400876 257582 400932
rect 192882 400764 192892 400820
rect 192948 400764 265580 400820
rect 265636 400764 265646 400820
rect 187842 400652 187852 400708
rect 187908 400652 201404 400708
rect 201460 400652 201470 400708
rect 202626 400652 202636 400708
rect 202692 400652 277676 400708
rect 277732 400652 277742 400708
rect 83944 400316 88172 400372
rect 88228 400316 88238 400372
rect 201394 399868 201404 399924
rect 201460 399868 329644 399924
rect 329700 399868 329710 399924
rect 299842 399644 299852 399700
rect 299908 399644 339612 399700
rect 339668 399644 339678 399700
rect 297826 399532 297836 399588
rect 297892 399532 338044 399588
rect 338100 399532 338110 399588
rect 189410 399420 189420 399476
rect 189476 399420 258860 399476
rect 258916 399420 258926 399476
rect 289090 399420 289100 399476
rect 289156 399420 339164 399476
rect 339220 399420 339230 399476
rect 197810 399308 197820 399364
rect 197876 399308 270956 399364
rect 271012 399308 271022 399364
rect 337586 399308 337596 399364
rect 337652 399308 340088 399364
rect 189410 399196 189420 399252
rect 189476 399196 280364 399252
rect 280420 399196 280430 399252
rect 285730 399196 285740 399252
rect 285796 399196 338604 399252
rect 338660 399196 338670 399252
rect 187618 399084 187628 399140
rect 187684 399084 199276 399140
rect 199332 399084 199342 399140
rect 244738 399084 244748 399140
rect 244804 399084 338940 399140
rect 338996 399084 339006 399140
rect 184594 398972 184604 399028
rect 184660 398972 333564 399028
rect 333620 398972 333630 399028
rect 199266 398188 199276 398244
rect 199332 398188 330988 398244
rect 331044 398188 331054 398244
rect 197474 398076 197484 398132
rect 197540 398076 200508 398132
rect 200564 398076 200574 398132
rect 200946 398076 200956 398132
rect 201012 398076 202860 398132
rect 202916 398076 202926 398132
rect 204754 398076 204764 398132
rect 204820 398076 204988 398132
rect 205044 398076 228508 398132
rect 228564 398076 228574 398132
rect 188066 397964 188076 398020
rect 188132 397964 240044 398020
rect 240100 397964 240110 398020
rect 192994 397852 193004 397908
rect 193060 397852 245420 397908
rect 245476 397852 245486 397908
rect 199042 397740 199052 397796
rect 199108 397740 202636 397796
rect 202692 397740 202702 397796
rect 202850 397740 202860 397796
rect 202916 397740 272300 397796
rect 272356 397740 272366 397796
rect 201282 397628 201292 397684
rect 201348 397628 276332 397684
rect 276388 397628 276398 397684
rect 167122 397516 167132 397572
rect 167188 397516 192444 397572
rect 192500 397516 192510 397572
rect 203522 397516 203532 397572
rect 203588 397516 279020 397572
rect 279076 397516 279086 397572
rect 279682 397516 279692 397572
rect 279748 397516 339500 397572
rect 339556 397516 339566 397572
rect 83944 397404 93212 397460
rect 93268 397404 93278 397460
rect 94882 397404 94892 397460
rect 94948 397404 209132 397460
rect 209188 397404 209198 397460
rect 274306 397404 274316 397460
rect 274372 397404 340620 397460
rect 340676 397404 340686 397460
rect 85250 397292 85260 397348
rect 85316 397292 315308 397348
rect 315364 397292 315374 397348
rect 177202 397180 177212 397236
rect 177268 397180 205212 397236
rect 205268 397180 205278 397236
rect 198034 396396 198044 396452
rect 198100 396396 223356 396452
rect 223412 396396 223422 396452
rect 290434 396396 290444 396452
rect 290500 396396 340284 396452
rect 340340 396396 340350 396452
rect 287746 396284 287756 396340
rect 287812 396284 337708 396340
rect 337764 396284 337774 396340
rect 283042 396172 283052 396228
rect 283108 396172 340060 396228
rect 340116 396172 340126 396228
rect 281026 396060 281036 396116
rect 281092 396060 339836 396116
rect 339892 396060 339902 396116
rect 184594 395948 184604 396004
rect 184660 395948 194908 396004
rect 194964 395948 194974 396004
rect 197922 395948 197932 396004
rect 197988 395948 266924 396004
rect 266980 395948 266990 396004
rect 275650 395948 275660 396004
rect 275716 395948 338828 396004
rect 338884 395948 338894 396004
rect 165554 395836 165564 395892
rect 165620 395836 198044 395892
rect 198100 395836 198110 395892
rect 250114 395836 250124 395892
rect 250180 395836 340508 395892
rect 340564 395836 340574 395892
rect 152002 395724 152012 395780
rect 152068 395724 205772 395780
rect 205828 395724 205838 395780
rect 223346 395724 223356 395780
rect 223412 395724 330316 395780
rect 330372 395724 330382 395780
rect 196354 395612 196364 395668
rect 196420 395612 340620 395668
rect 340676 395612 340686 395668
rect 194898 394828 194908 394884
rect 194964 394828 196252 394884
rect 196308 394828 333116 394884
rect 333172 394828 333182 394884
rect 585442 394828 585452 394884
rect 585508 394828 590604 394884
rect 590660 394828 590670 394884
rect 186274 394604 186284 394660
rect 186340 394604 201068 394660
rect 201124 394604 201134 394660
rect 83944 394492 277228 394548
rect 277284 394492 277294 394548
rect 186386 394380 186396 394436
rect 186452 394380 201740 394436
rect 201796 394380 201806 394436
rect 202514 394380 202524 394436
rect 202580 394380 229404 394436
rect 229460 394380 229470 394436
rect 160402 394268 160412 394324
rect 160468 394268 206444 394324
rect 206500 394268 206510 394324
rect 289874 394268 289884 394324
rect 289940 394268 335356 394324
rect 335412 394268 335422 394324
rect 186274 394156 186284 394212
rect 186340 394156 333452 394212
rect 333508 394156 333518 394212
rect 88274 394044 88284 394100
rect 88340 394044 313964 394100
rect 314020 394044 314030 394100
rect 85026 393932 85036 393988
rect 85092 393932 317324 393988
rect 317380 393932 317390 393988
rect 192434 393260 192444 393316
rect 192500 393260 334460 393316
rect 334516 393260 334526 393316
rect 187170 393148 187180 393204
rect 187236 393148 334348 393204
rect 334404 393148 334414 393204
rect 292450 392924 292460 392980
rect 292516 392924 339948 392980
rect 340004 392924 340014 392980
rect 295138 392812 295148 392868
rect 295204 392812 336924 392868
rect 336980 392812 336990 392868
rect 337138 392812 337148 392868
rect 337204 392812 337484 392868
rect 337540 392812 340088 392868
rect 258178 392700 258188 392756
rect 258244 392700 339276 392756
rect 339332 392700 339342 392756
rect 192322 392588 192332 392644
rect 192388 392588 227612 392644
rect 227668 392588 227678 392644
rect 256834 392588 256844 392644
rect 256900 392588 340396 392644
rect 340452 392588 340462 392644
rect 184482 392476 184492 392532
rect 184548 392476 191548 392532
rect 191604 392476 191614 392532
rect 193106 392476 193116 392532
rect 193172 392476 229628 392532
rect 229684 392476 229694 392532
rect 248770 392476 248780 392532
rect 248836 392476 339052 392532
rect 339108 392476 339118 392532
rect 90066 392364 90076 392420
rect 90132 392364 315980 392420
rect 316036 392364 316046 392420
rect 86818 392252 86828 392308
rect 86884 392252 314636 392308
rect 314692 392252 314702 392308
rect 83346 391804 83356 391860
rect 83412 391804 309260 391860
rect 309316 391804 309326 391860
rect 196466 391692 196476 391748
rect 196532 391692 336700 391748
rect 336756 391692 336766 391748
rect 83944 391580 86604 391636
rect 86660 391580 86670 391636
rect 89842 391580 89852 391636
rect 89908 391580 237356 391636
rect 237412 391580 237422 391636
rect 336690 391468 336700 391524
rect 336756 391468 337372 391524
rect 337428 391468 337438 391524
rect 186386 390908 186396 390964
rect 186452 390908 199612 390964
rect 199668 390908 199678 390964
rect 183026 390796 183036 390852
rect 183092 390796 201068 390852
rect 201124 390796 201134 390852
rect 277330 390796 277340 390852
rect 277396 390796 278012 390852
rect 278068 390796 278078 390852
rect 191426 390684 191436 390740
rect 191492 390684 229852 390740
rect 229908 390684 229918 390740
rect 299954 390684 299964 390740
rect 300020 390684 335468 390740
rect 335524 390684 335534 390740
rect 52882 390572 52892 390628
rect 52948 390572 207116 390628
rect 207172 390572 207182 390628
rect 284722 390572 284732 390628
rect 284788 390572 335244 390628
rect 335300 390572 335310 390628
rect 201282 390460 201292 390516
rect 201348 390460 277340 390516
rect 277396 390460 277406 390516
rect 595560 390404 597000 390600
rect 4162 390348 4172 390404
rect 4228 390348 199500 390404
rect 199556 390348 321692 390404
rect 321748 390348 321758 390404
rect 590482 390348 590492 390404
rect 590548 390376 597000 390404
rect 590548 390348 595672 390376
rect 199378 390236 199388 390292
rect 199444 390236 330316 390292
rect 330372 390236 330382 390292
rect 99922 390124 99932 390180
rect 99988 390124 236684 390180
rect 236740 390124 236750 390180
rect 37986 390012 37996 390068
rect 38052 390012 219884 390068
rect 219940 390012 219950 390068
rect 192546 389900 192556 389956
rect 192612 389900 330204 389956
rect 330260 389900 330270 389956
rect -960 389620 480 389816
rect 53106 389788 53116 389844
rect 53172 389788 305228 389844
rect 305284 389788 305294 389844
rect -960 389592 4284 389620
rect 392 389564 4284 389592
rect 4340 389564 4350 389620
rect 295810 389228 295820 389284
rect 295876 389228 337036 389284
rect 337092 389228 337102 389284
rect 288418 389116 288428 389172
rect 288484 389116 338492 389172
rect 338548 389116 338558 389172
rect 200498 389004 200508 389060
rect 200564 389004 217532 389060
rect 217588 389004 217598 389060
rect 287074 389004 287084 389060
rect 287140 389004 338716 389060
rect 338772 389004 338782 389060
rect 182242 388892 182252 388948
rect 182308 388892 316652 388948
rect 316708 388892 316718 388948
rect 201170 388780 201180 388836
rect 201236 388780 329756 388836
rect 329812 388780 329822 388836
rect 95106 388668 95116 388724
rect 95172 388668 233996 388724
rect 234052 388668 234062 388724
rect 94882 388556 94892 388612
rect 94948 388556 235340 388612
rect 235396 388556 235406 388612
rect 91522 388444 91532 388500
rect 91588 388444 232652 388500
rect 232708 388444 232718 388500
rect 196018 388332 196028 388388
rect 196084 388332 337820 388388
rect 337876 388332 337886 388388
rect 69682 388220 69692 388276
rect 69748 388220 307916 388276
rect 307972 388220 307982 388276
rect 316082 388220 316092 388276
rect 316148 388220 317436 388276
rect 317492 388220 336812 388276
rect 336868 388220 336878 388276
rect 20850 388108 20860 388164
rect 20916 388108 331100 388164
rect 331156 388108 331166 388164
rect 197474 387996 197484 388052
rect 197540 387996 207452 388052
rect 207508 387996 207518 388052
rect 331510 387996 331548 388052
rect 331604 387996 332556 388052
rect 332612 387996 332622 388052
rect 202626 387212 202636 387268
rect 202692 387212 218204 387268
rect 218260 387212 218270 387268
rect 277218 387212 277228 387268
rect 277284 387212 311948 387268
rect 312004 387212 312014 387268
rect 178882 387100 178892 387156
rect 178948 387100 228620 387156
rect 228676 387100 228686 387156
rect 96562 386988 96572 387044
rect 96628 386988 229964 387044
rect 230020 386988 230030 387044
rect 177202 386876 177212 386932
rect 177268 386876 311276 386932
rect 311332 386876 311342 386932
rect 163762 386764 163772 386820
rect 163828 386764 197484 386820
rect 197540 386764 197932 386820
rect 197988 386764 197998 386820
rect 204530 386764 204540 386820
rect 204596 386764 339500 386820
rect 339556 386764 339566 386820
rect 95330 386652 95340 386708
rect 95396 386652 231980 386708
rect 232036 386652 232046 386708
rect 91522 386540 91532 386596
rect 91588 386540 230636 386596
rect 230692 386540 230702 386596
rect 73490 386428 73500 386484
rect 73556 386428 308588 386484
rect 308644 386428 308654 386484
rect 337026 386316 337036 386372
rect 337092 386316 337484 386372
rect 337540 386316 340088 386372
rect 294802 386092 294812 386148
rect 294868 386092 332108 386148
rect 332164 386092 332174 386148
rect 268706 385980 268716 386036
rect 268772 385980 330092 386036
rect 330148 385980 330158 386036
rect 183922 385868 183932 385924
rect 183988 385868 312620 385924
rect 312676 385868 312686 385924
rect 180562 385756 180572 385812
rect 180628 385756 317996 385812
rect 318052 385756 318062 385812
rect 86482 385644 86492 385700
rect 86548 385644 318668 385700
rect 318724 385644 318734 385700
rect 84802 385532 84812 385588
rect 84868 385532 319340 385588
rect 319396 385532 319406 385588
rect 204418 385196 204428 385252
rect 204484 385196 326396 385252
rect 326452 385196 327404 385252
rect 327460 385196 327470 385252
rect 103282 385084 103292 385140
rect 103348 385084 234668 385140
rect 234724 385084 234734 385140
rect 91746 384972 91756 385028
rect 91812 384972 229292 385028
rect 229348 384972 229358 385028
rect 38434 384860 38444 384916
rect 38500 384860 219212 384916
rect 219268 384860 219278 384916
rect 40226 384748 40236 384804
rect 40292 384748 225932 384804
rect 225988 384748 225998 384804
rect 217522 384636 217532 384692
rect 217588 384636 225148 384692
rect 225204 384636 225214 384692
rect 208226 384188 208236 384244
rect 208292 384188 208348 384244
rect 208404 384188 208414 384244
rect 24322 384076 24332 384132
rect 24388 384076 212492 384132
rect 212548 384076 212558 384132
rect 34402 383964 34412 384020
rect 34468 383964 211820 384020
rect 211876 383964 211886 384020
rect 227602 383964 227612 384020
rect 227668 383964 266252 384020
rect 266308 383964 266318 384020
rect 306786 383964 306796 384020
rect 306852 383964 335580 384020
rect 335636 383964 335646 384020
rect 59602 383852 59612 383908
rect 59668 383852 209804 383908
rect 209860 383852 209870 383908
rect 243394 383852 243404 383908
rect 243460 383852 336588 383908
rect 336644 383852 336654 383908
rect 199042 383740 199052 383796
rect 199108 383740 227276 383796
rect 227332 383740 227342 383796
rect 179106 383628 179116 383684
rect 179172 383628 227948 383684
rect 228004 383628 228014 383684
rect 113474 383516 113484 383572
rect 113540 383516 210476 383572
rect 210532 383516 210542 383572
rect 335906 383516 335916 383572
rect 335972 383516 336924 383572
rect 336980 383516 336990 383572
rect 176978 383404 176988 383460
rect 177044 383404 306572 383460
rect 306628 383404 306638 383460
rect 177426 383292 177436 383348
rect 177492 383292 307244 383348
rect 307300 383292 307310 383348
rect 197362 383180 197372 383236
rect 197428 383180 226604 383236
rect 226660 383180 226670 383236
rect 274642 383180 274652 383236
rect 274708 383180 335132 383236
rect 335188 383180 335198 383236
rect 208898 383068 208908 383124
rect 208964 383068 334908 383124
rect 334964 383068 334974 383124
rect 206658 382956 206668 383012
rect 206724 382956 207788 383012
rect 207844 382956 207854 383012
rect 229842 382956 229852 383012
rect 229908 382956 237692 383012
rect 237748 382956 237758 383012
rect 189522 382844 189532 382900
rect 189588 382844 199724 382900
rect 199780 382844 199790 382900
rect 229618 382844 229628 382900
rect 229684 382844 251468 382900
rect 251524 382844 251534 382900
rect 229394 382732 229404 382788
rect 229460 382732 254156 382788
rect 254212 382732 254222 382788
rect 202850 382620 202860 382676
rect 202916 382620 217868 382676
rect 217924 382620 217934 382676
rect 225138 382620 225148 382676
rect 225204 382620 268940 382676
rect 268996 382620 269006 382676
rect 218194 382508 218204 382564
rect 218260 382508 263564 382564
rect 263620 382508 263630 382564
rect 276994 382508 277004 382564
rect 277060 382508 339052 382564
rect 339108 382508 339118 382564
rect 201506 382396 201516 382452
rect 201572 382396 268268 382452
rect 268324 382396 268334 382452
rect 270274 382396 270284 382452
rect 270340 382396 338604 382452
rect 338660 382396 338670 382452
rect 198370 382284 198380 382340
rect 198436 382284 199836 382340
rect 199892 382284 199902 382340
rect 239362 382284 239372 382340
rect 239428 382284 338828 382340
rect 338884 382284 338894 382340
rect 197026 382172 197036 382228
rect 197092 382172 197708 382228
rect 197764 382172 197774 382228
rect 198118 382172 198156 382228
rect 198212 382172 198222 382228
rect 199042 382172 199052 382228
rect 199108 382172 199724 382228
rect 199780 382172 199790 382228
rect 199910 382172 199948 382228
rect 200004 382172 200014 382228
rect 204082 382172 204092 382228
rect 204148 382172 206556 382228
rect 206612 382172 331884 382228
rect 331940 382172 331950 382228
rect 111682 382060 111692 382116
rect 111748 382060 236012 382116
rect 236068 382060 236078 382116
rect 237682 382060 237692 382116
rect 237748 382060 246092 382116
rect 246148 382060 246158 382116
rect 301186 382060 301196 382116
rect 301252 382060 302316 382116
rect 302372 382060 302382 382116
rect 303202 382060 303212 382116
rect 303268 382060 303884 382116
rect 303940 382060 303950 382116
rect 160402 381948 160412 382004
rect 160468 381948 222572 382004
rect 222628 381948 222638 382004
rect 242722 381948 242732 382004
rect 242788 381948 243516 382004
rect 243572 381948 243582 382004
rect 262210 381948 262220 382004
rect 262276 381948 263676 382004
rect 263732 381948 263742 382004
rect 278758 381948 278796 382004
rect 278852 381948 278862 382004
rect 297154 381948 297164 382004
rect 297220 381948 297276 382004
rect 297332 381948 297342 382004
rect 298918 381948 298956 382004
rect 299012 381948 299022 382004
rect 300514 381948 300524 382004
rect 300580 381948 300636 382004
rect 300692 381948 300702 382004
rect 302166 381948 302204 382004
rect 302260 381948 302270 382004
rect 303874 381948 303884 382004
rect 303940 381948 303996 382004
rect 304052 381948 304062 382004
rect 313282 381948 313292 382004
rect 313348 381948 313404 382004
rect 313460 381948 313470 382004
rect 118402 381836 118412 381892
rect 118468 381836 221900 381892
rect 221956 381836 221966 381892
rect 116722 381724 116732 381780
rect 116788 381724 223916 381780
rect 223972 381724 223982 381780
rect 113362 381612 113372 381668
rect 113428 381612 220556 381668
rect 220612 381612 220622 381668
rect 260866 381612 260876 381668
rect 260932 381612 261996 381668
rect 262052 381612 262062 381668
rect 294466 381612 294476 381668
rect 294532 381612 295596 381668
rect 295652 381612 295662 381668
rect 304546 381612 304556 381668
rect 304612 381612 305676 381668
rect 305732 381612 305742 381668
rect 104962 381500 104972 381556
rect 105028 381500 225260 381556
rect 225316 381500 225326 381556
rect 214470 381388 214508 381444
rect 214564 381388 214574 381444
rect 216486 381388 216524 381444
rect 216580 381388 216590 381444
rect 293122 381388 293132 381444
rect 293188 381388 293916 381444
rect 293972 381388 293982 381444
rect 215012 380828 231868 380884
rect 321682 380828 321692 380884
rect 321748 380828 330652 380884
rect 330708 380828 330718 380884
rect 215012 380660 215068 380828
rect 231812 380660 231868 380828
rect 311602 380716 311612 380772
rect 311668 380716 330428 380772
rect 330484 380716 330494 380772
rect 197698 380604 197708 380660
rect 197764 380604 215068 380660
rect 216626 380604 216636 380660
rect 216692 380604 226828 380660
rect 231812 380604 274652 380660
rect 274708 380604 274718 380660
rect 278002 380604 278012 380660
rect 278068 380604 330204 380660
rect 330260 380604 330270 380660
rect 226772 380548 226828 380604
rect 189522 380492 189532 380548
rect 189588 380492 208908 380548
rect 208964 380492 208974 380548
rect 209122 380492 209132 380548
rect 209188 380492 223244 380548
rect 223300 380492 223310 380548
rect 226772 380492 328636 380548
rect 328692 380492 328702 380548
rect 162082 380380 162092 380436
rect 162148 380380 231308 380436
rect 231364 380380 231374 380436
rect 96786 380268 96796 380324
rect 96852 380268 233324 380324
rect 233380 380268 233390 380324
rect 38210 380156 38220 380212
rect 38276 380156 221228 380212
rect 221284 380156 221294 380212
rect 40114 380044 40124 380100
rect 40180 380044 209132 380100
rect 209188 380044 209198 380100
rect 215012 380044 224140 380100
rect 224196 380044 224206 380100
rect 215012 379988 215068 380044
rect 38322 379932 38332 379988
rect 38388 379932 215068 379988
rect 215814 379932 215852 379988
rect 215908 379932 215918 379988
rect 81106 379820 81116 379876
rect 81172 379820 309932 379876
rect 309988 379820 309998 379876
rect 336914 379820 336924 379876
rect 336980 379820 340088 379876
rect 58258 379708 58268 379764
rect 58324 379708 305900 379764
rect 305956 379708 305966 379764
rect 44482 379596 44492 379652
rect 44548 379596 211148 379652
rect 211204 379596 211214 379652
rect 218502 379596 218540 379652
rect 218596 379596 218606 379652
rect 328626 379596 328636 379652
rect 328692 379596 329084 379652
rect 329140 379596 338492 379652
rect 338548 379596 338558 379652
rect 190726 379484 190764 379540
rect 190820 379484 190830 379540
rect 191286 379484 191324 379540
rect 191380 379484 191390 379540
rect 192070 379484 192108 379540
rect 192164 379484 192174 379540
rect 192630 379484 192668 379540
rect 192724 379484 192734 379540
rect 193302 379484 193340 379540
rect 193396 379484 193406 379540
rect 194646 379484 194684 379540
rect 194740 379484 194750 379540
rect 195206 379484 195244 379540
rect 195300 379484 195310 379540
rect 196354 379484 196364 379540
rect 196420 379484 282380 379540
rect 282436 379484 282446 379540
rect 84914 379372 84924 379428
rect 84980 379372 310604 379428
rect 310660 379372 310670 379428
rect 192966 379260 193004 379316
rect 193060 379260 193070 379316
rect 195010 379260 195020 379316
rect 195076 379260 196140 379316
rect 196196 379260 196206 379316
rect 213126 379260 213164 379316
rect 213220 379260 213230 379316
rect 213798 379260 213836 379316
rect 213892 379260 213902 379316
rect 215142 379260 215180 379316
rect 215236 379260 215246 379316
rect 217158 379260 217196 379316
rect 217252 379260 217262 379316
rect 204306 378700 204316 378756
rect 204372 378700 330092 378756
rect 330148 378700 330158 378756
rect 587122 377356 587132 377412
rect 587188 377384 595672 377412
rect 587188 377356 597000 377384
rect 4274 377132 4284 377188
rect 4340 377132 165452 377188
rect 165508 377132 165518 377188
rect 595560 377160 597000 377356
rect 392 375704 4172 375732
rect -960 375676 4172 375704
rect 4228 375676 4238 375732
rect -960 375480 480 375676
rect 88162 374556 88172 374612
rect 88228 374556 88956 374612
rect 89012 374556 89022 374612
rect 171378 374556 171388 374612
rect 171444 374556 172172 374612
rect 172228 374556 172238 374612
rect 329896 373996 337820 374052
rect 337876 373996 337886 374052
rect 88946 373772 88956 373828
rect 89012 373772 171388 373828
rect 171444 373772 171454 373828
rect 337362 373324 337372 373380
rect 337428 373324 340088 373380
rect 329896 373100 330428 373156
rect 330484 373100 330494 373156
rect 329410 372204 329420 372260
rect 329476 372204 329486 372260
rect 329896 371308 340508 371364
rect 340564 371308 340574 371364
rect 329896 370412 333340 370468
rect 333396 370412 333406 370468
rect 329896 369516 337708 369572
rect 337764 369516 337774 369572
rect 177874 368620 177884 368676
rect 177940 368620 180040 368676
rect 329896 368620 340284 368676
rect 340340 368620 340350 368676
rect 329896 367724 339612 367780
rect 339668 367724 339678 367780
rect 177762 367500 177772 367556
rect 177828 367500 180040 367556
rect 93202 367052 93212 367108
rect 93268 367052 168028 367108
rect 168084 367052 168812 367108
rect 168868 367052 168878 367108
rect 177986 366380 177996 366436
rect 178052 366380 180040 366436
rect 329532 366324 329588 366856
rect 332546 366828 332556 366884
rect 332612 366828 340088 366884
rect 329522 366268 329532 366324
rect 329588 366268 329598 366324
rect 166338 366156 166348 366212
rect 166404 366156 167132 366212
rect 167188 366156 167198 366212
rect 329896 365932 340620 365988
rect 340676 365932 340686 365988
rect 86482 365372 86492 365428
rect 86548 365372 166348 365428
rect 166404 365372 166414 365428
rect 177650 365260 177660 365316
rect 177716 365260 180040 365316
rect 329896 365036 331212 365092
rect 331268 365036 331278 365092
rect 50642 364476 50652 364532
rect 50708 364476 53116 364532
rect 53172 364476 53182 364532
rect 77298 363916 77308 363972
rect 77364 363916 83356 363972
rect 83412 363916 83422 363972
rect 88722 363916 88732 363972
rect 88788 363916 177212 363972
rect 177268 363916 177278 363972
rect 65874 363804 65884 363860
rect 65940 363804 177436 363860
rect 177492 363804 177502 363860
rect 62066 363692 62076 363748
rect 62132 363692 176988 363748
rect 177044 363692 177054 363748
rect 180012 363300 180068 364168
rect 329896 364140 338044 364196
rect 338100 364140 338110 364196
rect 590594 364140 590604 364196
rect 590660 364168 595672 364196
rect 590660 364140 597000 364168
rect 595560 363944 597000 364140
rect 160860 363244 180068 363300
rect 160860 363048 160916 363244
rect 174738 363020 174748 363076
rect 174804 363020 180040 363076
rect 329420 362964 329476 363272
rect 54450 362908 54460 362964
rect 54516 362908 86492 362964
rect 86548 362908 86558 362964
rect 329410 362908 329420 362964
rect 329476 362908 329486 362964
rect 329896 362348 338044 362404
rect 338100 362348 338110 362404
rect 174850 361900 174860 361956
rect 174916 361900 180040 361956
rect -960 361396 480 361592
rect 329896 361452 331772 361508
rect 331828 361452 331838 361508
rect -960 361368 113484 361396
rect 392 361340 113484 361368
rect 113540 361340 113550 361396
rect 176194 360780 176204 360836
rect 176260 360780 180040 360836
rect 329896 360556 334572 360612
rect 334628 360556 334638 360612
rect 86482 360332 86492 360388
rect 86548 360332 89964 360388
rect 90020 360332 90030 360388
rect 336354 360332 336364 360388
rect 336420 360332 340088 360388
rect 88946 359884 88956 359940
rect 89012 359884 92428 359940
rect 92484 359884 92494 359940
rect 161252 359772 174748 359828
rect 174804 359772 174814 359828
rect 161252 359716 161308 359772
rect 160888 359660 161308 359716
rect 171378 359660 171388 359716
rect 171444 359660 180040 359716
rect 329896 359660 333228 359716
rect 333284 359660 333294 359716
rect 329896 358764 339500 358820
rect 339556 358764 339566 358820
rect 177202 358540 177212 358596
rect 177268 358540 180040 358596
rect 329896 357868 338492 357924
rect 338548 357868 338558 357924
rect 165666 357420 165676 357476
rect 165732 357420 180040 357476
rect 329896 356972 340172 357028
rect 340228 356972 340238 357028
rect 160888 356300 174860 356356
rect 174916 356300 174926 356356
rect 177202 356300 177212 356356
rect 177268 356300 180040 356356
rect 329896 356076 330988 356132
rect 331044 356076 331054 356132
rect 166226 355180 166236 355236
rect 166292 355180 180040 355236
rect 329896 355180 339836 355236
rect 339892 355180 339902 355236
rect 329896 354284 333452 354340
rect 333508 354284 333518 354340
rect 167794 354060 167804 354116
rect 167860 354060 180040 354116
rect 330642 353836 330652 353892
rect 330708 353836 340088 353892
rect 329868 353108 329924 353416
rect 161252 353052 176204 353108
rect 176260 353052 176270 353108
rect 329868 353052 340396 353108
rect 340452 353052 340462 353108
rect 161252 352996 161308 353052
rect 160888 352940 161308 352996
rect 171266 352940 171276 352996
rect 171332 352940 180040 352996
rect 329896 352492 337932 352548
rect 337988 352492 337998 352548
rect 180124 351316 180180 351848
rect 329896 351596 334460 351652
rect 334516 351596 334526 351652
rect 180114 351260 180124 351316
rect 180180 351260 180190 351316
rect 595560 350756 597000 350952
rect 176306 350700 176316 350756
rect 176372 350700 180040 350756
rect 329896 350700 338604 350756
rect 338660 350700 338670 350756
rect 590594 350700 590604 350756
rect 590660 350728 597000 350756
rect 590660 350700 595672 350728
rect 329896 349804 331996 349860
rect 332052 349804 332062 349860
rect 160888 349580 171388 349636
rect 171444 349580 171454 349636
rect 179442 349580 179452 349636
rect 179508 349580 180040 349636
rect 329896 348908 336028 348964
rect 336084 348908 336094 348964
rect 172722 348460 172732 348516
rect 172788 348460 180040 348516
rect 329896 348012 332220 348068
rect 332276 348012 332286 348068
rect -960 347284 480 347480
rect 167906 347340 167916 347396
rect 167972 347340 180040 347396
rect 336802 347340 336812 347396
rect 336868 347340 337484 347396
rect 337540 347340 340088 347396
rect -960 347256 4284 347284
rect 392 347228 4284 347256
rect 4340 347228 4350 347284
rect 329756 346612 329812 347144
rect 329746 346556 329756 346612
rect 329812 346556 329822 346612
rect 160888 346220 161308 346276
rect 161364 346220 163100 346276
rect 163156 346220 163166 346276
rect 169586 346220 169596 346276
rect 169652 346220 180040 346276
rect 329896 346220 333340 346276
rect 333396 346220 333406 346276
rect 329896 345324 338716 345380
rect 338772 345324 338782 345380
rect 167682 345100 167692 345156
rect 167748 345100 180040 345156
rect 329896 344428 333452 344484
rect 333508 344428 333518 344484
rect 171154 343980 171164 344036
rect 171220 343980 180040 344036
rect 329896 343532 332668 343588
rect 332724 343532 332734 343588
rect 160888 342860 162988 342916
rect 163044 342860 163054 342916
rect 169362 342860 169372 342916
rect 169428 342860 180040 342916
rect 329896 342636 334012 342692
rect 334068 342636 334078 342692
rect 169474 341740 169484 341796
rect 169540 341740 180040 341796
rect 329896 341740 333788 341796
rect 333844 341740 333854 341796
rect 163090 340956 163100 341012
rect 163156 340956 163772 341012
rect 163828 340956 163838 341012
rect 330418 340956 330428 341012
rect 330484 340956 336812 341012
rect 336868 340956 340116 341012
rect 329896 340844 333004 340900
rect 333060 340844 333070 340900
rect 340060 340872 340116 340956
rect 172386 340620 172396 340676
rect 172452 340620 180040 340676
rect 329896 339948 333900 340004
rect 333956 339948 333966 340004
rect 160748 339332 160804 339528
rect 170930 339500 170940 339556
rect 170996 339500 180040 339556
rect 161084 339388 163100 339444
rect 163156 339388 163166 339444
rect 161084 339332 161140 339388
rect 160748 339276 161140 339332
rect 329896 339052 333116 339108
rect 333172 339052 333182 339108
rect 163762 338492 163772 338548
rect 163828 338492 177212 338548
rect 177268 338492 177278 338548
rect 176194 338380 176204 338436
rect 176260 338380 180040 338436
rect 329896 338156 332332 338212
rect 332388 338156 332398 338212
rect 595560 337652 597000 337736
rect 590706 337596 590716 337652
rect 590772 337596 597000 337652
rect 595560 337512 597000 337596
rect 171042 337260 171052 337316
rect 171108 337260 180040 337316
rect 329896 337260 339724 337316
rect 339780 337260 339790 337316
rect 329896 336364 334684 336420
rect 334740 336364 334750 336420
rect 160888 336140 171388 336196
rect 171444 336140 171454 336196
rect 174514 336140 174524 336196
rect 174580 336140 180040 336196
rect 329896 335468 340620 335524
rect 340676 335468 340686 335524
rect 172274 335020 172284 335076
rect 172340 335020 180040 335076
rect 329896 334572 332108 334628
rect 332164 334572 332174 334628
rect 334562 334348 334572 334404
rect 334628 334348 334796 334404
rect 334852 334348 334862 334404
rect 335570 334348 335580 334404
rect 335636 334348 336924 334404
rect 336980 334348 340088 334404
rect 172610 333900 172620 333956
rect 172676 333900 180040 333956
rect 329522 333676 329532 333732
rect 329588 333676 329598 333732
rect 392 333368 4172 333396
rect -960 333340 4172 333368
rect 4228 333340 4238 333396
rect -960 333144 480 333340
rect 160888 332780 168028 332836
rect 168084 332780 168094 332836
rect 174626 332780 174636 332836
rect 174692 332780 180040 332836
rect 329896 332780 334572 332836
rect 334628 332780 334638 332836
rect 329746 331884 329756 331940
rect 329812 331884 329822 331940
rect 179330 331660 179340 331716
rect 179396 331660 180040 331716
rect 329896 330988 331100 331044
rect 331156 330988 331166 331044
rect 89954 330876 89964 330932
rect 90020 330876 92540 330932
rect 92596 330876 92606 330932
rect 170818 330540 170828 330596
rect 170884 330540 180040 330596
rect 329896 330092 337932 330148
rect 337988 330092 337998 330148
rect 160888 329420 166348 329476
rect 166404 329420 166414 329476
rect 172498 329420 172508 329476
rect 172564 329420 180040 329476
rect 329746 329196 329756 329252
rect 329812 329196 329822 329252
rect 166114 328300 166124 328356
rect 166180 328300 180040 328356
rect 329896 328300 334460 328356
rect 334516 328300 334526 328356
rect 340060 327684 340116 327880
rect 335458 327628 335468 327684
rect 335524 327628 336812 327684
rect 336868 327628 340116 327684
rect 329896 327404 338604 327460
rect 338660 327404 338670 327460
rect 167570 327180 167580 327236
rect 167636 327180 180040 327236
rect 329298 326508 329308 326564
rect 329364 326508 329374 326564
rect 160888 326060 163772 326116
rect 163828 326060 163838 326116
rect 174402 326060 174412 326116
rect 174468 326060 180040 326116
rect 329896 325612 338492 325668
rect 338548 325612 338558 325668
rect 166002 324940 166012 324996
rect 166068 324940 180040 324996
rect 329896 324716 338716 324772
rect 338772 324716 338782 324772
rect 590482 324492 590492 324548
rect 590548 324520 595672 324548
rect 590548 324492 597000 324520
rect 595560 324296 597000 324492
rect 169250 323820 169260 323876
rect 169316 323820 180040 323876
rect 329298 323820 329308 323876
rect 329364 323820 329374 323876
rect 160300 323372 165564 323428
rect 165620 323372 165630 323428
rect 160300 322084 160356 323372
rect 329896 322924 335580 322980
rect 335636 322924 335646 322980
rect 174290 322700 174300 322756
rect 174356 322700 180040 322756
rect 149492 322028 160356 322084
rect 329896 322028 332332 322084
rect 332388 322028 332398 322084
rect 149492 321748 149548 322028
rect 106642 321692 106652 321748
rect 106708 321692 149548 321748
rect 176082 321580 176092 321636
rect 176148 321580 180040 321636
rect 332098 321356 332108 321412
rect 332164 321356 340088 321412
rect 329298 321132 329308 321188
rect 329364 321132 329374 321188
rect 93314 320796 93324 320852
rect 93380 320796 163100 320852
rect 163156 320796 163166 320852
rect 169586 320460 169596 320516
rect 169652 320460 180040 320516
rect 329896 320236 331996 320292
rect 332052 320236 332062 320292
rect 147746 320012 147756 320068
rect 147812 320012 177212 320068
rect 177268 320012 177278 320068
rect 177090 319340 177100 319396
rect 177156 319340 180040 319396
rect 329896 319340 334684 319396
rect 334740 319340 334750 319396
rect -960 319060 480 319256
rect 330306 319116 330316 319172
rect 330372 319116 334124 319172
rect 334180 319116 334190 319172
rect -960 319032 44492 319060
rect 392 319004 44492 319032
rect 44548 319004 44558 319060
rect 329896 318444 334460 318500
rect 334516 318444 334526 318500
rect 160514 318220 160524 318276
rect 160580 318220 180040 318276
rect 329896 317548 336476 317604
rect 336532 317548 336542 317604
rect 179554 317100 179564 317156
rect 179620 317100 180040 317156
rect 332546 316988 332556 317044
rect 332612 316988 333340 317044
rect 333396 316988 333406 317044
rect 329868 316036 329924 316680
rect 180114 315980 180124 316036
rect 180180 315980 180190 316036
rect 329868 315980 332556 316036
rect 332612 315980 332622 316036
rect 329896 315756 333788 315812
rect 333844 315756 333854 315812
rect 335346 315756 335356 315812
rect 335412 315756 336364 315812
rect 336420 315756 336430 315812
rect 177538 314860 177548 314916
rect 177604 314860 180040 314916
rect 329896 314860 334796 314916
rect 334852 314860 334862 314916
rect 336354 314860 336364 314916
rect 336420 314860 340088 314916
rect 329298 313964 329308 314020
rect 329364 313964 329374 314020
rect 176194 313740 176204 313796
rect 176260 313740 180040 313796
rect 4274 313292 4284 313348
rect 4340 313292 160412 313348
rect 160468 313292 160478 313348
rect 329298 313068 329308 313124
rect 329364 313068 329374 313124
rect 177874 312620 177884 312676
rect 177940 312620 180040 312676
rect 329896 312172 340172 312228
rect 340228 312172 340238 312228
rect 169474 311500 169484 311556
rect 169540 311500 180040 311556
rect 329896 311276 338156 311332
rect 338212 311276 338222 311332
rect 595560 311108 597000 311304
rect 590706 311052 590716 311108
rect 590772 311080 597000 311108
rect 590772 311052 595672 311080
rect 174514 310380 174524 310436
rect 174580 310380 180040 310436
rect 329896 310380 340284 310436
rect 340340 310380 340350 310436
rect 329896 309484 339388 309540
rect 339444 309484 339454 309540
rect 174290 309260 174300 309316
rect 174356 309260 180040 309316
rect 330530 309148 330540 309204
rect 330596 309148 331212 309204
rect 331268 309148 331278 309204
rect 329970 308924 329980 308980
rect 330036 308924 335020 308980
rect 335076 308924 335086 308980
rect 330194 308812 330204 308868
rect 330260 308812 332220 308868
rect 332276 308812 332286 308868
rect 329896 308588 333676 308644
rect 333732 308588 333742 308644
rect 329522 308364 329532 308420
rect 329588 308364 332108 308420
rect 332164 308364 332174 308420
rect 335234 308364 335244 308420
rect 335300 308364 337596 308420
rect 337652 308364 340088 308420
rect 330418 308252 330428 308308
rect 330484 308252 331100 308308
rect 331156 308252 331166 308308
rect 332658 308252 332668 308308
rect 332724 308252 333228 308308
rect 333284 308252 333294 308308
rect 171266 308140 171276 308196
rect 171332 308140 180040 308196
rect 330642 308140 330652 308196
rect 330708 308140 333340 308196
rect 333396 308140 333406 308196
rect 332770 308028 332780 308084
rect 332836 308028 333116 308084
rect 333172 308028 333182 308084
rect 329970 307916 329980 307972
rect 330036 307916 333228 307972
rect 333284 307916 333294 307972
rect 329896 307692 338044 307748
rect 338100 307692 338110 307748
rect 329746 307356 329756 307412
rect 329812 307356 334572 307412
rect 334628 307356 334638 307412
rect 180226 307020 180236 307076
rect 180292 307020 180302 307076
rect 329896 306796 334012 306852
rect 334068 306796 334078 306852
rect 179442 305900 179452 305956
rect 179508 305900 180040 305956
rect 329896 305900 335020 305956
rect 335076 305900 335086 305956
rect 332434 305676 332444 305732
rect 332500 305676 333788 305732
rect 333844 305676 333854 305732
rect 332322 305564 332332 305620
rect 332388 305564 333676 305620
rect 333732 305564 333742 305620
rect -960 304948 480 305144
rect 329896 305004 333116 305060
rect 333172 305004 333182 305060
rect -960 304920 155372 304948
rect 392 304892 155372 304920
rect 155428 304892 155438 304948
rect 167906 304780 167916 304836
rect 167972 304780 180040 304836
rect 333442 304444 333452 304500
rect 333508 304444 338828 304500
rect 338884 304444 338894 304500
rect 329896 304108 335468 304164
rect 335524 304108 335534 304164
rect 334786 303996 334796 304052
rect 334852 303996 335244 304052
rect 335300 303996 335310 304052
rect 334226 303884 334236 303940
rect 334292 303884 334796 303940
rect 334852 303884 334862 303940
rect 177762 303660 177772 303716
rect 177828 303660 180040 303716
rect 329896 303212 334348 303268
rect 334404 303212 334414 303268
rect 166226 302540 166236 302596
rect 166292 302540 180040 302596
rect 329896 302316 333228 302372
rect 333284 302316 333294 302372
rect 334002 302092 334012 302148
rect 334068 302092 336588 302148
rect 336644 302092 336654 302148
rect 330194 301868 330204 301924
rect 330260 301868 340088 301924
rect 172946 301420 172956 301476
rect 173012 301420 180040 301476
rect 329896 301420 331884 301476
rect 331940 301420 331950 301476
rect 333666 300860 333676 300916
rect 333732 300860 338100 300916
rect 337026 300748 337036 300804
rect 337092 300748 337820 300804
rect 337876 300748 337886 300804
rect 338044 300580 338100 300860
rect 329896 300524 331772 300580
rect 331828 300524 331838 300580
rect 337810 300524 337820 300580
rect 337876 300524 338100 300580
rect 174402 300300 174412 300356
rect 174468 300300 180040 300356
rect 329896 299628 331324 299684
rect 331380 299628 331390 299684
rect 330866 299292 330876 299348
rect 330932 299292 336476 299348
rect 336532 299292 336542 299348
rect 177202 299180 177212 299236
rect 177268 299180 180040 299236
rect 331538 299180 331548 299236
rect 331604 299180 332556 299236
rect 332612 299180 332622 299236
rect 332210 299068 332220 299124
rect 332276 299068 332668 299124
rect 332724 299068 332734 299124
rect 329896 298732 331212 298788
rect 331268 298732 331278 298788
rect 332546 298508 332556 298564
rect 332612 298508 335356 298564
rect 335412 298508 335422 298564
rect 177314 298060 177324 298116
rect 177380 298060 180040 298116
rect 595560 297892 597000 298088
rect 329858 297836 329868 297892
rect 329924 297836 329934 297892
rect 590818 297836 590828 297892
rect 590884 297864 597000 297892
rect 590884 297836 595672 297864
rect 331874 297500 331884 297556
rect 331940 297500 336700 297556
rect 336756 297500 336766 297556
rect 332406 297388 332444 297444
rect 332500 297388 332510 297444
rect 334674 297164 334684 297220
rect 334740 297164 335916 297220
rect 335972 297164 335982 297220
rect 177426 296940 177436 296996
rect 177492 296940 180040 296996
rect 329634 296940 329644 296996
rect 329700 296940 329710 296996
rect 10994 296492 11004 296548
rect 11060 296492 168812 296548
rect 168868 296492 168878 296548
rect 332546 296492 332556 296548
rect 332612 296492 334348 296548
rect 334404 296492 334414 296548
rect 335682 296492 335692 296548
rect 335748 296492 337820 296548
rect 337876 296492 337886 296548
rect 338930 296492 338940 296548
rect 338996 296492 339724 296548
rect 339780 296492 339790 296548
rect 332770 296268 332780 296324
rect 332836 296268 333340 296324
rect 333396 296268 333406 296324
rect 329896 296044 332780 296100
rect 332836 296044 332846 296100
rect 177650 295820 177660 295876
rect 177716 295820 180040 295876
rect 329634 295596 329644 295652
rect 329700 295596 329710 295652
rect 334226 295596 334236 295652
rect 334292 295596 334796 295652
rect 334852 295596 334862 295652
rect 329644 295176 329700 295596
rect 335122 295372 335132 295428
rect 335188 295372 340088 295428
rect 156258 294812 156268 294868
rect 156324 294812 165676 294868
rect 165732 294812 165742 294868
rect 176082 294700 176092 294756
rect 176148 294700 180040 294756
rect 335570 294700 335580 294756
rect 335636 294700 340396 294756
rect 340452 294700 340462 294756
rect 329896 294252 330988 294308
rect 331044 294252 331054 294308
rect 72118 293916 72156 293972
rect 72212 293916 72222 293972
rect 84578 293916 84588 293972
rect 84644 293916 85596 293972
rect 85652 293916 85662 293972
rect 334226 293916 334236 293972
rect 334292 293916 334684 293972
rect 334740 293916 334750 293972
rect 334450 293804 334460 293860
rect 334516 293804 335468 293860
rect 335524 293804 335534 293860
rect 333218 293692 333228 293748
rect 333284 293692 335244 293748
rect 335300 293692 335310 293748
rect 59042 293132 59052 293188
rect 59108 293132 108332 293188
rect 108388 293132 108398 293188
rect 180236 293076 180292 293608
rect 329868 293188 329924 293384
rect 332770 293356 332780 293412
rect 332836 293356 334684 293412
rect 334740 293356 334750 293412
rect 329868 293132 332780 293188
rect 332836 293132 333340 293188
rect 333396 293132 333406 293188
rect 180226 293020 180236 293076
rect 180292 293020 180302 293076
rect 26002 292460 26012 292516
rect 26068 292460 180040 292516
rect 329896 292460 333564 292516
rect 333620 292460 333630 292516
rect 46834 292348 46844 292404
rect 46900 292348 137788 292404
rect 137844 292348 137854 292404
rect 333442 292236 333452 292292
rect 333508 292236 336028 292292
rect 336084 292236 336094 292292
rect 329896 291564 333004 291620
rect 333060 291564 333070 291620
rect 27682 291340 27692 291396
rect 27748 291340 180040 291396
rect -960 290836 480 291032
rect 335346 291004 335356 291060
rect 335412 291004 339948 291060
rect 340004 291004 340014 291060
rect -960 290808 4172 290836
rect 392 290780 4172 290808
rect 4228 290780 4238 290836
rect 329896 290668 332780 290724
rect 332836 290668 332846 290724
rect 335010 290332 335020 290388
rect 335076 290332 338268 290388
rect 338324 290332 338334 290388
rect 10882 290220 10892 290276
rect 10948 290220 180040 290276
rect 329896 289772 332892 289828
rect 332948 289772 332958 289828
rect 4274 289212 4284 289268
rect 4340 289212 96012 289268
rect 96068 289212 96078 289268
rect 29362 289100 29372 289156
rect 29428 289100 180040 289156
rect 330866 289100 330876 289156
rect 330932 289100 336252 289156
rect 336308 289100 336318 289156
rect 139206 288988 139244 289044
rect 139300 288988 139310 289044
rect 330082 288988 330092 289044
rect 330148 288988 335636 289044
rect 335794 288988 335804 289044
rect 335860 288988 338044 289044
rect 338100 288988 338110 289044
rect 335580 288932 335636 288988
rect 90888 288876 162540 288932
rect 162596 288876 162606 288932
rect 329896 288876 332668 288932
rect 332724 288876 332734 288932
rect 335580 288876 340088 288932
rect 123442 287980 123452 288036
rect 123508 287980 180040 288036
rect 329896 287980 337036 288036
rect 337092 287980 337102 288036
rect 336690 287756 336700 287812
rect 336756 287756 339612 287812
rect 339668 287756 339678 287812
rect 332098 287420 332108 287476
rect 332164 287420 334796 287476
rect 334852 287420 334862 287476
rect 337362 287420 337372 287476
rect 337428 287420 338940 287476
rect 338996 287420 339006 287476
rect 330418 287308 330428 287364
rect 330484 287308 330988 287364
rect 331044 287308 331054 287364
rect 329896 287084 332668 287140
rect 332724 287084 332734 287140
rect 108322 286860 108332 286916
rect 108388 286860 180040 286916
rect 335346 286748 335356 286804
rect 335412 286748 338156 286804
rect 338212 286748 338222 286804
rect 329896 286188 336140 286244
rect 336196 286188 336206 286244
rect 178882 285964 178892 286020
rect 178948 285964 180572 286020
rect 180628 285964 180638 286020
rect 96002 285740 96012 285796
rect 96068 285740 180040 285796
rect 330530 285740 330540 285796
rect 330596 285740 334908 285796
rect 334964 285740 334974 285796
rect 93650 285628 93660 285684
rect 93716 285628 163884 285684
rect 163940 285628 163950 285684
rect 330306 285628 330316 285684
rect 330372 285628 330876 285684
rect 330932 285628 330942 285684
rect 335234 285516 335244 285572
rect 335300 285516 335580 285572
rect 335636 285516 335646 285572
rect 155362 285292 155372 285348
rect 155428 285292 180068 285348
rect 329896 285292 330316 285348
rect 330372 285292 330382 285348
rect 93426 284732 93436 284788
rect 93492 284732 161308 284788
rect 161364 284732 161374 284788
rect 90888 284620 161868 284676
rect 161924 284620 161934 284676
rect 180012 284648 180068 285292
rect 595560 284676 597000 284872
rect 585442 284620 585452 284676
rect 585508 284648 597000 284676
rect 585508 284620 595672 284648
rect 329896 284396 333900 284452
rect 333956 284396 333966 284452
rect 160888 283948 180460 284004
rect 180516 283948 180526 284004
rect 334114 283836 334124 283892
rect 334180 283836 335020 283892
rect 335076 283836 335086 283892
rect 335346 283836 335356 283892
rect 335412 283836 336140 283892
rect 336196 283836 336206 283892
rect 332434 283724 332444 283780
rect 332500 283724 334348 283780
rect 334404 283724 334414 283780
rect 160402 283500 160412 283556
rect 160468 283500 180040 283556
rect 329896 283500 334908 283556
rect 334964 283500 334974 283556
rect 329298 282604 329308 282660
rect 329364 282604 329374 282660
rect 165442 282380 165452 282436
rect 165508 282380 180040 282436
rect 336690 282380 336700 282436
rect 336756 282380 340088 282436
rect 162530 282156 162540 282212
rect 162596 282156 163436 282212
rect 163492 282156 163502 282212
rect 332098 282156 332108 282212
rect 332164 282156 333116 282212
rect 333172 282156 333182 282212
rect 335318 282156 335356 282212
rect 335412 282156 335422 282212
rect 160888 281932 178892 281988
rect 178948 281932 178958 281988
rect 329896 281708 334460 281764
rect 334516 281708 334526 281764
rect 332658 281372 332668 281428
rect 332724 281372 334796 281428
rect 334852 281372 334862 281428
rect 162082 281260 162092 281316
rect 162148 281260 180040 281316
rect 329868 280644 329924 280840
rect 334534 280812 334572 280868
rect 334628 280812 334638 280868
rect 329868 280588 335020 280644
rect 335076 280588 335086 280644
rect 161858 280476 161868 280532
rect 161924 280476 163996 280532
rect 164052 280476 164062 280532
rect 90888 280364 93660 280420
rect 93716 280364 93726 280420
rect 170482 280140 170492 280196
rect 170548 280140 180040 280196
rect 160888 279916 179900 279972
rect 179956 279916 179966 279972
rect 329896 279916 333116 279972
rect 333172 279916 333182 279972
rect 329868 279580 330092 279636
rect 330148 279580 330158 279636
rect 168802 279020 168812 279076
rect 168868 279020 180040 279076
rect 329868 279048 329924 279580
rect 329896 278124 339500 278180
rect 339556 278124 339566 278180
rect 160860 278012 168924 278068
rect 168980 278012 168990 278068
rect 160860 277928 160916 278012
rect 167122 277900 167132 277956
rect 167188 277900 180040 277956
rect 329868 277788 337708 277844
rect 337764 277788 337774 277844
rect 329868 277256 329924 277788
rect 330530 277564 330540 277620
rect 330596 277564 338940 277620
rect 338996 277564 339006 277620
rect 335682 277452 335692 277508
rect 335748 277452 336532 277508
rect 336476 277396 336532 277452
rect 335122 277340 335132 277396
rect 335188 277340 336028 277396
rect 336084 277340 336094 277396
rect 336476 277340 337932 277396
rect 337988 277340 337998 277396
rect 335570 277228 335580 277284
rect 335636 277228 336700 277284
rect 336756 277228 336766 277284
rect -960 276724 480 276920
rect 168802 276780 168812 276836
rect 168868 276780 180040 276836
rect -960 276696 34412 276724
rect 392 276668 34412 276696
rect 34468 276668 34478 276724
rect 334226 276556 334236 276612
rect 334292 276556 337820 276612
rect 337876 276556 337886 276612
rect 329896 276332 332668 276388
rect 332724 276332 332734 276388
rect 90888 276108 93996 276164
rect 94052 276108 94062 276164
rect 160888 275884 164108 275940
rect 164164 275884 164174 275940
rect 333106 275884 333116 275940
rect 333172 275884 334572 275940
rect 334628 275884 334638 275940
rect 336578 275884 336588 275940
rect 336644 275884 337596 275940
rect 337652 275884 340088 275940
rect 165442 275660 165452 275716
rect 165508 275660 180040 275716
rect 333442 275660 333452 275716
rect 333508 275660 337708 275716
rect 337764 275660 337774 275716
rect 163762 275548 163772 275604
rect 163828 275548 168476 275604
rect 168532 275548 168542 275604
rect 330642 275548 330652 275604
rect 330708 275548 332108 275604
rect 332164 275548 332174 275604
rect 334114 275548 334124 275604
rect 334180 275548 334572 275604
rect 334628 275548 334638 275604
rect 329868 275268 329924 275464
rect 329868 275212 340396 275268
rect 340452 275212 340462 275268
rect 170482 274540 170492 274596
rect 170548 274540 180040 274596
rect 329896 274540 330988 274596
rect 331044 274540 331054 274596
rect 160888 273868 169036 273924
rect 169092 273868 169102 273924
rect 332546 273868 332556 273924
rect 332612 273868 334348 273924
rect 334404 273868 334414 273924
rect 329896 273644 333564 273700
rect 333620 273644 333630 273700
rect 179666 273420 179676 273476
rect 179732 273420 180040 273476
rect 329868 273308 330876 273364
rect 330932 273308 330942 273364
rect 329868 272776 329924 273308
rect 330754 272636 330764 272692
rect 330820 272636 332892 272692
rect 332948 272636 332958 272692
rect 179554 272300 179564 272356
rect 179620 272300 180040 272356
rect 90888 271852 93436 271908
rect 93492 271852 93502 271908
rect 160888 271852 165564 271908
rect 165620 271852 165630 271908
rect 329896 271852 332892 271908
rect 332948 271852 332958 271908
rect 595560 271460 597000 271656
rect 590930 271404 590940 271460
rect 590996 271432 597000 271460
rect 590996 271404 595672 271432
rect 179666 271180 179676 271236
rect 179732 271180 180040 271236
rect 329532 270564 329588 270984
rect 332434 270956 332444 271012
rect 332500 270956 334348 271012
rect 334404 270956 334414 271012
rect 329522 270508 329532 270564
rect 329588 270508 329598 270564
rect 180002 270396 180012 270452
rect 180068 270396 180078 270452
rect 334114 270396 334124 270452
rect 334180 270396 335132 270452
rect 335188 270396 335198 270452
rect 180012 270088 180068 270396
rect 329896 270060 337932 270116
rect 337988 270060 337998 270116
rect 160888 269836 167244 269892
rect 167300 269836 167310 269892
rect 337250 269388 337260 269444
rect 337316 269388 340088 269444
rect 329896 269164 334348 269220
rect 334404 269164 334414 269220
rect 172946 268940 172956 268996
rect 173012 268940 180040 268996
rect 334786 268940 334796 268996
rect 334852 268940 337820 268996
rect 337876 268940 337886 268996
rect 335458 268828 335468 268884
rect 335524 268828 337708 268884
rect 337764 268828 337774 268884
rect 331538 268716 331548 268772
rect 331604 268716 332108 268772
rect 332164 268716 332174 268772
rect 329896 268268 332780 268324
rect 332836 268268 332846 268324
rect 332322 268044 332332 268100
rect 332388 268044 338156 268100
rect 338212 268044 338222 268100
rect 160888 267820 163436 267876
rect 163492 267820 163502 267876
rect 172834 267820 172844 267876
rect 172900 267820 180040 267876
rect 90888 267596 106652 267652
rect 106708 267596 106718 267652
rect 335906 267596 335916 267652
rect 335972 267596 338940 267652
rect 338996 267596 339006 267652
rect 329868 267204 329924 267400
rect 329868 267148 330540 267204
rect 330596 267148 330606 267204
rect 174626 266700 174636 266756
rect 174692 266700 180040 266756
rect 329896 266476 332668 266532
rect 332724 266476 332734 266532
rect 334226 266252 334236 266308
rect 334292 266252 336140 266308
rect 336196 266252 336206 266308
rect 160888 265804 163996 265860
rect 164052 265804 164062 265860
rect 176306 265580 176316 265636
rect 176372 265580 180040 265636
rect 329298 265580 329308 265636
rect 329364 265580 329374 265636
rect 330194 265468 330204 265524
rect 330260 265468 331884 265524
rect 331940 265468 331950 265524
rect 335010 265468 335020 265524
rect 335076 265468 337372 265524
rect 337428 265468 337438 265524
rect 180562 265020 180572 265076
rect 180628 265020 180638 265076
rect 180572 264488 180628 265020
rect 329896 264684 333340 264740
rect 333396 264684 333406 264740
rect 335346 264684 335356 264740
rect 335412 264684 340396 264740
rect 340452 264684 340462 264740
rect 331650 264572 331660 264628
rect 331716 264572 337932 264628
rect 337988 264572 337998 264628
rect 329858 264236 329868 264292
rect 329924 264236 333004 264292
rect 333060 264236 333070 264292
rect 332322 264124 332332 264180
rect 332388 264124 336028 264180
rect 336084 264124 336094 264180
rect 329756 264012 330148 264068
rect 330530 264012 330540 264068
rect 330596 264012 331324 264068
rect 331380 264012 331390 264068
rect 332770 264012 332780 264068
rect 332836 264012 336252 264068
rect 336308 264012 336318 264068
rect 160888 263788 163884 263844
rect 163940 263788 163950 263844
rect 329756 263816 329812 264012
rect 330092 263956 330148 264012
rect 330092 263900 336028 263956
rect 336084 263900 336094 263956
rect 330530 263788 330540 263844
rect 330596 263788 330764 263844
rect 330820 263788 330830 263844
rect 333554 263788 333564 263844
rect 333620 263788 335132 263844
rect 335188 263788 335198 263844
rect 334114 263676 334124 263732
rect 334180 263676 338380 263732
rect 338436 263676 338446 263732
rect 90888 263340 93436 263396
rect 93492 263340 93502 263396
rect 180002 263340 180012 263396
rect 180068 263340 180078 263396
rect 329896 262892 333788 262948
rect 333844 262892 333854 262948
rect 336914 262892 336924 262948
rect 336980 262892 337484 262948
rect 337540 262892 340088 262948
rect 392 262808 4284 262836
rect -960 262780 4284 262808
rect 4340 262780 4350 262836
rect -960 262584 480 262780
rect 180002 262220 180012 262276
rect 180068 262220 180078 262276
rect 329896 261996 332668 262052
rect 332724 261996 332734 262052
rect 160328 261800 163772 261828
rect 160300 261772 163772 261800
rect 163828 261772 163838 261828
rect 160300 261716 160356 261772
rect 138674 261660 138684 261716
rect 138740 261660 160356 261716
rect 332322 261436 332332 261492
rect 332388 261436 332612 261492
rect 332556 261380 332612 261436
rect 332546 261324 332556 261380
rect 332612 261324 332622 261380
rect 180674 261100 180684 261156
rect 180740 261100 180750 261156
rect 329896 261100 333340 261156
rect 333396 261100 333406 261156
rect 330082 260876 330092 260932
rect 330148 260876 333452 260932
rect 333508 260876 333518 260932
rect 335906 260428 335916 260484
rect 335972 260428 337708 260484
rect 337764 260428 337774 260484
rect 330306 260316 330316 260372
rect 330372 260316 333228 260372
rect 333284 260316 333294 260372
rect 334226 260316 334236 260372
rect 334292 260316 335468 260372
rect 335524 260316 335534 260372
rect 180674 259980 180684 260036
rect 180740 259980 180750 260036
rect 329868 259700 329924 260232
rect 330082 259868 330092 259924
rect 330148 259868 334684 259924
rect 334740 259868 334750 259924
rect 329868 259644 338380 259700
rect 338436 259644 338446 259700
rect 329410 259532 329420 259588
rect 329476 259532 335244 259588
rect 335300 259532 335310 259588
rect 332322 259420 332332 259476
rect 332388 259420 335020 259476
rect 335076 259420 335086 259476
rect 329896 259308 336476 259364
rect 336532 259308 336542 259364
rect 90888 259084 163212 259140
rect 163268 259084 163278 259140
rect 180674 258860 180684 258916
rect 180740 258860 180750 258916
rect 332770 258860 332780 258916
rect 332836 258860 334572 258916
rect 334628 258860 334638 258916
rect 333666 258748 333676 258804
rect 333732 258748 334908 258804
rect 334964 258748 334974 258804
rect 329970 258636 329980 258692
rect 330036 258636 330876 258692
rect 330932 258636 330942 258692
rect 330866 258524 330876 258580
rect 330932 258524 331660 258580
rect 331716 258524 331726 258580
rect 329896 258412 332780 258468
rect 332836 258412 332846 258468
rect 595560 258244 597000 258440
rect 591042 258188 591052 258244
rect 591108 258216 597000 258244
rect 591108 258188 595672 258216
rect 180572 257236 180628 257768
rect 329896 257516 336252 257572
rect 336308 257516 336318 257572
rect 180562 257180 180572 257236
rect 180628 257180 180638 257236
rect 336018 257180 336028 257236
rect 336084 257180 337932 257236
rect 337988 257180 337998 257236
rect 333666 257068 333676 257124
rect 333732 257068 334796 257124
rect 334852 257068 334862 257124
rect 335906 257068 335916 257124
rect 335972 257068 336140 257124
rect 336196 257068 336206 257124
rect 338370 257068 338380 257124
rect 338436 257068 339500 257124
rect 339556 257068 339566 257124
rect 331202 256956 331212 257012
rect 331268 256956 332668 257012
rect 332724 256956 332734 257012
rect 179666 256620 179676 256676
rect 179732 256620 180040 256676
rect 329868 256116 329924 256648
rect 331874 256396 331884 256452
rect 331940 256396 337596 256452
rect 337652 256396 340088 256452
rect 332994 256172 333004 256228
rect 333060 256172 334348 256228
rect 334404 256172 334414 256228
rect 329868 256060 330204 256116
rect 330260 256060 330270 256116
rect 329896 255724 333116 255780
rect 333172 255724 333182 255780
rect 180338 255500 180348 255556
rect 180404 255500 180414 255556
rect 334226 255276 334236 255332
rect 334292 255276 335692 255332
rect 335748 255276 335758 255332
rect 337922 254940 337932 254996
rect 337988 254940 338044 254996
rect 338100 254940 338110 254996
rect 90888 254828 93324 254884
rect 93380 254828 93390 254884
rect 329896 254828 333228 254884
rect 333284 254828 333294 254884
rect 332434 254604 332444 254660
rect 332500 254604 337708 254660
rect 337764 254604 337774 254660
rect 176978 254380 176988 254436
rect 177044 254380 180040 254436
rect 329896 253932 336252 253988
rect 336308 253932 336318 253988
rect 332210 253708 332220 253764
rect 332276 253708 334908 253764
rect 334964 253708 334974 253764
rect 333778 253596 333788 253652
rect 333844 253596 334684 253652
rect 334740 253596 334750 253652
rect 337810 253596 337820 253652
rect 337876 253596 339052 253652
rect 339108 253596 339118 253652
rect 336466 253484 336476 253540
rect 336532 253484 339724 253540
rect 339780 253484 339790 253540
rect 180572 252756 180628 253288
rect 332658 253148 332668 253204
rect 332724 253148 336252 253204
rect 336308 253148 336318 253204
rect 180562 252700 180572 252756
rect 180628 252700 180638 252756
rect 329868 252532 329924 253064
rect 329868 252476 330092 252532
rect 330148 252476 330158 252532
rect 329970 252364 329980 252420
rect 330036 252364 331212 252420
rect 331268 252364 331278 252420
rect 180674 252140 180684 252196
rect 180740 252140 180750 252196
rect 329896 252140 336028 252196
rect 336084 252140 336094 252196
rect 330418 252028 330428 252084
rect 330484 252028 333452 252084
rect 333508 252028 333518 252084
rect 329896 251244 333788 251300
rect 333844 251244 333854 251300
rect 177538 251020 177548 251076
rect 177604 251020 180040 251076
rect 330754 250684 330764 250740
rect 330820 250684 333564 250740
rect 333620 250684 333630 250740
rect 90888 250572 92428 250628
rect 92484 250572 93324 250628
rect 93380 250572 93390 250628
rect 329868 250572 333452 250628
rect 333508 250572 333518 250628
rect 329868 250376 329924 250572
rect 331650 250460 331660 250516
rect 331716 250460 334236 250516
rect 334292 250460 334302 250516
rect 330530 250348 330540 250404
rect 330596 250348 330764 250404
rect 330820 250348 330830 250404
rect 332434 250348 332444 250404
rect 332500 250348 332780 250404
rect 332836 250348 332846 250404
rect 336466 250236 336476 250292
rect 336532 250236 337260 250292
rect 337316 250236 337326 250292
rect 335906 250124 335916 250180
rect 335972 250124 338044 250180
rect 338100 250124 338110 250180
rect 332658 249900 332668 249956
rect 332724 249900 340088 249956
rect 329868 248948 329924 249480
rect 332322 249452 332332 249508
rect 332388 249452 332780 249508
rect 332836 249452 332846 249508
rect 329868 248892 333004 248948
rect 333060 248892 333070 248948
rect 335878 248780 335916 248836
rect 335972 248780 335982 248836
rect -960 248500 480 248696
rect 331174 248668 331212 248724
rect 331268 248668 331278 248724
rect 337894 248668 337932 248724
rect 337988 248668 337998 248724
rect 338258 248668 338268 248724
rect 338324 248668 338334 248724
rect 338268 248612 338324 248668
rect 329896 248556 332780 248612
rect 332836 248556 332846 248612
rect 338268 248556 339948 248612
rect 340004 248556 340014 248612
rect -960 248472 4620 248500
rect 392 248444 4620 248472
rect 4676 248444 4686 248500
rect 329868 247044 329924 247688
rect 337250 247100 337260 247156
rect 337316 247100 339500 247156
rect 339556 247100 339566 247156
rect 329868 246988 330988 247044
rect 331044 246988 331054 247044
rect 334898 246988 334908 247044
rect 334964 246988 336028 247044
rect 336084 246988 336094 247044
rect 336578 246988 336588 247044
rect 336644 246988 337372 247044
rect 337428 246988 337438 247044
rect 339042 246988 339052 247044
rect 339108 246988 339276 247044
rect 339332 246988 339342 247044
rect 330306 246876 330316 246932
rect 330372 246876 331884 246932
rect 331940 246876 331950 246932
rect 332434 246876 332444 246932
rect 332500 246876 334124 246932
rect 334180 246876 334190 246932
rect 337250 246876 337260 246932
rect 337316 246876 337596 246932
rect 337652 246876 337662 246932
rect 339462 246876 339500 246932
rect 339556 246876 339566 246932
rect 329896 246764 333452 246820
rect 333508 246764 333518 246820
rect 90888 246316 93212 246372
rect 93268 246316 93436 246372
rect 93492 246316 93502 246372
rect 329756 245364 329812 245896
rect 333218 245420 333228 245476
rect 333284 245420 337932 245476
rect 337988 245420 337998 245476
rect 329746 245308 329756 245364
rect 329812 245308 329822 245364
rect 333666 245308 333676 245364
rect 333732 245308 333742 245364
rect 334786 245308 334796 245364
rect 334852 245308 335916 245364
rect 335972 245308 335982 245364
rect 333676 245252 333732 245308
rect 331538 245196 331548 245252
rect 331604 245196 332108 245252
rect 332164 245196 332174 245252
rect 333676 245196 336028 245252
rect 336084 245196 336094 245252
rect 595560 245028 597000 245224
rect 330530 244972 330540 245028
rect 330596 244972 332108 245028
rect 332164 244972 332174 245028
rect 587122 244972 587132 245028
rect 587188 245000 597000 245028
rect 587188 244972 595672 245000
rect 330866 244860 330876 244916
rect 330932 244860 334236 244916
rect 334292 244860 334302 244916
rect 335906 244076 335916 244132
rect 335972 244076 336476 244132
rect 336532 244076 336542 244132
rect 334226 243740 334236 243796
rect 334292 243740 337708 243796
rect 337764 243740 337774 243796
rect 332322 243628 332332 243684
rect 332388 243628 332398 243684
rect 332332 243572 332388 243628
rect 332332 243516 333228 243572
rect 333284 243516 333294 243572
rect 333442 243516 333452 243572
rect 333508 243516 333900 243572
rect 333956 243516 333966 243572
rect 336018 243516 336028 243572
rect 336084 243516 337820 243572
rect 337876 243516 337886 243572
rect 332658 243404 332668 243460
rect 332724 243404 332780 243460
rect 332836 243404 332846 243460
rect 333666 243404 333676 243460
rect 333732 243404 340088 243460
rect 334114 243180 334124 243236
rect 334180 243180 336924 243236
rect 336980 243180 336990 243236
rect 90888 242060 92596 242116
rect 330950 242060 330988 242116
rect 331044 242060 331054 242116
rect 92540 242004 92596 242060
rect 92530 241948 92540 242004
rect 92596 241948 93212 242004
rect 93268 241948 93278 242004
rect 329410 241948 329420 242004
rect 329476 241948 332892 242004
rect 332948 241948 332958 242004
rect 338930 241948 338940 242004
rect 338996 241948 339052 242004
rect 339108 241948 339118 242004
rect 335458 241164 335468 241220
rect 335524 241164 339500 241220
rect 339556 241164 339566 241220
rect 332434 240716 332444 240772
rect 332500 240716 338156 240772
rect 338212 240716 338222 240772
rect 48290 240604 48300 240660
rect 48356 240604 118412 240660
rect 118468 240604 118478 240660
rect 314132 240604 326508 240660
rect 326564 240604 332220 240660
rect 332276 240604 332286 240660
rect 314132 240548 314188 240604
rect 60834 240492 60844 240548
rect 60900 240492 197372 240548
rect 197428 240492 197438 240548
rect 202514 240492 202524 240548
rect 202580 240492 314188 240548
rect 327954 240492 327964 240548
rect 328020 240492 337708 240548
rect 337764 240492 337774 240548
rect 44706 240380 44716 240436
rect 44772 240380 113372 240436
rect 113428 240380 113438 240436
rect 199154 240380 199164 240436
rect 199220 240380 294812 240436
rect 294868 240380 294878 240436
rect 327506 240380 327516 240436
rect 327572 240380 329980 240436
rect 330036 240380 330046 240436
rect 53666 240268 53676 240324
rect 53732 240268 116732 240324
rect 116788 240268 116798 240324
rect 328514 240268 328524 240324
rect 328580 240268 329196 240324
rect 329252 240268 329262 240324
rect 330194 240268 330204 240324
rect 330260 240268 331212 240324
rect 331268 240268 331278 240324
rect 332434 240268 332444 240324
rect 332500 240268 336364 240324
rect 336420 240268 336430 240324
rect 50082 240156 50092 240212
rect 50148 240156 160412 240212
rect 160468 240156 160478 240212
rect 334562 240156 334572 240212
rect 334628 240156 335132 240212
rect 335188 240156 335198 240212
rect 66210 240044 66220 240100
rect 66276 240044 178892 240100
rect 178948 240044 178958 240100
rect 184818 240044 184828 240100
rect 184884 240044 184940 240100
rect 184996 240044 185006 240100
rect 202402 240044 202412 240100
rect 202468 240044 334460 240100
rect 334516 240044 334526 240100
rect 335010 240044 335020 240100
rect 335076 240044 335356 240100
rect 335412 240044 335422 240100
rect 334460 239988 334516 240044
rect 4162 239932 4172 239988
rect 4228 239932 204428 239988
rect 204484 239932 208348 239988
rect 334460 239932 335580 239988
rect 335636 239932 335646 239988
rect 208292 239876 208348 239932
rect 57250 239820 57260 239876
rect 57316 239820 104972 239876
rect 105028 239820 105038 239876
rect 208292 239820 270172 239876
rect 270228 239820 270238 239876
rect 321794 239820 321804 239876
rect 321860 239820 329420 239876
rect 329476 239820 329486 239876
rect 334226 239820 334236 239876
rect 334292 239820 339836 239876
rect 339892 239820 339902 239876
rect 85922 239708 85932 239764
rect 85988 239708 111692 239764
rect 111748 239708 111758 239764
rect 177538 239708 177548 239764
rect 177604 239708 268044 239764
rect 268100 239708 268110 239764
rect 284722 239708 284732 239764
rect 284788 239708 333340 239764
rect 333396 239708 333406 239764
rect 177202 239596 177212 239652
rect 177268 239596 275660 239652
rect 275716 239596 275726 239652
rect 278114 239596 278124 239652
rect 278180 239596 333564 239652
rect 333620 239596 333630 239652
rect 177650 239484 177660 239540
rect 177716 239484 278348 239540
rect 278404 239484 278414 239540
rect 281362 239484 281372 239540
rect 281428 239484 331660 239540
rect 331716 239484 331726 239540
rect 77298 239372 77308 239428
rect 77364 239372 179116 239428
rect 179172 239372 179182 239428
rect 186274 239372 186284 239428
rect 186340 239372 204316 239428
rect 204372 239372 334460 239428
rect 334516 239372 334526 239428
rect 186386 239260 186396 239316
rect 186452 239260 335356 239316
rect 335412 239260 335422 239316
rect 314132 238812 335132 238868
rect 335188 238812 335198 238868
rect 228508 238700 287308 238756
rect 287364 238700 287374 238756
rect 37986 238476 37996 238532
rect 38052 238476 42924 238532
rect 42980 238476 42990 238532
rect 87714 238476 87724 238532
rect 87780 238476 99932 238532
rect 99988 238476 99998 238532
rect 184930 238476 184940 238532
rect 184996 238476 186396 238532
rect 186452 238476 186462 238532
rect 228508 238420 228564 238700
rect 314132 238644 314188 238812
rect 329074 238700 329084 238756
rect 329140 238700 332668 238756
rect 332724 238700 332734 238756
rect 243572 238588 314188 238644
rect 331510 238588 331548 238644
rect 331604 238588 331614 238644
rect 332322 238588 332332 238644
rect 332388 238588 335468 238644
rect 335524 238588 335534 238644
rect 243572 238532 243628 238588
rect 38210 238364 38220 238420
rect 38276 238364 46508 238420
rect 46564 238364 46574 238420
rect 64418 238364 64428 238420
rect 64484 238364 77308 238420
rect 77364 238364 77374 238420
rect 80546 238364 80556 238420
rect 80612 238364 95116 238420
rect 95172 238364 95182 238420
rect 138562 238364 138572 238420
rect 138628 238364 204764 238420
rect 204820 238364 228564 238420
rect 231812 238476 243628 238532
rect 251234 238476 251244 238532
rect 251300 238476 281820 238532
rect 281876 238476 281886 238532
rect 332658 238476 332668 238532
rect 332724 238476 334684 238532
rect 334740 238476 334750 238532
rect 231812 238308 231868 238476
rect 239586 238364 239596 238420
rect 239652 238364 272188 238420
rect 272244 238364 272254 238420
rect 307682 238364 307692 238420
rect 307748 238364 325388 238420
rect 325444 238364 325454 238420
rect 40114 238252 40124 238308
rect 40180 238252 51884 238308
rect 51940 238252 51950 238308
rect 84130 238252 84140 238308
rect 84196 238252 94892 238308
rect 94948 238252 94958 238308
rect 187506 238252 187516 238308
rect 187572 238252 231868 238308
rect 243170 238252 243180 238308
rect 243236 238252 275884 238308
rect 275940 238252 275950 238308
rect 295250 238252 295260 238308
rect 295316 238252 302428 238308
rect 305890 238252 305900 238308
rect 305956 238252 324268 238308
rect 324324 238252 324334 238308
rect 325826 238252 325836 238308
rect 325892 238252 330316 238308
rect 330372 238252 330382 238308
rect 38322 238140 38332 238196
rect 38388 238140 55468 238196
rect 55524 238140 55534 238196
rect 75170 238140 75180 238196
rect 75236 238140 95340 238196
rect 95396 238140 95406 238196
rect 237794 238140 237804 238196
rect 237860 238140 270620 238196
rect 270676 238140 270686 238196
rect 282034 238140 282044 238196
rect 282100 238140 297836 238196
rect 297892 238140 297902 238196
rect 302372 238084 302428 238252
rect 304098 238140 304108 238196
rect 304164 238140 325164 238196
rect 325220 238140 325230 238196
rect 325714 238140 325724 238196
rect 325780 238140 330876 238196
rect 330932 238140 330942 238196
rect 78754 238028 78764 238084
rect 78820 238028 96796 238084
rect 96852 238028 96862 238084
rect 236002 238028 236012 238084
rect 236068 238028 268828 238084
rect 268884 238028 268894 238084
rect 294242 238028 294252 238084
rect 294308 238028 298284 238084
rect 298340 238028 298350 238084
rect 302372 238028 318444 238084
rect 318500 238028 318510 238084
rect 324482 238028 324492 238084
rect 324548 238028 336140 238084
rect 336196 238028 336206 238084
rect 40226 237916 40236 237972
rect 40292 237916 59052 237972
rect 59108 237916 59118 237972
rect 73378 237916 73388 237972
rect 73444 237916 162092 237972
rect 162148 237916 162158 237972
rect 242274 237916 242284 237972
rect 242340 237916 275660 237972
rect 275716 237916 275726 237972
rect 280354 237916 280364 237972
rect 280420 237916 291564 237972
rect 291620 237916 291630 237972
rect 296034 237916 296044 237972
rect 296100 237916 324940 237972
rect 324996 237916 325006 237972
rect 325826 237916 325836 237972
rect 325892 237916 337260 237972
rect 337316 237916 337326 237972
rect 69794 237804 69804 237860
rect 69860 237804 96572 237860
rect 96628 237804 96638 237860
rect 240482 237804 240492 237860
rect 240548 237804 273868 237860
rect 273924 237804 273934 237860
rect 287298 237804 287308 237860
rect 287364 237804 296548 237860
rect 298274 237804 298284 237860
rect 298340 237804 326732 237860
rect 326788 237804 326798 237860
rect 327506 237804 327516 237860
rect 327572 237804 337932 237860
rect 337988 237804 337998 237860
rect 296492 237748 296548 237804
rect 67974 237692 68012 237748
rect 68068 237692 68078 237748
rect 82338 237692 82348 237748
rect 82404 237692 103292 237748
rect 103348 237692 103358 237748
rect 238690 237692 238700 237748
rect 238756 237692 272636 237748
rect 272692 237692 272702 237748
rect 288866 237692 288876 237748
rect 288932 237692 292460 237748
rect 292516 237692 292526 237748
rect 296492 237692 327236 237748
rect 327394 237692 327404 237748
rect 327460 237692 330092 237748
rect 330148 237692 330158 237748
rect 327180 237636 327236 237692
rect 71558 237580 71596 237636
rect 71652 237580 71662 237636
rect 76962 237580 76972 237636
rect 77028 237580 91532 237636
rect 91588 237580 91598 237636
rect 252130 237580 252140 237636
rect 252196 237580 274764 237636
rect 274820 237580 274830 237636
rect 321122 237580 321132 237636
rect 321188 237580 326060 237636
rect 326116 237580 326126 237636
rect 327180 237580 327852 237636
rect 327908 237580 328972 237636
rect 329028 237580 329038 237636
rect 322914 237468 322924 237524
rect 322980 237468 325948 237524
rect 326004 237468 326014 237524
rect 285506 237356 285516 237412
rect 285572 237356 290668 237412
rect 290724 237356 290734 237412
rect 328850 237244 328860 237300
rect 328916 237244 335916 237300
rect 335972 237244 335982 237300
rect 235078 237132 235116 237188
rect 235172 237132 235182 237188
rect 280466 237132 280476 237188
rect 280532 237132 287980 237188
rect 288036 237132 288046 237188
rect 234182 237020 234220 237076
rect 234276 237020 234286 237076
rect 264450 237020 264460 237076
rect 264516 237020 265244 237076
rect 265300 237020 265310 237076
rect 268034 237020 268044 237076
rect 268100 237020 268716 237076
rect 268772 237020 268782 237076
rect 269826 237020 269836 237076
rect 269892 237020 270396 237076
rect 270452 237020 270462 237076
rect 275202 237020 275212 237076
rect 275268 237020 275324 237076
rect 275380 237020 275390 237076
rect 277890 237020 277900 237076
rect 277956 237020 278796 237076
rect 278852 237020 278862 237076
rect 282146 237020 282156 237076
rect 282212 237020 287084 237076
rect 287140 237020 287150 237076
rect 293906 237020 293916 237076
rect 293972 237020 296940 237076
rect 296996 237020 297006 237076
rect 226678 236908 226716 236964
rect 226772 236908 226782 236964
rect 231718 236908 231756 236964
rect 231812 236908 231822 236964
rect 233314 236908 233324 236964
rect 233380 236908 233436 236964
rect 233492 236908 233502 236964
rect 265318 236908 265356 236964
rect 265412 236908 265422 236964
rect 266242 236908 266252 236964
rect 266308 236908 266812 236964
rect 266868 236908 266878 236964
rect 266998 236908 267036 236964
rect 267092 236908 267102 236964
rect 268566 236908 268604 236964
rect 268660 236908 268670 236964
rect 270246 236908 270284 236964
rect 270340 236908 270350 236964
rect 272038 236908 272076 236964
rect 272132 236908 272142 236964
rect 275398 236908 275436 236964
rect 275492 236908 275502 236964
rect 276994 236908 277004 236964
rect 277060 236908 277116 236964
rect 277172 236908 277182 236964
rect 278646 236908 278684 236964
rect 278740 236908 278750 236964
rect 283826 236908 283836 236964
rect 283892 236908 288876 236964
rect 288932 236908 288942 236964
rect 290434 236908 290444 236964
rect 290500 236908 290556 236964
rect 290612 236908 290622 236964
rect 293766 236908 293804 236964
rect 293860 236908 293870 236964
rect 295334 236908 295372 236964
rect 295428 236908 295438 236964
rect 298918 236908 298956 236964
rect 299012 236908 299022 236964
rect 305638 236908 305676 236964
rect 305732 236908 305742 236964
rect 328962 236908 328972 236964
rect 329028 236908 340088 236964
rect 178882 236796 178892 236852
rect 178948 236796 191548 236852
rect 191604 236796 191614 236852
rect 325042 236796 325052 236852
rect 325108 236796 328636 236852
rect 328692 236796 328702 236852
rect 197698 236684 197708 236740
rect 197764 236684 282604 236740
rect 282660 236684 282670 236740
rect 289762 236684 289772 236740
rect 289828 236684 332668 236740
rect 332724 236684 332734 236740
rect 337362 236684 337372 236740
rect 337428 236684 339948 236740
rect 340004 236684 340014 236740
rect 187394 236572 187404 236628
rect 187460 236572 276556 236628
rect 276612 236572 276622 236628
rect 288082 236572 288092 236628
rect 288148 236572 329924 236628
rect 330082 236572 330092 236628
rect 330148 236572 337708 236628
rect 337764 236572 337774 236628
rect 329868 236516 329924 236572
rect 199378 236460 199388 236516
rect 199444 236460 308252 236516
rect 308308 236460 308318 236516
rect 324370 236460 324380 236516
rect 324436 236460 329812 236516
rect 329868 236460 332668 236516
rect 332724 236460 332734 236516
rect 329756 236404 329812 236460
rect 202962 236348 202972 236404
rect 203028 236348 326844 236404
rect 326900 236348 326910 236404
rect 329756 236348 337148 236404
rect 337204 236348 337214 236404
rect 191538 236236 191548 236292
rect 191604 236236 192556 236292
rect 192612 236236 330540 236292
rect 330596 236236 330606 236292
rect 38210 236124 38220 236180
rect 38276 236124 198380 236180
rect 198436 236124 198446 236180
rect 198930 236124 198940 236180
rect 198996 236124 330316 236180
rect 330372 236124 330382 236180
rect 36866 236012 36876 236068
rect 36932 236012 199276 236068
rect 199332 236012 199342 236068
rect 203298 236012 203308 236068
rect 203364 236012 204540 236068
rect 204596 236012 332668 236068
rect 332724 236012 332734 236068
rect 204082 235900 204092 235956
rect 204148 235900 280588 235956
rect 280644 235900 280654 235956
rect 326498 235900 326508 235956
rect 326564 235900 327404 235956
rect 327460 235900 327470 235956
rect 328962 235900 328972 235956
rect 329028 235900 332444 235956
rect 332500 235900 332510 235956
rect 189410 235788 189420 235844
rect 189476 235788 333676 235844
rect 333732 235788 333742 235844
rect 188066 235676 188076 235732
rect 188132 235676 203308 235732
rect 203364 235676 203374 235732
rect 183922 235116 183932 235172
rect 183988 235116 202524 235172
rect 202580 235116 202748 235172
rect 202804 235116 202814 235172
rect 225250 235116 225260 235172
rect 225316 235116 267260 235172
rect 267316 235116 267326 235172
rect 290098 235116 290108 235172
rect 290164 235116 326844 235172
rect 326900 235116 326910 235172
rect 224354 235004 224364 235060
rect 224420 235004 266924 235060
rect 266980 235004 266990 235060
rect 270162 235004 270172 235060
rect 270228 235004 280140 235060
rect 280196 235004 280206 235060
rect 285954 235004 285964 235060
rect 286020 235004 330092 235060
rect 330148 235004 330158 235060
rect 189298 234892 189308 234948
rect 189364 234892 289660 234948
rect 289716 234892 289726 234948
rect 289874 234892 289884 234948
rect 289940 234892 327516 234948
rect 327572 234892 327582 234948
rect 169250 234780 169260 234836
rect 169316 234780 290444 234836
rect 290500 234780 290510 234836
rect 172386 234668 172396 234724
rect 172452 234668 307244 234724
rect 307300 234668 307310 234724
rect -960 234388 480 234584
rect 41346 234556 41356 234612
rect 41412 234556 196588 234612
rect 196644 234556 196654 234612
rect 213602 234556 213612 234612
rect 213668 234556 271516 234612
rect 271572 234556 271582 234612
rect 291442 234556 291452 234612
rect 291508 234556 336140 234612
rect 336196 234556 336206 234612
rect 40002 234444 40012 234500
rect 40068 234444 195692 234500
rect 195748 234444 195758 234500
rect 200162 234444 200172 234500
rect 200228 234444 275772 234500
rect 275828 234444 275838 234500
rect 284722 234444 284732 234500
rect 284788 234444 333788 234500
rect 333844 234444 333854 234500
rect -960 234360 24332 234388
rect 392 234332 24332 234360
rect 24388 234332 24398 234388
rect 41234 234332 41244 234388
rect 41300 234332 197484 234388
rect 197540 234332 197550 234388
rect 202514 234332 202524 234388
rect 202580 234332 308476 234388
rect 308532 234332 308542 234388
rect 230626 234220 230636 234276
rect 230692 234220 254492 234276
rect 254548 234220 254558 234276
rect 285058 234220 285068 234276
rect 285124 234220 313964 234276
rect 314020 234220 314030 234276
rect 285170 234108 285180 234164
rect 285236 234108 313068 234164
rect 313124 234108 313134 234164
rect 42802 233436 42812 233492
rect 42868 233436 197820 233492
rect 197876 233436 198044 233492
rect 198100 233436 198110 233492
rect 202850 233436 202860 233492
rect 202916 233436 274092 233492
rect 274148 233436 274158 233492
rect 291554 233436 291564 233492
rect 291620 233436 327964 233492
rect 328020 233436 328030 233492
rect 62626 233324 62636 233380
rect 62692 233324 199052 233380
rect 199108 233324 199118 233380
rect 201954 233324 201964 233380
rect 202020 233324 275548 233380
rect 275604 233324 275614 233380
rect 288418 233324 288428 233380
rect 288484 233324 328748 233380
rect 328804 233324 328814 233380
rect 177874 233212 177884 233268
rect 177940 233212 269500 233268
rect 269556 233212 269566 233268
rect 281586 233212 281596 233268
rect 281652 233212 328412 233268
rect 328468 233212 328478 233268
rect 167570 233100 167580 233156
rect 167636 233100 293804 233156
rect 293860 233100 293870 233156
rect 172274 232988 172284 233044
rect 172340 232988 301644 233044
rect 301700 232988 301710 233044
rect 172722 232876 172732 232932
rect 172788 232876 315084 232932
rect 315140 232876 315150 232932
rect 325266 232876 325276 232932
rect 325332 232876 330988 232932
rect 331044 232876 331054 232932
rect 35186 232764 35196 232820
rect 35252 232764 191212 232820
rect 191268 232764 191278 232820
rect 198034 232764 198044 232820
rect 198100 232764 272300 232820
rect 272356 232764 272366 232820
rect 279794 232764 279804 232820
rect 279860 232764 330204 232820
rect 330260 232764 330270 232820
rect 22754 232652 22764 232708
rect 22820 232652 186732 232708
rect 186788 232652 186798 232708
rect 195682 232652 195692 232708
rect 195748 232652 335468 232708
rect 335524 232652 335534 232708
rect 208226 232540 208236 232596
rect 208292 232540 277452 232596
rect 277508 232540 277518 232596
rect 595560 231924 597000 232008
rect 591154 231868 591164 231924
rect 591220 231868 597000 231924
rect 209122 231756 209132 231812
rect 209188 231756 267484 231812
rect 267540 231756 267550 231812
rect 288194 231756 288204 231812
rect 288260 231756 328300 231812
rect 328356 231756 328366 231812
rect 595560 231784 597000 231868
rect 197586 231644 197596 231700
rect 197652 231644 275996 231700
rect 276052 231644 276062 231700
rect 286626 231644 286636 231700
rect 286692 231644 333228 231700
rect 333284 231644 333294 231700
rect 167906 231532 167916 231588
rect 167972 231532 272300 231588
rect 272356 231532 272366 231588
rect 281474 231532 281484 231588
rect 281540 231532 329532 231588
rect 329588 231532 329598 231588
rect 176194 231420 176204 231476
rect 176260 231420 305004 231476
rect 305060 231420 305070 231476
rect 166114 231308 166124 231364
rect 166180 231308 294924 231364
rect 294980 231308 294990 231364
rect 171266 231196 171276 231252
rect 171332 231196 319564 231252
rect 319620 231196 319630 231252
rect 41010 231084 41020 231140
rect 41076 231084 194796 231140
rect 194852 231084 194862 231140
rect 201058 231084 201068 231140
rect 201124 231084 330988 231140
rect 331044 231084 331054 231140
rect 41122 230972 41132 231028
rect 41188 230972 223468 231028
rect 223524 230972 223534 231028
rect 227042 230972 227052 231028
rect 227108 230972 268940 231028
rect 268996 230972 269006 231028
rect 284834 230972 284844 231028
rect 284900 230972 335804 231028
rect 335860 230972 335870 231028
rect 214498 230860 214508 230916
rect 214564 230860 271404 230916
rect 271460 230860 271470 230916
rect 289986 230860 289996 230916
rect 290052 230860 326620 230916
rect 326676 230860 326686 230916
rect 334562 230412 334572 230468
rect 334628 230412 340088 230468
rect 328626 230188 328636 230244
rect 328692 230188 334572 230244
rect 334628 230188 334638 230244
rect 207330 230076 207340 230132
rect 207396 230076 282268 230132
rect 282324 230076 282334 230132
rect 203746 229964 203756 230020
rect 203812 229964 278908 230020
rect 278964 229964 278974 230020
rect 166226 229852 166236 229908
rect 166292 229852 273308 229908
rect 273364 229852 273374 229908
rect 166002 229740 166012 229796
rect 166068 229740 291564 229796
rect 291620 229740 291630 229796
rect 174514 229628 174524 229684
rect 174580 229628 302764 229684
rect 302820 229628 302830 229684
rect 180114 229516 180124 229572
rect 180180 229516 318444 229572
rect 318500 229516 318510 229572
rect 37986 229404 37996 229460
rect 38052 229404 188524 229460
rect 188580 229404 188590 229460
rect 196130 229404 196140 229460
rect 196196 229404 325164 229460
rect 325220 229404 325230 229460
rect 186386 229292 186396 229348
rect 186452 229292 277228 229348
rect 277284 229292 277294 229348
rect 284946 229292 284956 229348
rect 285012 229292 339724 229348
rect 339780 229292 339790 229348
rect 212706 229180 212716 229236
rect 212772 229180 270844 229236
rect 270900 229180 270910 229236
rect 210914 228396 210924 228452
rect 210980 228396 268940 228452
rect 268996 228396 269006 228452
rect 176082 228284 176092 228340
rect 176148 228284 288204 228340
rect 288260 228284 288270 228340
rect 179330 228172 179340 228228
rect 179396 228172 298284 228228
rect 298340 228172 298350 228228
rect 170930 228060 170940 228116
rect 170996 228060 306124 228116
rect 306180 228060 306190 228116
rect 167794 227948 167804 228004
rect 167860 227948 320684 228004
rect 320740 227948 320750 228004
rect 39778 227836 39788 227892
rect 39844 227836 193900 227892
rect 193956 227836 193966 227892
rect 210018 227836 210028 227892
rect 210084 227836 268828 227892
rect 268884 227836 268894 227892
rect 13234 227724 13244 227780
rect 13300 227724 185836 227780
rect 185892 227724 185902 227780
rect 211810 227724 211820 227780
rect 211876 227724 271068 227780
rect 271124 227724 271134 227780
rect 39890 227612 39900 227668
rect 39956 227612 222572 227668
rect 222628 227612 222638 227668
rect 228834 227612 228844 227668
rect 228900 227612 270508 227668
rect 270564 227612 270574 227668
rect 279906 227612 279916 227668
rect 279972 227612 326732 227668
rect 326788 227612 326798 227668
rect 227938 227500 227948 227556
rect 228004 227500 269052 227556
rect 269108 227500 269118 227556
rect 202850 226492 202860 226548
rect 202916 226492 271292 226548
rect 271348 226492 271358 226548
rect 204642 226380 204652 226436
rect 204708 226380 278012 226436
rect 278068 226380 278078 226436
rect 177762 226268 177772 226324
rect 177828 226268 273980 226324
rect 274036 226268 274046 226324
rect 170818 226156 170828 226212
rect 170884 226156 297164 226212
rect 297220 226156 297230 226212
rect 201170 226044 201180 226100
rect 201236 226044 333788 226100
rect 333844 226044 333854 226100
rect 192882 225932 192892 225988
rect 192948 225932 330092 225988
rect 330148 225932 330158 225988
rect 201058 225036 201068 225092
rect 201124 225036 274204 225092
rect 274260 225036 274270 225092
rect 177314 224924 177324 224980
rect 177380 224924 270620 224980
rect 270676 224924 270686 224980
rect 172610 224812 172620 224868
rect 172676 224812 300412 224868
rect 300468 224812 300478 224868
rect 197922 224700 197932 224756
rect 197988 224700 337260 224756
rect 337316 224700 337326 224756
rect 171154 224588 171164 224644
rect 171220 224588 310604 224644
rect 310660 224588 310670 224644
rect 166226 224476 166236 224532
rect 166292 224476 321804 224532
rect 321860 224476 321870 224532
rect 41906 224364 41916 224420
rect 41972 224364 220780 224420
rect 220836 224364 220846 224420
rect 232418 224364 232428 224420
rect 232484 224364 274316 224420
rect 274372 224364 274382 224420
rect 93314 224252 93324 224308
rect 93380 224252 276332 224308
rect 276388 224252 276398 224308
rect 206434 224140 206444 224196
rect 206500 224140 279132 224196
rect 279188 224140 279198 224196
rect 333442 223916 333452 223972
rect 333508 223916 337372 223972
rect 337428 223916 340088 223972
rect 177426 223356 177436 223412
rect 177492 223356 275772 223412
rect 275828 223356 275838 223412
rect 172498 223244 172508 223300
rect 172564 223244 296044 223300
rect 296100 223244 296110 223300
rect 171042 223132 171052 223188
rect 171108 223132 303884 223188
rect 303940 223132 303950 223188
rect 167682 223020 167692 223076
rect 167748 223020 311724 223076
rect 311780 223020 311790 223076
rect 39666 222908 39676 222964
rect 39732 222908 189420 222964
rect 189476 222908 189486 222964
rect 194674 222908 194684 222964
rect 194740 222908 274988 222964
rect 275044 222908 275054 222964
rect 30370 222796 30380 222852
rect 30436 222796 187628 222852
rect 187684 222796 187694 222852
rect 202290 222796 202300 222852
rect 202356 222796 293356 222852
rect 293412 222796 293422 222852
rect 34402 222684 34412 222740
rect 34468 222684 216300 222740
rect 216356 222684 216366 222740
rect 247650 222684 247660 222740
rect 247716 222684 269836 222740
rect 269892 222684 269902 222740
rect 93426 222572 93436 222628
rect 93492 222572 326956 222628
rect 327012 222572 327022 222628
rect 250338 222460 250348 222516
rect 250404 222460 269612 222516
rect 269668 222460 269678 222516
rect 229730 221676 229740 221732
rect 229796 221676 270732 221732
rect 270788 221676 270798 221732
rect 205538 221564 205548 221620
rect 205604 221564 274428 221620
rect 274484 221564 274494 221620
rect 198146 221452 198156 221508
rect 198212 221452 282380 221508
rect 282436 221452 282446 221508
rect 199490 221340 199500 221396
rect 199556 221340 290668 221396
rect 290724 221340 290734 221396
rect 177650 221228 177660 221284
rect 177716 221228 273868 221284
rect 273924 221228 273934 221284
rect 174402 221116 174412 221172
rect 174468 221116 292684 221172
rect 292740 221116 292750 221172
rect 200722 221004 200732 221060
rect 200788 221004 326732 221060
rect 326788 221004 326798 221060
rect 167906 220892 167916 220948
rect 167972 220892 313964 220948
rect 314020 220892 314030 220948
rect -960 220276 480 220472
rect -960 220248 108332 220276
rect 392 220220 108332 220248
rect 108388 220220 108398 220276
rect 204866 219996 204876 220052
rect 204932 219996 276444 220052
rect 276500 219996 276510 220052
rect 174290 219884 174300 219940
rect 174356 219884 272524 219940
rect 272580 219884 272590 219940
rect 174290 219772 174300 219828
rect 174356 219772 289324 219828
rect 289380 219772 289390 219828
rect 176306 219660 176316 219716
rect 176372 219660 317324 219716
rect 317380 219660 317390 219716
rect 40898 219548 40908 219604
rect 40964 219548 190316 219604
rect 190372 219548 190382 219604
rect 192434 219548 192444 219604
rect 192500 219548 323932 219604
rect 323988 219548 323998 219604
rect 38546 219436 38556 219492
rect 38612 219436 217196 219492
rect 217252 219436 217262 219492
rect 260194 219436 260204 219492
rect 260260 219436 278124 219492
rect 278180 219436 278190 219492
rect 41458 219324 41468 219380
rect 41524 219324 221676 219380
rect 221732 219324 221742 219380
rect 258402 219324 258412 219380
rect 258468 219324 278348 219380
rect 278404 219324 278414 219380
rect 26562 219212 26572 219268
rect 26628 219212 323372 219268
rect 323428 219212 323438 219268
rect 261986 219100 261996 219156
rect 262052 219100 279692 219156
rect 279748 219100 279758 219156
rect 595560 218596 597000 218792
rect 591266 218540 591276 218596
rect 591332 218568 597000 218596
rect 591332 218540 595672 218568
rect 195794 218316 195804 218372
rect 195860 218316 293244 218372
rect 293300 218316 293310 218372
rect 171266 218204 171276 218260
rect 171332 218204 273196 218260
rect 273252 218204 273262 218260
rect 179666 218092 179676 218148
rect 179732 218092 283276 218148
rect 283332 218092 283342 218148
rect 174626 217980 174636 218036
rect 174692 217980 299404 218036
rect 299460 217980 299470 218036
rect 179442 217868 179452 217924
rect 179508 217868 316204 217924
rect 316260 217868 316270 217924
rect 169362 217756 169372 217812
rect 169428 217756 309372 217812
rect 309428 217756 309438 217812
rect 38434 217644 38444 217700
rect 38500 217644 219884 217700
rect 219940 217644 219950 217700
rect 244962 217644 244972 217700
rect 245028 217644 276444 217700
rect 276500 217644 276510 217700
rect 93202 217532 93212 217588
rect 93268 217532 323148 217588
rect 323204 217532 323214 217588
rect 326834 217532 326844 217588
rect 326900 217532 337148 217588
rect 337204 217532 340116 217588
rect 204642 217420 204652 217476
rect 204708 217420 277340 217476
rect 277396 217420 277406 217476
rect 340060 217448 340116 217532
rect 154914 216748 154924 216804
rect 154980 216748 160524 216804
rect 160580 216748 160590 216804
rect 244066 216636 244076 216692
rect 244132 216636 285852 216692
rect 285908 216636 285918 216692
rect 193330 216524 193340 216580
rect 193396 216524 281708 216580
rect 281764 216524 281774 216580
rect 179442 216412 179452 216468
rect 179508 216412 272636 216468
rect 272692 216412 272702 216468
rect 177090 216300 177100 216356
rect 177156 216300 271516 216356
rect 271572 216300 271582 216356
rect 169474 216188 169484 216244
rect 169540 216188 272860 216244
rect 272916 216188 272926 216244
rect 177874 216076 177884 216132
rect 177940 216076 288652 216132
rect 288708 216076 288718 216132
rect 169474 215964 169484 216020
rect 169540 215964 308364 216020
rect 308420 215964 308430 216020
rect 169586 215852 169596 215908
rect 169652 215852 312844 215908
rect 312900 215852 312910 215908
rect 256610 215740 256620 215796
rect 256676 215740 280028 215796
rect 280084 215740 280094 215796
rect 202626 214956 202636 215012
rect 202692 214956 285292 215012
rect 285348 214956 285358 215012
rect 192994 214844 193004 214900
rect 193060 214844 278236 214900
rect 278292 214844 278302 214900
rect 180338 214732 180348 214788
rect 180404 214732 271740 214788
rect 271796 214732 271806 214788
rect 187282 214620 187292 214676
rect 187348 214620 280252 214676
rect 280308 214620 280318 214676
rect 177762 214508 177772 214564
rect 177828 214508 285068 214564
rect 285124 214508 285134 214564
rect 40226 214396 40236 214452
rect 40292 214396 193004 214452
rect 193060 214396 193070 214452
rect 196354 214396 196364 214452
rect 196420 214396 323372 214452
rect 323428 214396 323438 214452
rect 38322 214284 38332 214340
rect 38388 214284 218092 214340
rect 218148 214284 218158 214340
rect 248546 214284 248556 214340
rect 248612 214284 278012 214340
rect 278068 214284 278078 214340
rect 33506 214172 33516 214228
rect 33572 214172 218988 214228
rect 219044 214172 219054 214228
rect 246754 214172 246764 214228
rect 246820 214172 283052 214228
rect 283108 214172 283118 214228
rect 337026 213948 337036 214004
rect 337092 213948 337148 214004
rect 337204 213948 337214 214004
rect 36082 213388 36092 213444
rect 36148 213388 337148 213444
rect 337204 213388 337214 213444
rect 177510 213276 177548 213332
rect 177604 213276 177614 213332
rect 255714 213276 255724 213332
rect 255780 213276 279804 213332
rect 279860 213276 279870 213332
rect 253922 213164 253932 213220
rect 253988 213164 278236 213220
rect 278292 213164 278302 213220
rect 236898 213052 236908 213108
rect 236964 213052 270508 213108
rect 270564 213052 270574 213108
rect 180226 212940 180236 212996
rect 180292 212940 269052 212996
rect 269108 212940 269118 212996
rect 177986 212828 177996 212884
rect 178052 212828 280028 212884
rect 280084 212828 280094 212884
rect 180002 212716 180012 212772
rect 180068 212716 293132 212772
rect 293188 212716 293198 212772
rect 40114 212604 40124 212660
rect 40180 212604 192108 212660
rect 192164 212604 192174 212660
rect 199266 212604 199276 212660
rect 199332 212604 281596 212660
rect 281652 212604 281662 212660
rect 24658 212492 24668 212548
rect 24724 212492 215404 212548
rect 215460 212492 215470 212548
rect 245858 212492 245868 212548
rect 245924 212492 325052 212548
rect 325108 212492 325118 212548
rect 261090 212380 261100 212436
rect 261156 212380 283052 212436
rect 283108 212380 283118 212436
rect 257506 211596 257516 211652
rect 257572 211596 267932 211652
rect 267988 211596 267998 211652
rect 273634 211596 273644 211652
rect 273700 211596 274876 211652
rect 274932 211596 274942 211652
rect 262882 211484 262892 211540
rect 262948 211484 281372 211540
rect 281428 211484 281438 211540
rect 254818 211372 254828 211428
rect 254884 211372 267708 211428
rect 267764 211372 267774 211428
rect 267922 211372 267932 211428
rect 267988 211372 274652 211428
rect 274708 211372 274718 211428
rect 253026 211260 253036 211316
rect 253092 211260 267932 211316
rect 267988 211260 267998 211316
rect 272738 211260 272748 211316
rect 272804 211260 278684 211316
rect 278740 211260 278750 211316
rect 249442 211148 249452 211204
rect 249508 211148 276780 211204
rect 276836 211148 276846 211204
rect 180226 211036 180236 211092
rect 180292 211036 273420 211092
rect 273476 211036 273486 211092
rect 267698 210924 267708 210980
rect 267764 210924 276556 210980
rect 276612 210924 276622 210980
rect 284946 210924 284956 210980
rect 285012 210924 312172 210980
rect 312228 210924 312238 210980
rect 337250 210924 337260 210980
rect 337316 210924 340088 210980
rect 4274 210812 4284 210868
rect 4340 210812 123452 210868
rect 123508 210812 123518 210868
rect 169586 210812 169596 210868
rect 169652 210812 327628 210868
rect 327684 210812 327694 210868
rect 259298 210700 259308 210756
rect 259364 210700 266756 210756
rect 267922 210700 267932 210756
rect 267988 210700 278460 210756
rect 278516 210700 278526 210756
rect 266700 210644 266756 210700
rect 176082 210588 176092 210644
rect 176148 210588 262108 210644
rect 266700 210588 271292 210644
rect 271348 210588 271358 210644
rect 262052 210532 262108 210588
rect 262052 210476 272524 210532
rect 272580 210476 272590 210532
rect 241350 210028 241388 210084
rect 241444 210028 241454 210084
rect 189522 209916 189532 209972
rect 189588 209916 273868 209972
rect 179554 209804 179564 209860
rect 179620 209804 269500 209860
rect 269556 209804 269566 209860
rect 272290 209804 272300 209860
rect 272356 209804 273196 209860
rect 273252 209804 273262 209860
rect 273812 209748 273868 209916
rect 176194 209692 176204 209748
rect 176260 209692 272412 209748
rect 272468 209692 272478 209748
rect 273812 209692 275548 209748
rect 275604 209692 275614 209748
rect 174514 209580 174524 209636
rect 174580 209580 272748 209636
rect 272804 209580 272814 209636
rect 174402 209468 174412 209524
rect 174468 209468 272748 209524
rect 272804 209468 272814 209524
rect 172946 209356 172956 209412
rect 173012 209356 272860 209412
rect 272916 209356 272926 209412
rect 273074 209132 273084 209188
rect 273140 209132 273308 209188
rect 273364 209132 273374 209188
rect 180114 209020 180124 209076
rect 180180 209020 269612 209076
rect 269668 209020 269678 209076
rect 241378 208908 241388 208964
rect 241444 208908 273980 208964
rect 274036 208908 274046 208964
rect 269490 207564 269500 207620
rect 269556 207564 269566 207620
rect 269500 207032 269556 207564
rect 392 206360 4060 206388
rect -960 206332 4060 206360
rect 4116 206332 4126 206388
rect 272934 206332 272972 206388
rect 273028 206332 273038 206388
rect -960 206136 480 206332
rect 595560 205380 597000 205576
rect 585554 205324 585564 205380
rect 585620 205352 597000 205380
rect 585620 205324 595672 205352
rect 269602 204764 269612 204820
rect 269668 204764 269678 204820
rect 269612 204120 269668 204764
rect 314132 204428 328636 204484
rect 328692 204428 340088 204484
rect 314132 204148 314188 204428
rect 276322 204092 276332 204148
rect 276388 204092 314188 204148
rect 270498 203308 270508 203364
rect 270564 203308 270574 203364
rect 270508 203140 270564 203308
rect 272178 203196 272188 203252
rect 272244 203196 272860 203252
rect 272916 203196 272926 203252
rect 270508 203084 270732 203140
rect 270788 203084 270798 203140
rect 295138 202748 295148 202804
rect 295204 202748 309484 202804
rect 309540 202748 309550 202804
rect 306786 202636 306796 202692
rect 306852 202636 325388 202692
rect 325444 202636 325454 202692
rect 308242 202524 308252 202580
rect 308308 202524 328412 202580
rect 328468 202524 328478 202580
rect 308466 202412 308476 202468
rect 308532 202412 335804 202468
rect 335860 202412 335870 202468
rect 269602 201404 269612 201460
rect 269668 201404 269678 201460
rect 269612 201208 269668 201404
rect 299404 200060 300300 200116
rect 300356 200060 300366 200116
rect 299404 199892 299460 200060
rect 299618 199948 299628 200004
rect 299684 199948 299694 200004
rect 301158 199948 301196 200004
rect 301252 199948 301262 200004
rect 301410 199948 301420 200004
rect 301476 199948 301514 200004
rect 320226 199948 320236 200004
rect 320292 199948 320302 200004
rect 322018 199948 322028 200004
rect 322084 199948 322094 200004
rect 326946 199948 326956 200004
rect 327012 199948 328524 200004
rect 328580 199948 328590 200004
rect 293682 199836 293692 199892
rect 293748 199836 299460 199892
rect 299628 199892 299684 199948
rect 299628 199836 319172 199892
rect 284610 199724 284620 199780
rect 284676 199724 314860 199780
rect 314916 199724 314926 199780
rect 283602 199612 283612 199668
rect 283668 199612 315756 199668
rect 315812 199612 315822 199668
rect 283714 199500 283724 199556
rect 283780 199500 316652 199556
rect 316708 199500 316718 199556
rect 319116 199444 319172 199836
rect 320236 199780 320292 199948
rect 322028 199892 322084 199948
rect 322028 199836 324604 199892
rect 324660 199836 324670 199892
rect 320236 199724 324268 199780
rect 324324 199724 324334 199780
rect 323810 199612 323820 199668
rect 323876 199612 326284 199668
rect 326340 199612 326350 199668
rect 319330 199500 319340 199556
rect 319396 199500 326508 199556
rect 326564 199500 326574 199556
rect 283378 199388 283388 199444
rect 283444 199388 302428 199444
rect 303202 199388 303212 199444
rect 303268 199388 303492 199444
rect 308550 199388 308588 199444
rect 308644 199388 308654 199444
rect 310370 199388 310380 199444
rect 310436 199388 310828 199444
rect 310884 199388 310894 199444
rect 311798 199388 311836 199444
rect 311892 199388 311902 199444
rect 314132 199388 317548 199444
rect 317604 199388 317614 199444
rect 319116 199388 325276 199444
rect 325332 199388 325342 199444
rect 272290 199164 272300 199220
rect 272356 199164 273756 199220
rect 273812 199164 273822 199220
rect 302372 199108 302428 199388
rect 303436 199332 303492 199388
rect 303436 199276 310268 199332
rect 310324 199276 310334 199332
rect 314132 199220 314188 199388
rect 303436 199164 314188 199220
rect 303436 199108 303492 199164
rect 290434 199052 290444 199108
rect 290500 199052 301420 199108
rect 301476 199052 301486 199108
rect 302372 199052 303492 199108
rect 310594 199052 310604 199108
rect 310660 199052 324044 199108
rect 324100 199052 324110 199108
rect 310818 198940 310828 198996
rect 310884 198940 323260 198996
rect 323316 198940 323326 198996
rect 292226 198828 292236 198884
rect 292292 198828 308588 198884
rect 308644 198828 308654 198884
rect 311826 198828 311836 198884
rect 311892 198828 326844 198884
rect 326900 198828 326910 198884
rect 301186 198604 301196 198660
rect 301252 198604 326620 198660
rect 326676 198604 326686 198660
rect 269864 198268 272412 198324
rect 272468 198268 272478 198324
rect 324146 198268 324156 198324
rect 324212 198268 324380 198324
rect 324436 198268 324446 198324
rect 337250 198268 337260 198324
rect 337316 198268 337708 198324
rect 337764 198268 337774 198324
rect 332658 198156 332668 198212
rect 332724 198156 333900 198212
rect 333956 198156 333966 198212
rect 326946 198044 326956 198100
rect 327012 198044 336140 198100
rect 336196 198044 336206 198100
rect 305666 197820 305676 197876
rect 305732 197820 329980 197876
rect 330036 197820 330046 197876
rect 276322 197708 276332 197764
rect 276388 197708 321804 197764
rect 321860 197708 321870 197764
rect 323362 197708 323372 197764
rect 323428 197708 339164 197764
rect 339220 197708 339230 197764
rect 289650 197596 289660 197652
rect 289716 197596 339388 197652
rect 339444 197596 339454 197652
rect 324940 197428 324996 197512
rect 332612 197428 332668 197540
rect 332724 197484 332734 197540
rect 340060 197428 340116 197960
rect 271506 197372 271516 197428
rect 271572 197372 272300 197428
rect 272356 197372 272366 197428
rect 272738 197372 272748 197428
rect 272804 197372 273420 197428
rect 273476 197372 273486 197428
rect 324940 197372 332668 197428
rect 336130 197372 336140 197428
rect 336196 197372 340116 197428
rect 339378 197260 339388 197316
rect 339444 197260 340060 197316
rect 340116 197260 340126 197316
rect 339490 197148 339500 197204
rect 339556 197148 340620 197204
rect 340676 197148 340686 197204
rect 269490 195356 269500 195412
rect 269556 195356 269566 195412
rect 324370 195132 324380 195188
rect 324436 195132 324446 195188
rect 324380 194600 324436 195132
rect 269864 192444 272188 192500
rect 272244 192444 272254 192500
rect -960 192052 480 192248
rect 324706 192220 324716 192276
rect 324772 192220 324782 192276
rect -960 192024 31052 192052
rect 392 191996 31052 192024
rect 31108 191996 31118 192052
rect 324716 191716 324772 192220
rect 595560 192164 597000 192360
rect 590370 192108 590380 192164
rect 590436 192136 597000 192164
rect 590436 192108 595672 192136
rect 324716 191688 324968 191716
rect 324744 191660 324996 191688
rect 324940 191604 324996 191660
rect 324940 191548 328524 191604
rect 328580 191548 328590 191604
rect 335346 191548 335356 191604
rect 335412 191548 336028 191604
rect 336084 191548 336094 191604
rect 336018 191436 336028 191492
rect 336084 191436 337036 191492
rect 337092 191436 340088 191492
rect 271394 190652 271404 190708
rect 271460 190652 272412 190708
rect 272468 190652 272478 190708
rect 272850 190652 272860 190708
rect 272916 190652 272972 190708
rect 273028 190652 273038 190708
rect 330754 189756 330764 189812
rect 330820 189756 334796 189812
rect 334852 189756 334862 189812
rect 335906 189756 335916 189812
rect 335972 189756 337932 189812
rect 337988 189756 337998 189812
rect 269864 189532 272972 189588
rect 273028 189532 273038 189588
rect 329074 188972 329084 189028
rect 329140 188972 338940 189028
rect 338996 188972 339006 189028
rect 324940 188860 327628 188916
rect 327684 188860 327852 188916
rect 327908 188860 327918 188916
rect 324940 188776 324996 188860
rect 327058 188076 327068 188132
rect 327124 188076 328412 188132
rect 328468 188076 328478 188132
rect 334114 188076 334124 188132
rect 334180 188076 334460 188132
rect 334516 188076 334526 188132
rect 269864 186620 272524 186676
rect 272580 186620 272590 186676
rect 272402 186396 272412 186452
rect 272468 186396 272636 186452
rect 272692 186396 272702 186452
rect 327394 186396 327404 186452
rect 327460 186396 328636 186452
rect 328692 186396 328702 186452
rect 272962 185948 272972 186004
rect 273028 185948 277452 186004
rect 277508 185948 277518 186004
rect 324940 185332 324996 185864
rect 324940 185276 327404 185332
rect 327460 185276 327470 185332
rect 334114 184940 334124 184996
rect 334180 184940 340088 184996
rect 269864 183708 273196 183764
rect 273252 183708 273262 183764
rect 337362 183708 337372 183764
rect 337428 183708 340620 183764
rect 340676 183708 340686 183764
rect 324940 183036 333452 183092
rect 333508 183036 333518 183092
rect 324940 182952 324996 183036
rect 337362 182252 337372 182308
rect 337428 182252 338044 182308
rect 338100 182252 338110 182308
rect 336018 181356 336028 181412
rect 336084 181356 337148 181412
rect 337204 181356 339276 181412
rect 339332 181356 339342 181412
rect 269864 180796 272748 180852
rect 272804 180796 272814 180852
rect 324940 180124 336028 180180
rect 336084 180124 336094 180180
rect 324940 180040 324996 180124
rect 337250 179676 337260 179732
rect 337316 179676 337820 179732
rect 337876 179676 337886 179732
rect 595560 178948 597000 179144
rect 590370 178892 590380 178948
rect 590436 178920 597000 178948
rect 590436 178892 595672 178920
rect 273634 178444 273644 178500
rect 273700 178444 275996 178500
rect 276052 178444 276062 178500
rect 333890 178444 333900 178500
rect 333956 178444 340088 178500
rect -960 178052 480 178136
rect -960 177996 4284 178052
rect 4340 177996 4350 178052
rect 336018 177996 336028 178052
rect 336084 177996 337372 178052
rect 337428 177996 338380 178052
rect 338436 177996 338446 178052
rect -960 177912 480 177996
rect 269864 177884 272636 177940
rect 272692 177884 272702 177940
rect 324940 177044 324996 177128
rect 324940 176988 336028 177044
rect 336084 176988 336094 177044
rect 271842 176316 271852 176372
rect 271908 176316 273420 176372
rect 273476 176316 273486 176372
rect 269864 174972 273196 175028
rect 273252 174972 273262 175028
rect 324940 174636 328636 174692
rect 328692 174636 336028 174692
rect 336084 174636 336094 174692
rect 324940 174216 324996 174636
rect 269864 172060 273980 172116
rect 274036 172060 274046 172116
rect 339154 171948 339164 172004
rect 339220 171948 340088 172004
rect 324940 171220 324996 171304
rect 324940 171164 336140 171220
rect 336196 171164 336206 171220
rect 269864 169148 273084 169204
rect 273140 169148 273150 169204
rect 324940 168308 324996 168392
rect 324940 168252 336028 168308
rect 336084 168252 337036 168308
rect 337092 168252 337102 168308
rect 269864 166236 272860 166292
rect 272916 166236 272926 166292
rect 324940 166012 327628 166068
rect 327684 166012 327694 166068
rect 324940 165480 324996 166012
rect 595560 165704 597000 165928
rect 337586 165452 337596 165508
rect 337652 165452 340088 165508
rect -960 163828 480 164024
rect -960 163800 39452 163828
rect 392 163772 39452 163800
rect 39508 163772 39518 163828
rect 269864 163324 272748 163380
rect 272804 163324 272814 163380
rect 324940 161924 324996 162568
rect 324940 161868 327628 161924
rect 327684 161868 327694 161924
rect 339266 161084 339276 161140
rect 339332 161084 422604 161140
rect 422660 161084 422670 161140
rect 338370 160972 338380 161028
rect 338436 160972 422828 161028
rect 422884 160972 422894 161028
rect 467842 160860 467852 160916
rect 467908 160860 587132 160916
rect 587188 160860 587198 160916
rect 271730 160636 271740 160692
rect 271796 160636 590380 160692
rect 590436 160636 590446 160692
rect 284946 160524 284956 160580
rect 285012 160524 286188 160580
rect 286244 160524 286254 160580
rect 286412 160524 590716 160580
rect 590772 160524 590782 160580
rect 286412 160468 286468 160524
rect 269864 160412 275660 160468
rect 275716 160412 275726 160468
rect 280242 160412 280252 160468
rect 280308 160412 286468 160468
rect 290612 160412 523292 160468
rect 523348 160412 523358 160468
rect 290612 160356 290668 160412
rect 279906 160300 279916 160356
rect 279972 160300 290668 160356
rect 297490 160300 297500 160356
rect 297556 160300 298060 160356
rect 298116 160300 298126 160356
rect 335234 160300 335244 160356
rect 335300 160300 491932 160356
rect 491988 160300 491998 160356
rect 307682 160188 307692 160244
rect 307748 160188 325948 160244
rect 326004 160188 326014 160244
rect 338930 160188 338940 160244
rect 338996 160188 506716 160244
rect 506772 160188 506782 160244
rect 304098 160076 304108 160132
rect 304164 160076 326060 160132
rect 326116 160076 326126 160132
rect 330418 160076 330428 160132
rect 330484 160076 543676 160132
rect 543732 160076 543742 160132
rect 330642 159964 330652 160020
rect 330708 159964 351148 160020
rect 351204 159964 351214 160020
rect 422566 159964 422604 160020
rect 422660 159964 422670 160020
rect 422790 159964 422828 160020
rect 422884 159964 422894 160020
rect 467814 159964 467852 160020
rect 467908 159964 467918 160020
rect 591238 159628 591276 159684
rect 591332 159628 591342 159684
rect 335122 159516 335132 159572
rect 335188 159516 358876 159572
rect 358932 159516 358942 159572
rect 283266 159404 283276 159460
rect 283332 159404 591164 159460
rect 591220 159404 591230 159460
rect 293234 159292 293244 159348
rect 293300 159292 590940 159348
rect 590996 159292 591006 159348
rect 311266 159180 311276 159236
rect 311332 159180 324492 159236
rect 324548 159180 324558 159236
rect 357858 159180 357868 159236
rect 357924 159180 590380 159236
rect 590436 159180 590446 159236
rect 335570 159068 335580 159124
rect 335636 159068 528892 159124
rect 528948 159068 528958 159124
rect 332098 158956 332108 159012
rect 332164 158956 521500 159012
rect 521556 158956 521566 159012
rect 341506 158844 341516 158900
rect 341572 158844 575372 158900
rect 575428 158844 575438 158900
rect 324258 158732 324268 158788
rect 324324 158732 578172 158788
rect 578228 158732 578238 158788
rect 281474 158620 281484 158676
rect 281540 158620 590604 158676
rect 590660 158620 590670 158676
rect 327506 158508 327516 158564
rect 327572 158508 373660 158564
rect 373716 158508 373726 158564
rect 284610 157836 284620 157892
rect 284676 157836 291564 157892
rect 291620 157836 291630 157892
rect 309474 157836 309484 157892
rect 309540 157836 326284 157892
rect 326340 157836 326350 157892
rect 338706 157836 338716 157892
rect 338772 157836 344092 157892
rect 344148 157836 344158 157892
rect 283602 157724 283612 157780
rect 283668 157724 293356 157780
rect 293412 157724 293422 157780
rect 302306 157724 302316 157780
rect 302372 157724 324268 157780
rect 324324 157724 324334 157780
rect 338482 157724 338492 157780
rect 338548 157724 447580 157780
rect 447636 157724 447646 157780
rect 305890 157612 305900 157668
rect 305956 157612 324604 157668
rect 324660 157612 324670 157668
rect 331986 157612 331996 157668
rect 332052 157612 381052 157668
rect 381108 157612 381118 157668
rect 558422 157612 558460 157668
rect 558516 157612 558526 157668
rect 269864 157500 270620 157556
rect 270676 157500 270686 157556
rect 283378 157500 283388 157556
rect 283444 157500 296940 157556
rect 296996 157500 297006 157556
rect 316642 157500 316652 157556
rect 316708 157500 333116 157556
rect 333172 157500 333182 157556
rect 420802 157500 420812 157556
rect 420868 157500 454972 157556
rect 455028 157500 455038 157556
rect 457762 157500 457772 157556
rect 457828 157500 477148 157556
rect 477204 157500 477214 157556
rect 514098 157500 514108 157556
rect 514164 157500 514202 157556
rect 320226 157388 320236 157444
rect 320292 157388 333004 157444
rect 333060 157388 574812 157444
rect 574868 157388 574878 157444
rect 283714 157276 283724 157332
rect 283780 157276 295148 157332
rect 295204 157276 295214 157332
rect 323810 157276 323820 157332
rect 323876 157276 334012 157332
rect 334068 157276 574588 157332
rect 574644 157276 574654 157332
rect 300514 157164 300524 157220
rect 300580 157164 326508 157220
rect 326564 157164 326574 157220
rect 332658 157164 332668 157220
rect 332724 157164 333900 157220
rect 333956 157164 576492 157220
rect 576548 157164 576558 157220
rect 322018 157052 322028 157108
rect 322084 157052 333788 157108
rect 333844 157052 576268 157108
rect 576324 157052 576334 157108
rect 324482 156940 324492 156996
rect 324548 156940 333900 156996
rect 333956 156940 333966 156996
rect 335794 156940 335804 156996
rect 335860 156940 499324 156996
rect 499380 156940 499390 156996
rect 332210 156828 332220 156884
rect 332276 156828 366268 156884
rect 366324 156828 366334 156884
rect 318434 156716 318444 156772
rect 318500 156716 332668 156772
rect 332724 156716 332734 156772
rect 333554 156380 333564 156436
rect 333620 156380 335356 156436
rect 335412 156380 335422 156436
rect 333106 156268 333116 156324
rect 333172 156268 333676 156324
rect 333732 156268 333742 156324
rect 457986 156268 457996 156324
rect 458052 156268 462364 156324
rect 462420 156268 462430 156324
rect 328850 156156 328860 156212
rect 328916 156156 573244 156212
rect 573300 156156 573310 156212
rect 313058 156044 313068 156100
rect 313124 156044 333228 156100
rect 333284 156044 333294 156100
rect 337362 156044 337372 156100
rect 337428 156044 551068 156100
rect 551124 156044 551134 156100
rect 314850 155932 314860 155988
rect 314916 155932 333564 155988
rect 333620 155932 333630 155988
rect 340274 155932 340284 155988
rect 340340 155932 536284 155988
rect 536340 155932 536350 155988
rect 328066 155820 328076 155876
rect 328132 155820 484540 155876
rect 484596 155820 484606 155876
rect 278674 155708 278684 155764
rect 278740 155708 514892 155764
rect 514948 155708 514958 155764
rect 337250 155596 337260 155652
rect 337316 155596 578508 155652
rect 578564 155596 578574 155652
rect 285394 155484 285404 155540
rect 285460 155484 548044 155540
rect 548100 155484 548110 155540
rect 295138 155372 295148 155428
rect 295204 155372 574028 155428
rect 574084 155372 574094 155428
rect 341170 155260 341180 155316
rect 341236 155260 341516 155316
rect 341572 155260 341582 155316
rect 349412 155260 388444 155316
rect 388500 155260 388510 155316
rect 469522 155260 469532 155316
rect 469588 155260 585452 155316
rect 585508 155260 585518 155316
rect 349412 155204 349468 155260
rect 338594 155148 338604 155204
rect 338660 155148 349468 155204
rect 269864 154588 275772 154644
rect 275828 154588 275838 154644
rect 293122 154476 293132 154532
rect 293188 154476 591276 154532
rect 591332 154476 591342 154532
rect 334226 154364 334236 154420
rect 334292 154364 425404 154420
rect 425460 154364 425470 154420
rect 285282 154028 285292 154084
rect 285348 154028 516908 154084
rect 516964 154028 516974 154084
rect 293794 153916 293804 153972
rect 293860 153916 535052 153972
rect 535108 153916 535118 153972
rect 325378 153804 325388 153860
rect 325444 153804 574700 153860
rect 574756 153804 574766 153860
rect 281586 153692 281596 153748
rect 281652 153692 590828 153748
rect 590884 153692 590894 153748
rect 458210 153020 458220 153076
rect 458276 153020 574476 153076
rect 574532 153020 574542 153076
rect 333666 152908 333676 152964
rect 333732 152908 336028 152964
rect 336084 152908 479052 152964
rect 479108 152908 479118 152964
rect 338818 152796 338828 152852
rect 338884 152796 580636 152852
rect 580692 152796 580702 152852
rect 340386 152684 340396 152740
rect 340452 152684 410620 152740
rect 410676 152684 410686 152740
rect 590034 152684 590044 152740
rect 590100 152712 595672 152740
rect 590100 152684 597000 152712
rect 335682 152572 335692 152628
rect 335748 152572 403228 152628
rect 403284 152572 403294 152628
rect 457874 152572 457884 152628
rect 457940 152572 565852 152628
rect 565908 152572 565918 152628
rect 334786 152460 334796 152516
rect 334852 152460 395836 152516
rect 395892 152460 395902 152516
rect 466498 152460 466508 152516
rect 466564 152460 585564 152516
rect 585620 152460 585630 152516
rect 595560 152488 597000 152684
rect 284386 152348 284396 152404
rect 284452 152348 510636 152404
rect 510692 152348 510702 152404
rect 326722 152236 326732 152292
rect 326788 152236 562156 152292
rect 562212 152236 562222 152292
rect 333554 152124 333564 152180
rect 333620 152124 574700 152180
rect 574756 152124 574766 152180
rect 292226 152012 292236 152068
rect 292292 152012 574924 152068
rect 574980 152012 574990 152068
rect 269864 151676 273868 151732
rect 273924 151676 273934 151732
rect 336578 151228 336588 151284
rect 336644 151228 486892 151284
rect 486948 151228 486958 151284
rect 331650 151116 331660 151172
rect 331716 151116 432796 151172
rect 432852 151116 432862 151172
rect 324930 151004 324940 151060
rect 324996 151004 565292 151060
rect 565348 151004 565358 151060
rect 333218 150892 333228 150948
rect 333284 150892 576604 150948
rect 576660 150892 576670 150948
rect 328514 150780 328524 150836
rect 328580 150780 578396 150836
rect 578452 150780 578462 150836
rect 275314 150668 275324 150724
rect 275380 150668 527660 150724
rect 527716 150668 527726 150724
rect 278786 150556 278796 150612
rect 278852 150556 532364 150612
rect 532420 150556 532430 150612
rect 277106 150444 277116 150500
rect 277172 150444 530796 150500
rect 530852 150444 530862 150500
rect 275426 150332 275436 150388
rect 275492 150332 529228 150388
rect 529284 150332 529294 150388
rect 392 149912 7532 149940
rect -960 149884 7532 149912
rect 7588 149884 7598 149940
rect -960 149688 480 149884
rect 462914 149660 462924 149716
rect 462980 149660 499436 149716
rect 499492 149660 499502 149716
rect 337474 149548 337484 149604
rect 337540 149548 483756 149604
rect 483812 149548 483822 149604
rect 329746 149436 329756 149492
rect 329812 149436 469756 149492
rect 469812 149436 469822 149492
rect 338818 149324 338828 149380
rect 338884 149324 418012 149380
rect 418068 149324 418078 149380
rect 272066 148988 272076 149044
rect 272132 148988 512428 149044
rect 512484 148988 512494 149044
rect 278674 148876 278684 148932
rect 278740 148876 524524 148932
rect 524580 148876 524590 148932
rect 269864 148764 272524 148820
rect 272580 148764 272590 148820
rect 326834 148764 326844 148820
rect 326900 148764 575148 148820
rect 575204 148764 575214 148820
rect 282034 148652 282044 148708
rect 282100 148652 568428 148708
rect 568484 148652 568494 148708
rect 463698 148092 463708 148148
rect 463764 148092 575036 148148
rect 575092 148092 575102 148148
rect 465378 147980 465388 148036
rect 465444 147980 578396 148036
rect 578452 147980 578462 148036
rect 336018 147868 336028 147924
rect 336084 147868 337596 147924
rect 337652 147868 494732 147924
rect 494788 147868 494798 147924
rect 341394 147756 341404 147812
rect 341460 147756 422716 147812
rect 422772 147756 422782 147812
rect 333890 147644 333900 147700
rect 333956 147644 575260 147700
rect 575316 147644 575326 147700
rect 274866 147532 274876 147588
rect 274932 147532 526092 147588
rect 526148 147532 526158 147588
rect 283826 147420 283836 147476
rect 283892 147420 552748 147476
rect 552804 147420 552814 147476
rect 288866 147308 288876 147364
rect 288932 147308 559020 147364
rect 559076 147308 559086 147364
rect 285506 147196 285516 147252
rect 285572 147196 555884 147252
rect 555940 147196 555950 147252
rect 280466 147084 280476 147140
rect 280532 147084 551180 147140
rect 551236 147084 551246 147140
rect 280354 146972 280364 147028
rect 280420 146972 557452 147028
rect 557508 146972 557518 147028
rect 466386 146300 466396 146356
rect 466452 146300 488460 146356
rect 488516 146300 488526 146356
rect 462802 146188 462812 146244
rect 462868 146188 493164 146244
rect 493220 146188 493230 146244
rect 273634 146076 273644 146132
rect 273700 146076 327628 146132
rect 327684 146076 505596 146132
rect 505652 146076 505662 146132
rect 333666 145964 333676 146020
rect 333732 145964 579628 146020
rect 579684 145964 579694 146020
rect 269864 145852 272636 145908
rect 272692 145852 273644 145908
rect 273700 145852 273710 145908
rect 280802 145740 280812 145796
rect 280868 145740 538636 145796
rect 538692 145740 538702 145796
rect 281698 145628 281708 145684
rect 281764 145628 540204 145684
rect 540260 145628 540270 145684
rect 282594 145516 282604 145572
rect 282660 145516 541772 145572
rect 541828 145516 541838 145572
rect 283490 145404 283500 145460
rect 283556 145404 543340 145460
rect 543396 145404 543406 145460
rect 293906 145292 293916 145348
rect 293972 145292 566860 145348
rect 566916 145292 566926 145348
rect 341282 145180 341292 145236
rect 341348 145180 422380 145236
rect 422436 145180 422446 145236
rect 270274 145068 270284 145124
rect 270340 145068 519820 145124
rect 519876 145068 519886 145124
rect 458434 144508 458444 144564
rect 458500 144508 521388 144564
rect 521444 144508 521454 144564
rect 325826 144396 325836 144452
rect 325892 144396 420812 144452
rect 420868 144396 420878 144452
rect 332658 144284 332668 144340
rect 332724 144284 336028 144340
rect 336084 144284 336094 144340
rect 324146 144060 324156 144116
rect 324212 144060 327628 144116
rect 327684 144060 327694 144116
rect 422706 144060 422716 144116
rect 422772 144060 423276 144116
rect 423332 144060 423342 144116
rect 512418 144060 512428 144116
rect 512484 144060 522956 144116
rect 523012 144060 523022 144116
rect 337026 143948 337036 144004
rect 337092 143948 337484 144004
rect 337540 143948 504140 144004
rect 504196 143948 504206 144004
rect 505586 143948 505596 144004
rect 505652 143948 516684 144004
rect 516740 143948 516750 144004
rect 516898 143948 516908 144004
rect 516964 143948 520156 144004
rect 520212 143948 520222 144004
rect 523282 143948 523292 144004
rect 523348 143948 537068 144004
rect 537124 143948 537134 144004
rect 422370 143836 422380 143892
rect 422436 143836 466508 143892
rect 466564 143836 466574 143892
rect 514882 143836 514892 143892
rect 514948 143836 533932 143892
rect 533988 143836 533998 143892
rect 535042 143836 535052 143892
rect 535108 143836 560588 143892
rect 560644 143836 560654 143892
rect 422594 143724 422604 143780
rect 422660 143724 423164 143780
rect 423220 143724 423230 143780
rect 423378 143724 423388 143780
rect 423444 143724 469532 143780
rect 469588 143724 469598 143780
rect 502292 143724 515116 143780
rect 515172 143724 515182 143780
rect 519932 143724 544908 143780
rect 544964 143724 544974 143780
rect 502292 143668 502348 143724
rect 519932 143668 519988 143724
rect 269836 143612 270620 143668
rect 270676 143612 328524 143668
rect 328580 143612 502348 143668
rect 510626 143612 510636 143668
rect 510692 143612 519988 143668
rect 520146 143612 520156 143668
rect 520212 143612 546476 143668
rect 546532 143612 546542 143668
rect 269836 142968 269892 143612
rect 422818 143500 422828 143556
rect 422884 143500 471212 143556
rect 471268 143500 471278 143556
rect 507490 143500 507500 143556
rect 507556 143500 563724 143556
rect 563780 143500 563790 143556
rect 273186 143388 273196 143444
rect 273252 143388 273420 143444
rect 273476 143388 510412 143444
rect 510468 143388 510478 143444
rect 422258 143276 422268 143332
rect 422324 143276 467852 143332
rect 467908 143276 467918 143332
rect 510738 143276 510748 143332
rect 510804 143276 535500 143332
rect 535556 143276 535566 143332
rect 423154 143164 423164 143220
rect 423220 143164 472108 143220
rect 472164 143164 472174 143220
rect 472882 143164 472892 143220
rect 472948 143164 576492 143220
rect 576548 143164 576558 143220
rect 468626 143052 468636 143108
rect 468692 143052 578284 143108
rect 578340 143052 578350 143108
rect 501666 142940 501676 142996
rect 501732 142940 554316 142996
rect 554372 142940 554382 142996
rect 458322 142828 458332 142884
rect 458388 142828 474348 142884
rect 474404 142828 474414 142884
rect 489990 142828 490028 142884
rect 490084 142828 490094 142884
rect 497830 142828 497868 142884
rect 497924 142828 497934 142884
rect 505670 142828 505708 142884
rect 505764 142828 505774 142884
rect 507238 142828 507276 142884
rect 507332 142828 507342 142884
rect 508806 142828 508844 142884
rect 508900 142828 508910 142884
rect 511942 142828 511980 142884
rect 512036 142828 512046 142884
rect 513510 142828 513548 142884
rect 513604 142828 513614 142884
rect 279010 142716 279020 142772
rect 279076 142716 510748 142772
rect 510804 142716 510814 142772
rect 318546 142604 318556 142660
rect 318612 142604 330988 142660
rect 331044 142604 335020 142660
rect 335076 142604 335086 142660
rect 340610 142604 340620 142660
rect 340676 142604 463708 142660
rect 463764 142604 463774 142660
rect 323362 142492 323372 142548
rect 323428 142492 336028 142548
rect 336084 142492 336094 142548
rect 318322 142380 318332 142436
rect 318388 142380 336588 142436
rect 336644 142380 336654 142436
rect 309922 142268 309932 142324
rect 309988 142268 328860 142324
rect 328916 142268 335916 142324
rect 335972 142268 335982 142324
rect 338930 142268 338940 142324
rect 338996 142268 578732 142324
rect 578788 142268 578798 142324
rect 270386 142156 270396 142212
rect 270452 142156 518252 142212
rect 518308 142156 518318 142212
rect 325378 142044 325388 142100
rect 325444 142044 578284 142100
rect 578340 142044 578350 142100
rect 282146 141932 282156 141988
rect 282212 141932 549612 141988
rect 549668 141932 549678 141988
rect 468514 141708 468524 141764
rect 468580 141708 479612 141764
rect 479668 141708 479678 141764
rect 455252 141596 475916 141652
rect 475972 141596 475982 141652
rect 455252 141540 455308 141596
rect 425842 141484 425852 141540
rect 425908 141484 455308 141540
rect 472444 141484 472836 141540
rect 472444 141428 472500 141484
rect 463026 141372 463036 141428
rect 463092 141372 472500 141428
rect 472780 141316 472836 141484
rect 473732 141484 485548 141540
rect 473732 141428 473788 141484
rect 473116 141372 473788 141428
rect 485492 141428 485548 141484
rect 485492 141372 491596 141428
rect 491652 141372 491662 141428
rect 473116 141316 473172 141372
rect 466274 141260 466284 141316
rect 466340 141260 468524 141316
rect 468580 141260 468590 141316
rect 472780 141260 473172 141316
rect 479602 141260 479612 141316
rect 479668 141260 502572 141316
rect 502628 141260 502638 141316
rect 466610 141148 466620 141204
rect 466676 141148 485324 141204
rect 485380 141148 485390 141204
rect 295362 141036 295372 141092
rect 295428 141036 507500 141092
rect 507556 141036 507566 141092
rect 330194 140924 330204 140980
rect 330260 140924 465388 140980
rect 465444 140924 465454 140980
rect 329970 140812 329980 140868
rect 330036 140812 576828 140868
rect 576884 140812 576894 140868
rect 324034 140700 324044 140756
rect 324100 140700 575596 140756
rect 575652 140700 575662 140756
rect 325154 140588 325164 140644
rect 325220 140588 577948 140644
rect 578004 140588 578014 140644
rect 323250 140476 323260 140532
rect 323316 140476 576716 140532
rect 576772 140476 576782 140532
rect 293682 140364 293692 140420
rect 293748 140364 576940 140420
rect 576996 140364 577006 140420
rect 290434 140252 290444 140308
rect 290500 140252 581308 140308
rect 581364 140252 581374 140308
rect 269864 140028 336140 140084
rect 336196 140028 336206 140084
rect 480582 139692 480620 139748
rect 480676 139692 480686 139748
rect 466162 139580 466172 139636
rect 466228 139580 477484 139636
rect 477540 139580 477550 139636
rect 482150 139580 482188 139636
rect 482244 139580 482254 139636
rect 467058 139468 467068 139524
rect 467124 139468 501004 139524
rect 501060 139468 501070 139524
rect 501638 139468 501676 139524
rect 501732 139468 501742 139524
rect 595560 139412 597000 139496
rect 590146 139356 590156 139412
rect 590212 139356 597000 139412
rect 337652 139244 496300 139300
rect 496356 139244 496366 139300
rect 595560 139272 597000 139356
rect 311602 139132 311612 139188
rect 311668 139132 337260 139188
rect 337316 139132 337326 139188
rect 337652 139076 337708 139244
rect 273074 139020 273084 139076
rect 273140 139020 332668 139076
rect 332724 139020 332734 139076
rect 332892 139020 337708 139076
rect 338482 139020 338492 139076
rect 338548 139020 578172 139076
rect 578228 139020 578238 139076
rect 332892 138964 332948 139020
rect 314132 138908 328972 138964
rect 329028 138908 332948 138964
rect 333554 138908 333564 138964
rect 333620 138908 576380 138964
rect 576436 138908 576446 138964
rect 314132 138852 314188 138908
rect 308242 138796 308252 138852
rect 308308 138796 314188 138852
rect 330530 138796 330540 138852
rect 330596 138796 578060 138852
rect 578116 138796 578126 138852
rect 325266 138684 325276 138740
rect 325332 138684 575484 138740
rect 575540 138684 575550 138740
rect 323922 138572 323932 138628
rect 323988 138572 578620 138628
rect 578676 138572 578686 138628
rect 290546 138460 290556 138516
rect 290612 138460 501676 138516
rect 501732 138460 501742 138516
rect 270946 137676 270956 137732
rect 271012 137676 458444 137732
rect 458500 137676 458510 137732
rect 329858 137564 329868 137620
rect 329924 137564 457996 137620
rect 458052 137564 458062 137620
rect 339042 137452 339052 137508
rect 339108 137452 458220 137508
rect 458276 137452 458286 137508
rect 269864 137116 272188 137172
rect 272244 137116 272254 137172
rect 333442 136892 333452 136948
rect 333508 136892 422380 136948
rect 422436 136892 422446 136948
rect 330418 135996 330428 136052
rect 330484 135996 457996 136052
rect 458052 135996 458062 136052
rect 331762 135884 331772 135940
rect 331828 135884 457772 135940
rect 457828 135884 457838 135940
rect -960 135604 480 135800
rect 340162 135772 340172 135828
rect 340228 135772 440188 135828
rect 440244 135772 440254 135828
rect 422370 135660 422380 135716
rect 422436 135660 422604 135716
rect 422660 135660 458332 135716
rect 458388 135660 458398 135716
rect -960 135576 29372 135604
rect 392 135548 29372 135576
rect 29428 135548 29438 135604
rect 339938 135436 339948 135492
rect 340004 135436 459396 135492
rect 574952 135436 577948 135492
rect 578004 135436 578014 135492
rect 459340 135380 460040 135436
rect 329074 134316 329084 134372
rect 329140 134316 332668 134372
rect 332724 134316 333340 134372
rect 333396 134316 333406 134372
rect 336802 134316 336812 134372
rect 336868 134316 336924 134372
rect 336980 134316 336990 134372
rect 269864 134204 273196 134260
rect 273252 134204 273262 134260
rect 327954 134092 327964 134148
rect 328020 134092 457884 134148
rect 457940 134092 457950 134148
rect 574578 133980 574588 134036
rect 574644 133980 574654 134036
rect 574588 133448 574644 133980
rect 330642 132076 330652 132132
rect 330708 132076 459396 132132
rect 459340 132020 460040 132076
rect 575026 131852 575036 131908
rect 575092 131852 575596 131908
rect 575652 131852 575662 131908
rect 574952 131404 576268 131460
rect 576324 131404 576334 131460
rect 269864 131292 273196 131348
rect 273252 131292 273262 131348
rect 341506 130956 341516 131012
rect 341572 130956 421708 131012
rect 421764 130956 422268 131012
rect 422324 130956 422334 131012
rect 574802 129948 574812 130004
rect 574868 129948 574878 130004
rect 574812 129416 574868 129948
rect 335682 128716 335692 128772
rect 335748 128716 459396 128772
rect 459340 128660 460040 128716
rect 287746 128604 287756 128660
rect 287812 128604 337036 128660
rect 337092 128604 337102 128660
rect 281810 128492 281820 128548
rect 281876 128492 386204 128548
rect 386260 128492 386270 128548
rect 269864 128380 280140 128436
rect 280196 128380 280206 128436
rect 336802 127596 336812 127652
rect 336868 127596 337148 127652
rect 337204 127596 337214 127652
rect 574952 127372 576492 127428
rect 576548 127372 576558 127428
rect 595560 126056 597000 126280
rect 269864 125468 272972 125524
rect 273028 125468 273038 125524
rect 332546 125356 332556 125412
rect 332612 125356 459396 125412
rect 574952 125356 579628 125412
rect 579684 125356 579694 125412
rect 459340 125300 460040 125356
rect 274754 125132 274764 125188
rect 274820 125132 387772 125188
rect 387828 125132 387838 125188
rect 574952 123340 576380 123396
rect 576436 123340 576446 123396
rect 323474 122668 323484 122724
rect 323540 122668 324156 122724
rect 324212 122668 423276 122724
rect 423332 122668 423342 122724
rect 421820 122612 421876 122668
rect 269864 122556 287756 122612
rect 287812 122556 287822 122612
rect 421810 122556 421820 122612
rect 421876 122556 421886 122612
rect 335234 121996 335244 122052
rect 335300 121996 459396 122052
rect 459340 121940 460040 121996
rect 272850 121772 272860 121828
rect 272916 121772 333900 121828
rect 333956 121772 333966 121828
rect -960 121492 480 121688
rect -960 121464 36092 121492
rect 392 121436 36092 121464
rect 36148 121436 36158 121492
rect 574952 121324 576604 121380
rect 576660 121324 576670 121380
rect 269864 119644 272860 119700
rect 272916 119644 272926 119700
rect 574952 119308 575260 119364
rect 575316 119308 575326 119364
rect 331874 118636 331884 118692
rect 331940 118636 459396 118692
rect 459340 118580 460040 118636
rect 326722 117516 326732 117572
rect 326788 117516 327404 117572
rect 327460 117516 327470 117572
rect 425058 117516 425068 117572
rect 425124 117516 425852 117572
rect 425908 117516 425918 117572
rect 574952 117292 575148 117348
rect 575204 117292 575214 117348
rect 269864 116732 304892 116788
rect 304948 116732 304958 116788
rect 326722 116732 326732 116788
rect 326788 116732 425068 116788
rect 425124 116732 425134 116788
rect 331762 115276 331772 115332
rect 331828 115276 459396 115332
rect 574952 115276 576716 115332
rect 576772 115276 576782 115332
rect 459340 115220 460040 115276
rect 269864 113820 306572 113876
rect 306628 113820 306638 113876
rect 574924 113820 575148 113876
rect 575204 113820 575214 113876
rect 269938 113484 269948 113540
rect 270004 113484 379820 113540
rect 379876 113484 379886 113540
rect 271618 113372 271628 113428
rect 271684 113372 411180 113428
rect 411236 113372 411246 113428
rect 574924 113288 574980 113820
rect 590818 113036 590828 113092
rect 590884 113064 595672 113092
rect 590884 113036 597000 113064
rect 595560 112840 597000 113036
rect 332098 111916 332108 111972
rect 332164 111916 459396 111972
rect 459340 111860 460040 111916
rect 574914 111804 574924 111860
rect 574980 111804 574990 111860
rect 574924 111272 574980 111804
rect 269864 110908 293132 110964
rect 293188 110908 293198 110964
rect 280018 110572 280028 110628
rect 280084 110572 395500 110628
rect 395556 110572 395566 110628
rect 278338 110460 278348 110516
rect 278404 110460 398636 110516
rect 398692 110460 398702 110516
rect 335794 110348 335804 110404
rect 335860 110348 458108 110404
rect 458164 110348 458174 110404
rect 278114 110236 278124 110292
rect 278180 110236 401772 110292
rect 401828 110236 401838 110292
rect 328402 110124 328412 110180
rect 328468 110124 457884 110180
rect 457940 110124 457950 110180
rect 274866 110012 274876 110068
rect 274932 110012 409612 110068
rect 409668 110012 409678 110068
rect 574952 109228 578284 109284
rect 578340 109228 578350 109284
rect 269602 108668 269612 108724
rect 269668 108668 384524 108724
rect 384580 108668 384590 108724
rect 327282 108556 327292 108612
rect 327348 108556 459396 108612
rect 459340 108500 460040 108556
rect 279682 108444 279692 108500
rect 279748 108444 404908 108500
rect 404964 108444 404974 108500
rect 271282 108332 271292 108388
rect 271348 108332 400204 108388
rect 400260 108332 400270 108388
rect 269864 107996 308252 108052
rect 308308 107996 308318 108052
rect -960 107380 480 107576
rect 574690 107436 574700 107492
rect 574756 107436 574766 107492
rect -960 107352 14252 107380
rect 392 107324 14252 107352
rect 14308 107324 14318 107380
rect 574700 107240 574756 107436
rect 334114 106988 334124 107044
rect 334180 106988 421820 107044
rect 421876 106988 421886 107044
rect 285842 106876 285852 106932
rect 285908 106876 373548 106932
rect 373604 106876 373614 106932
rect 276434 106764 276444 106820
rect 276500 106764 375116 106820
rect 375172 106764 375182 106820
rect 335458 106652 335468 106708
rect 335524 106652 457772 106708
rect 457828 106652 457838 106708
rect 269938 105308 269948 105364
rect 270004 105308 407484 105364
rect 407540 105308 407550 105364
rect 325714 105196 325724 105252
rect 325780 105196 459396 105252
rect 574952 105196 578172 105252
rect 578228 105196 578238 105252
rect 459340 105140 460040 105196
rect 269864 105084 323372 105140
rect 323428 105084 323438 105140
rect 270050 104972 270060 105028
rect 270116 104972 412188 105028
rect 412244 104972 412254 105028
rect 283042 104076 283052 104132
rect 283108 104076 378028 104132
rect 378084 104076 378094 104132
rect 413298 104076 413308 104132
rect 413364 104076 414092 104132
rect 414148 104076 414158 104132
rect 414978 104076 414988 104132
rect 415044 104076 415660 104132
rect 415716 104076 415726 104132
rect 278002 103964 278012 104020
rect 278068 103964 381388 104020
rect 381444 103964 381454 104020
rect 406662 103964 406700 104020
rect 406756 103964 406766 104020
rect 276770 103852 276780 103908
rect 276836 103852 383180 103908
rect 383236 103852 383246 103908
rect 403190 103852 403228 103908
rect 403284 103852 403294 103908
rect 278450 103740 278460 103796
rect 278516 103740 388668 103796
rect 388724 103740 388734 103796
rect 278226 103628 278236 103684
rect 278292 103628 390236 103684
rect 390292 103628 390302 103684
rect 279794 103516 279804 103572
rect 279860 103516 393372 103572
rect 393428 103516 393438 103572
rect 276546 103404 276556 103460
rect 276612 103404 391804 103460
rect 391860 103404 391870 103460
rect 274642 103292 274652 103348
rect 274708 103292 396508 103348
rect 396564 103292 396574 103348
rect 325042 103180 325052 103236
rect 325108 103180 376572 103236
rect 376628 103180 376638 103236
rect 574952 103180 576828 103236
rect 576884 103180 576894 103236
rect 269864 102172 280252 102228
rect 280308 102172 280318 102228
rect 329634 101836 329644 101892
rect 329700 101836 459396 101892
rect 459340 101780 460040 101836
rect 336914 101724 336924 101780
rect 336980 101724 458556 101780
rect 458612 101724 458622 101780
rect 574924 101724 575036 101780
rect 575092 101724 575102 101780
rect 332210 101612 332220 101668
rect 332276 101612 456988 101668
rect 457044 101612 457054 101668
rect 574924 101192 574980 101724
rect 334002 100156 334012 100212
rect 334068 100156 421708 100212
rect 421764 100156 421774 100212
rect 330530 100044 330540 100100
rect 330596 100044 458220 100100
rect 458276 100044 458286 100100
rect 330306 99932 330316 99988
rect 330372 99932 458444 99988
rect 458500 99932 458510 99988
rect 590706 99820 590716 99876
rect 590772 99848 595672 99876
rect 590772 99820 597000 99848
rect 595560 99624 597000 99820
rect 269864 99260 274988 99316
rect 275044 99260 275054 99316
rect 574952 99148 575372 99204
rect 575428 99148 575438 99204
rect 274642 99036 274652 99092
rect 274708 99036 336812 99092
rect 336868 99036 336878 99092
rect 337026 99036 337036 99092
rect 337092 99036 458556 99092
rect 458612 99036 458622 99092
rect 333442 98924 333452 98980
rect 333508 98924 458332 98980
rect 458388 98924 458398 98980
rect 330082 98812 330092 98868
rect 330148 98812 457772 98868
rect 457828 98812 457838 98868
rect 326722 98700 326732 98756
rect 326788 98700 457436 98756
rect 457492 98700 457502 98756
rect 325826 98588 325836 98644
rect 325892 98588 457548 98644
rect 457604 98588 457614 98644
rect 329858 98476 329868 98532
rect 329924 98476 459396 98532
rect 459340 98420 460040 98476
rect 295026 98364 295036 98420
rect 295092 98364 457660 98420
rect 457716 98364 457726 98420
rect 294802 98252 294812 98308
rect 294868 98252 457996 98308
rect 458052 98252 458062 98308
rect 456978 97580 456988 97636
rect 457044 97580 458444 97636
rect 458500 97580 458510 97636
rect 574952 97132 581308 97188
rect 581364 97132 581374 97188
rect 419944 97020 421820 97076
rect 421876 97020 424172 97076
rect 424228 97020 424238 97076
rect 269864 96348 318556 96404
rect 318612 96348 318622 96404
rect 457650 95116 457660 95172
rect 457716 95116 459396 95172
rect 574952 95116 576940 95172
rect 576996 95116 577006 95172
rect 459340 95060 460040 95116
rect 282146 93996 282156 94052
rect 282212 93996 366268 94052
rect 366324 93996 367052 94052
rect 367108 93996 367118 94052
rect 392 93464 10892 93492
rect -960 93436 10892 93464
rect 10948 93436 10958 93492
rect 269864 93436 280588 93492
rect 280644 93436 282156 93492
rect 282212 93436 282222 93492
rect -960 93240 480 93436
rect 574952 93100 575484 93156
rect 575540 93100 575550 93156
rect 419916 91588 419972 92120
rect 457426 91756 457436 91812
rect 457492 91756 459396 91812
rect 459340 91700 460040 91756
rect 273186 91532 273196 91588
rect 273252 91532 323484 91588
rect 323540 91532 323550 91588
rect 366258 91532 366268 91588
rect 366324 91532 369460 91588
rect 419916 91532 421708 91588
rect 421764 91532 427532 91588
rect 427588 91532 427598 91588
rect 369404 91476 370104 91532
rect 574952 91084 578844 91140
rect 578900 91084 578910 91140
rect 269864 90524 318332 90580
rect 318388 90524 318398 90580
rect 574924 89628 575036 89684
rect 575092 89628 575102 89684
rect 574924 89096 574980 89628
rect 458546 88396 458556 88452
rect 458612 88396 459396 88452
rect 459340 88340 460040 88396
rect 269864 87612 309932 87668
rect 309988 87612 309998 87668
rect 419944 87164 421820 87220
rect 421876 87164 421886 87220
rect 574952 87052 578508 87108
rect 578564 87052 578574 87108
rect 273298 86492 273308 86548
rect 273364 86492 326732 86548
rect 326788 86492 326798 86548
rect 595560 86408 597000 86632
rect 457538 85036 457548 85092
rect 457604 85036 459396 85092
rect 574952 85036 578732 85092
rect 578788 85036 578798 85092
rect 459340 84980 460040 85036
rect 276434 84812 276444 84868
rect 276500 84812 367052 84868
rect 367108 84812 367118 84868
rect 269864 84700 311612 84756
rect 311668 84700 311678 84756
rect 273410 83132 273420 83188
rect 273476 83132 332668 83188
rect 332724 83132 332734 83188
rect 574914 83020 574924 83076
rect 574980 83020 574990 83076
rect 419944 82236 425068 82292
rect 425124 82236 425134 82292
rect 269864 81788 274652 81844
rect 274708 81788 274718 81844
rect 458434 81676 458444 81732
rect 458500 81676 459396 81732
rect 459340 81620 460040 81676
rect 574802 81004 574812 81060
rect 574868 81004 574878 81060
rect -960 79156 480 79352
rect -960 79128 4284 79156
rect 392 79100 4284 79128
rect 4340 79100 4350 79156
rect 574952 78988 578396 79044
rect 578452 78988 578462 79044
rect 269864 78876 273420 78932
rect 273476 78876 273486 78932
rect 458546 78316 458556 78372
rect 458612 78316 459396 78372
rect 459340 78260 460040 78316
rect 419944 77308 420140 77364
rect 420196 77308 422604 77364
rect 422660 77308 422670 77364
rect 574952 76972 578060 77028
rect 578116 76972 578126 77028
rect 269864 75964 273084 76020
rect 273140 75964 273150 76020
rect 367042 74956 367052 75012
rect 367108 74956 369460 75012
rect 458322 74956 458332 75012
rect 458388 74956 459396 75012
rect 574690 74956 574700 75012
rect 574756 74956 574766 75012
rect 369404 74900 370104 74956
rect 459340 74900 460040 74956
rect 590594 73388 590604 73444
rect 590660 73416 595672 73444
rect 590660 73388 597000 73416
rect 595560 73192 597000 73388
rect 269864 73052 273196 73108
rect 273252 73052 273262 73108
rect 574952 72940 578620 72996
rect 578676 72940 578686 72996
rect 419944 72380 420140 72436
rect 420196 72380 423164 72436
rect 423220 72380 423230 72436
rect 457762 71596 457772 71652
rect 457828 71596 459396 71652
rect 459340 71540 460040 71596
rect 574952 70924 578284 70980
rect 578340 70924 578350 70980
rect 269864 70140 273308 70196
rect 273364 70140 273374 70196
rect 574952 68908 578060 68964
rect 578116 68908 578126 68964
rect 421810 68796 421820 68852
rect 421876 68796 422940 68852
rect 422996 68796 423006 68852
rect 458434 68236 458444 68292
rect 458500 68236 459396 68292
rect 459340 68180 460040 68236
rect 419944 67452 421820 67508
rect 421876 67452 421886 67508
rect 269864 67228 273084 67284
rect 273140 67228 273150 67284
rect 574952 66892 578172 66948
rect 578228 66892 578238 66948
rect -960 65044 480 65240
rect -960 65016 32732 65044
rect 392 64988 32732 65016
rect 32788 64988 32798 65044
rect 458210 64876 458220 64932
rect 458276 64876 459396 64932
rect 574578 64876 574588 64932
rect 574644 64876 574654 64932
rect 459340 64820 460040 64876
rect 269864 64316 273196 64372
rect 273252 64316 273262 64372
rect 574952 62860 578396 62916
rect 578452 62860 578462 62916
rect 419944 62524 420252 62580
rect 420308 62524 422716 62580
rect 422772 62524 422782 62580
rect 458098 61516 458108 61572
rect 458164 61516 459396 61572
rect 459340 61460 460040 61516
rect 269864 61404 276444 61460
rect 276500 61404 276510 61460
rect 574578 61068 574588 61124
rect 574644 61068 574654 61124
rect 574588 60872 574644 61068
rect 590482 60172 590492 60228
rect 590548 60200 595672 60228
rect 590548 60172 597000 60200
rect 595560 59976 597000 60172
rect 574952 58828 577948 58884
rect 578004 58828 578014 58884
rect 269864 58492 272860 58548
rect 272916 58492 272926 58548
rect 369404 58324 370104 58380
rect 367826 58268 367836 58324
rect 367892 58268 369460 58324
rect 457874 58156 457884 58212
rect 457940 58156 459396 58212
rect 459340 58100 460040 58156
rect 419944 57596 421708 57652
rect 421764 57596 421774 57652
rect 337586 57148 337596 57204
rect 337652 57148 367836 57204
rect 367892 57148 367902 57204
rect 574952 56812 576380 56868
rect 576436 56812 576446 56868
rect 269864 55580 288092 55636
rect 288148 55580 288158 55636
rect 457762 54796 457772 54852
rect 457828 54796 459396 54852
rect 574952 54796 576492 54852
rect 576548 54796 576558 54852
rect 459340 54740 460040 54796
rect 574466 52780 574476 52836
rect 574532 52780 574542 52836
rect 269864 52668 288988 52724
rect 289044 52668 289054 52724
rect 419272 52696 422492 52724
rect 419244 52668 422492 52696
rect 422548 52668 422558 52724
rect 419244 52164 419300 52668
rect 419234 52108 419244 52164
rect 419300 52108 419310 52164
rect 273074 51996 273084 52052
rect 273140 51996 420028 52052
rect 420084 51996 420094 52052
rect 272850 51884 272860 51940
rect 272916 51884 420252 51940
rect 420308 51884 420318 51940
rect 209346 51772 209356 51828
rect 209412 51772 275884 51828
rect 275940 51772 275950 51828
rect 288082 51772 288092 51828
rect 288148 51772 421708 51828
rect 421764 51772 421774 51828
rect 201730 51660 201740 51716
rect 201796 51660 272300 51716
rect 272356 51660 272366 51716
rect 288978 51660 288988 51716
rect 289044 51660 419244 51716
rect 419300 51660 419310 51716
rect 196018 51548 196028 51604
rect 196084 51548 270844 51604
rect 270900 51548 270910 51604
rect 190418 51436 190428 51492
rect 190484 51436 271068 51492
rect 271124 51436 271134 51492
rect 327394 51436 327404 51492
rect 327460 51436 459396 51492
rect 459340 51380 460040 51436
rect 173170 51324 173180 51380
rect 173236 51324 267484 51380
rect 267540 51324 267550 51380
rect 40002 51212 40012 51268
rect 40068 51212 87500 51268
rect 87556 51212 87566 51268
rect 89394 51212 89404 51268
rect 89460 51212 266924 51268
rect 266980 51212 266990 51268
rect -960 50932 480 51128
rect -960 50904 27692 50932
rect 392 50876 27692 50904
rect 27748 50876 27758 50932
rect 39666 50764 39676 50820
rect 39732 50764 45612 50820
rect 45668 50764 45678 50820
rect 574952 50764 577948 50820
rect 578004 50764 578014 50820
rect 41234 50652 41244 50708
rect 41300 50652 98924 50708
rect 98980 50652 98990 50708
rect 136994 50652 137004 50708
rect 137060 50652 325052 50708
rect 325108 50652 325118 50708
rect 41346 50540 41356 50596
rect 41412 50540 78988 50596
rect 87462 50540 87500 50596
rect 87556 50540 87566 50596
rect 89366 50540 89404 50596
rect 89460 50540 89470 50596
rect 173142 50540 173180 50596
rect 173236 50540 173246 50596
rect 178882 50540 178892 50596
rect 178948 50540 268828 50596
rect 268884 50540 268894 50596
rect 78932 50484 78988 50540
rect 40898 50428 40908 50484
rect 40964 50428 53228 50484
rect 53284 50428 53294 50484
rect 78932 50428 93212 50484
rect 93268 50428 93278 50484
rect 184594 50428 184604 50484
rect 184660 50428 268940 50484
rect 268996 50428 269006 50484
rect 45574 50316 45612 50372
rect 45668 50316 45678 50372
rect 190306 50316 190316 50372
rect 190372 50316 190428 50372
rect 190484 50316 190494 50372
rect 195990 50316 196028 50372
rect 196084 50316 196094 50372
rect 201702 50316 201740 50372
rect 201796 50316 201806 50372
rect 209318 50316 209356 50372
rect 209412 50316 209422 50372
rect 273186 50316 273196 50372
rect 273252 50316 420140 50372
rect 420196 50316 420206 50372
rect 276434 50204 276444 50260
rect 276500 50204 421820 50260
rect 421876 50204 421886 50260
rect 39778 50092 39788 50148
rect 39844 50092 76076 50148
rect 76132 50092 76142 50148
rect 39890 49980 39900 50036
rect 39956 49980 77980 50036
rect 78036 49980 78046 50036
rect 41010 49868 41020 49924
rect 41076 49868 81788 49924
rect 81844 49868 81854 49924
rect 167458 49868 167468 49924
rect 167524 49868 272972 49924
rect 273028 49868 273038 49924
rect 41122 49756 41132 49812
rect 41188 49756 83692 49812
rect 83748 49756 83758 49812
rect 152226 49756 152236 49812
rect 152292 49756 267372 49812
rect 267428 49756 267438 49812
rect 38210 49644 38220 49700
rect 38276 49644 104636 49700
rect 104692 49644 104702 49700
rect 156034 49644 156044 49700
rect 156100 49644 279132 49700
rect 279188 49644 279198 49700
rect 36866 49532 36876 49588
rect 36932 49532 110348 49588
rect 110404 49532 110414 49588
rect 114258 49532 114268 49588
rect 114324 49532 289996 49588
rect 290052 49532 290062 49588
rect 574952 48748 578620 48804
rect 578676 48748 578686 48804
rect 97346 48636 97356 48692
rect 97412 48636 277228 48692
rect 277284 48636 293580 48692
rect 293636 48636 337596 48692
rect 337652 48636 337662 48692
rect 207442 48524 207452 48580
rect 207508 48524 272412 48580
rect 272468 48524 272478 48580
rect 288642 48524 288652 48580
rect 288708 48524 322252 48580
rect 322308 48524 322318 48580
rect 280018 48412 280028 48468
rect 280084 48412 307916 48468
rect 307972 48412 307982 48468
rect 159842 48300 159852 48356
rect 159908 48300 275548 48356
rect 275604 48300 275614 48356
rect 285058 48300 285068 48356
rect 285124 48300 315084 48356
rect 315140 48300 315150 48356
rect 97010 48188 97020 48244
rect 97076 48188 288428 48244
rect 288484 48188 288494 48244
rect 74162 48076 74172 48132
rect 74228 48076 284844 48132
rect 284900 48076 284910 48132
rect 457986 48076 457996 48132
rect 458052 48076 459396 48132
rect 459340 48020 460040 48076
rect 91298 47964 91308 48020
rect 91364 47964 330092 48020
rect 330148 47964 330158 48020
rect 11330 47852 11340 47908
rect 11396 47852 97356 47908
rect 97412 47852 97422 47908
rect 102722 47852 102732 47908
rect 102788 47852 279804 47908
rect 279860 47852 279870 47908
rect 335570 47852 335580 47908
rect 335636 47852 457660 47908
rect 457716 47852 457726 47908
rect 212258 47740 212268 47796
rect 212324 47740 269052 47796
rect 269108 47740 269118 47796
rect 278338 47740 278348 47796
rect 278404 47740 300748 47796
rect 300804 47740 300814 47796
rect 188402 47628 188412 47684
rect 188468 47628 291564 47684
rect 291620 47628 291630 47684
rect 574952 46732 578508 46788
rect 578564 46732 578574 46788
rect 595560 46760 597000 46984
rect 161746 46396 161756 46452
rect 161812 46396 282268 46452
rect 282324 46396 282334 46452
rect 150322 46284 150332 46340
rect 150388 46284 274428 46340
rect 274484 46284 274494 46340
rect 100818 46172 100828 46228
rect 100884 46172 267596 46228
rect 267652 46172 267662 46228
rect 194114 45276 194124 45332
rect 194180 45276 281484 45332
rect 281540 45276 281550 45332
rect 171378 45164 171388 45220
rect 171444 45164 278124 45220
rect 278180 45164 278190 45220
rect 154130 45052 154140 45108
rect 154196 45052 284732 45108
rect 284788 45052 284798 45108
rect 148418 44940 148428 44996
rect 148484 44940 289884 44996
rect 289940 44940 289950 44996
rect 125570 44828 125580 44884
rect 125636 44828 279916 44884
rect 279972 44828 279982 44884
rect 131282 44716 131292 44772
rect 131348 44716 290108 44772
rect 290164 44716 290174 44772
rect 457650 44716 457660 44772
rect 457716 44716 459396 44772
rect 574952 44716 578172 44772
rect 578228 44716 578238 44772
rect 459340 44660 460040 44716
rect 119858 44604 119868 44660
rect 119924 44604 284956 44660
rect 285012 44604 285022 44660
rect 108434 44492 108444 44548
rect 108500 44492 291452 44548
rect 291508 44492 291518 44548
rect 335346 44492 335356 44548
rect 335412 44492 456988 44548
rect 457044 44492 457054 44548
rect 205538 44380 205548 44436
rect 205604 44380 282380 44436
rect 282436 44380 282446 44436
rect 203634 43372 203644 43428
rect 203700 43372 275660 43428
rect 275716 43372 275726 43428
rect 144610 43260 144620 43316
rect 144676 43260 277340 43316
rect 277396 43260 277406 43316
rect 112242 43148 112252 43204
rect 112308 43148 269052 43204
rect 269108 43148 269118 43204
rect 116050 43036 116060 43092
rect 116116 43036 275772 43092
rect 275828 43036 275838 43092
rect 106530 42924 106540 42980
rect 106596 42924 268940 42980
rect 268996 42924 269006 42980
rect 95106 42812 95116 42868
rect 95172 42812 267260 42868
rect 267316 42812 267326 42868
rect 335122 42812 335132 42868
rect 335188 42812 457100 42868
rect 457156 42812 457166 42868
rect 574952 42700 578172 42756
rect 578228 42700 578238 42756
rect 199938 41916 199948 41972
rect 200004 41916 276332 41972
rect 276388 41916 276398 41972
rect 175074 41804 175084 41860
rect 175140 41804 270620 41860
rect 270676 41804 270686 41860
rect 85698 41692 85708 41748
rect 85764 41692 286412 41748
rect 286468 41692 286478 41748
rect 79874 41580 79884 41636
rect 79940 41580 285964 41636
rect 286020 41580 286030 41636
rect 68450 41468 68460 41524
rect 68516 41468 284732 41524
rect 284788 41468 284798 41524
rect 62738 41356 62748 41412
rect 62804 41356 286636 41412
rect 286692 41356 286702 41412
rect 456978 41356 456988 41412
rect 457044 41356 459396 41412
rect 459340 41300 460040 41356
rect 57138 41244 57148 41300
rect 57204 41244 288316 41300
rect 288372 41244 288382 41300
rect 49410 41132 49420 41188
rect 49476 41132 289772 41188
rect 289828 41132 289838 41188
rect 574952 40684 576268 40740
rect 576324 40684 576334 40740
rect 135090 39676 135100 39732
rect 135156 39676 272860 39732
rect 272916 39676 272926 39732
rect 123666 39564 123676 39620
rect 123732 39564 270732 39620
rect 270788 39564 270798 39620
rect 117954 39452 117964 39508
rect 118020 39452 270508 39508
rect 270564 39452 270574 39508
rect 574952 38668 578284 38724
rect 578340 38668 578350 38724
rect 457090 37996 457100 38052
rect 457156 37996 459396 38052
rect 459340 37940 460040 37996
rect 211250 37884 211260 37940
rect 211316 37884 279692 37940
rect 279748 37884 279758 37940
rect 176978 37772 176988 37828
rect 177044 37772 288204 37828
rect 288260 37772 288270 37828
rect 424162 37772 424172 37828
rect 424228 37772 457660 37828
rect 457716 37772 457726 37828
rect -960 36820 480 37016
rect -960 36792 272636 36820
rect 392 36764 272636 36792
rect 272692 36764 272702 36820
rect 574952 36652 578060 36708
rect 578116 36652 578126 36708
rect 146514 36316 146524 36372
rect 146580 36316 273084 36372
rect 273140 36316 273150 36372
rect 140802 36204 140812 36260
rect 140868 36204 274316 36260
rect 274372 36204 274382 36260
rect 129378 36092 129388 36148
rect 129444 36092 272300 36148
rect 272356 36092 272366 36148
rect 457650 34636 457660 34692
rect 457716 34636 459396 34692
rect 574952 34636 578396 34692
rect 578452 34636 578462 34692
rect 459340 34580 460040 34636
rect 186498 34412 186508 34468
rect 186564 34412 272188 34468
rect 272244 34412 272254 34468
rect 589922 33740 589932 33796
rect 589988 33768 595672 33796
rect 589988 33740 597000 33768
rect 595560 33544 597000 33740
rect 138898 33068 138908 33124
rect 138964 33068 278908 33124
rect 278964 33068 278974 33124
rect 133186 32956 133196 33012
rect 133252 32956 274092 33012
rect 274148 32956 274158 33012
rect 127474 32844 127484 32900
rect 127540 32844 275548 32900
rect 275604 32844 275614 32900
rect 121762 32732 121772 32788
rect 121828 32732 274204 32788
rect 274260 32732 274270 32788
rect 574952 32620 578172 32676
rect 578228 32620 578238 32676
rect 427522 31276 427532 31332
rect 427588 31276 459396 31332
rect 459340 31220 460040 31276
rect 574952 30604 577948 30660
rect 578004 30604 578014 30660
rect 142818 29372 142828 29428
rect 142884 29372 288092 29428
rect 288148 29372 288158 29428
rect 574578 29260 574588 29316
rect 574644 29260 574654 29316
rect 574588 28616 574644 29260
rect 271506 27916 271516 27972
rect 271572 27916 459396 27972
rect 459340 27860 460040 27916
rect 182690 26124 182700 26180
rect 182756 26124 281372 26180
rect 281428 26124 281438 26180
rect 574588 26068 574644 26600
rect 165554 26012 165564 26068
rect 165620 26012 281596 26068
rect 281652 26012 281662 26068
rect 574578 26012 574588 26068
rect 574644 26012 574654 26068
rect 367826 24556 367836 24612
rect 367892 24556 459396 24612
rect 459340 24500 460040 24556
rect 574588 24052 574644 24584
rect 574578 23996 574588 24052
rect 574644 23996 574654 24052
rect 329186 22988 329196 23044
rect 329252 22988 578284 23044
rect 578340 22988 578350 23044
rect 392 22904 4172 22932
rect -960 22876 4172 22904
rect 4228 22876 4238 22932
rect 335906 22876 335916 22932
rect 335972 22876 574588 22932
rect 574644 22876 574654 22932
rect -960 22680 480 22876
rect 340274 22764 340284 22820
rect 340340 22764 578172 22820
rect 578228 22764 578238 22820
rect 328402 21756 328412 21812
rect 328468 21756 578508 21812
rect 578564 21756 578574 21812
rect 331874 21644 331884 21700
rect 331940 21644 578620 21700
rect 578676 21644 578686 21700
rect 340162 21532 340172 21588
rect 340228 21532 578060 21588
rect 578116 21532 578126 21588
rect 340386 21420 340396 21476
rect 340452 21420 578396 21476
rect 578452 21420 578462 21476
rect 340610 21308 340620 21364
rect 340676 21308 574588 21364
rect 574644 21308 574654 21364
rect 340946 21196 340956 21252
rect 341012 21196 577948 21252
rect 578004 21196 578014 21252
rect 595560 20356 597000 20552
rect 274754 20300 274764 20356
rect 274820 20328 597000 20356
rect 274820 20300 595672 20328
rect 327506 20076 327516 20132
rect 327572 20076 578172 20132
rect 578228 20076 578238 20132
rect 180786 19292 180796 19348
rect 180852 19292 272412 19348
rect 272468 19292 272478 19348
rect 192210 15932 192220 15988
rect 192276 15932 273868 15988
rect 273924 15932 273934 15988
rect 4162 12572 4172 12628
rect 4228 12572 26012 12628
rect 26068 12572 26078 12628
rect 163874 9212 163884 9268
rect 163940 9212 268828 9268
rect 268884 9212 268894 9268
rect 392 8792 4172 8820
rect -960 8764 4172 8792
rect 4228 8764 4238 8820
rect -960 8568 480 8764
rect 278002 7644 278012 7700
rect 278068 7644 582540 7700
rect 582596 7644 582606 7700
rect 158162 7532 158172 7588
rect 158228 7532 267148 7588
rect 267204 7532 267214 7588
rect 271394 7532 271404 7588
rect 271460 7532 580636 7588
rect 580692 7532 580702 7588
rect 595560 7140 597000 7336
rect 274642 7084 274652 7140
rect 274708 7112 597000 7140
rect 274708 7084 595672 7112
rect 271282 5852 271292 5908
rect 271348 5852 584444 5908
rect 584500 5852 584510 5908
rect 41580 5068 42084 5124
rect 41580 5012 41636 5068
rect 42028 5012 42084 5068
rect 38322 4956 38332 5012
rect 38388 4956 41636 5012
rect 41766 4956 41804 5012
rect 41860 4956 41870 5012
rect 42028 4956 47516 5012
rect 47572 4956 47582 5012
rect 33506 4844 33516 4900
rect 33572 4844 55132 4900
rect 55188 4844 55198 4900
rect 38434 4732 38444 4788
rect 38500 4732 60844 4788
rect 60900 4732 60910 4788
rect 35186 4620 35196 4676
rect 35252 4620 58940 4676
rect 58996 4620 59006 4676
rect 40114 4508 40124 4564
rect 40180 4508 64652 4564
rect 64708 4508 64718 4564
rect 41906 4396 41916 4452
rect 41972 4396 66556 4452
rect 66612 4396 66622 4452
rect 32498 4284 32508 4340
rect 32564 4284 34300 4340
rect 34356 4284 34366 4340
rect 40226 4284 40236 4340
rect 40292 4284 70364 4340
rect 70420 4284 70430 4340
rect 198146 4284 198156 4340
rect 198212 4284 273980 4340
rect 274036 4284 274046 4340
rect 15362 4172 15372 4228
rect 15428 4172 16716 4228
rect 16772 4172 16782 4228
rect 17266 4172 17276 4228
rect 17332 4172 18396 4228
rect 18452 4172 18462 4228
rect 19170 4172 19180 4228
rect 19236 4172 20076 4228
rect 20132 4172 20142 4228
rect 34402 4172 34412 4228
rect 34468 4172 35196 4228
rect 35252 4172 35262 4228
rect 38546 4172 38556 4228
rect 38612 4172 39900 4228
rect 39956 4172 39966 4228
rect 41458 4172 41468 4228
rect 41524 4172 72268 4228
rect 72324 4172 72334 4228
rect 169586 4172 169596 4228
rect 169652 4172 270508 4228
rect 270564 4172 270574 4228
<< via3 >>
rect 202972 591164 203028 591220
rect 203196 590828 203252 590884
rect 203084 590604 203140 590660
rect 188972 590156 189028 590212
rect 253708 590156 253764 590212
rect 341068 590156 341124 590212
rect 590492 588588 590548 588644
rect 202860 587244 202916 587300
rect 196476 587132 196532 587188
rect 529676 576492 529732 576548
rect 189420 576380 189476 576436
rect 532588 576380 532644 576436
rect 202748 576268 202804 576324
rect 189196 575372 189252 575428
rect 190428 575148 190484 575204
rect 478828 575148 478884 575204
rect 480620 575036 480676 575092
rect 189308 574812 189364 574868
rect 532812 574812 532868 574868
rect 201180 574700 201236 574756
rect 198044 574588 198100 574644
rect 478940 573804 478996 573860
rect 480508 573692 480564 573748
rect 199612 573580 199668 573636
rect 197820 573468 197876 573524
rect 197708 573356 197764 573412
rect 192892 573244 192948 573300
rect 529452 573244 529508 573300
rect 196252 573132 196308 573188
rect 193116 572124 193172 572180
rect 479052 572124 479108 572180
rect 200956 572012 201012 572068
rect 529564 572012 529620 572068
rect 201068 571900 201124 571956
rect 201292 571788 201348 571844
rect 533260 571788 533316 571844
rect 199388 571676 199444 571732
rect 197932 571564 197988 571620
rect 193004 571452 193060 571508
rect 199836 571340 199892 571396
rect 192668 571228 192724 571284
rect 479164 570332 479220 570388
rect 203532 570220 203588 570276
rect 533036 570220 533092 570276
rect 202524 570108 202580 570164
rect 532700 570108 532756 570164
rect 201516 569996 201572 570052
rect 192556 569884 192612 569940
rect 199500 569884 199556 569940
rect 196364 569772 196420 569828
rect 196028 568652 196084 568708
rect 202636 568540 202692 568596
rect 532924 568540 532980 568596
rect 195916 568428 195972 568484
rect 529340 568428 529396 568484
rect 196140 568316 196196 568372
rect 192780 568204 192836 568260
rect 200732 568092 200788 568148
rect 590716 568092 590772 568148
rect 198156 567980 198212 568036
rect 189532 567868 189588 567924
rect 199276 567308 199332 567364
rect 479276 567308 479332 567364
rect 191324 567196 191380 567252
rect 191436 567084 191492 567140
rect 190428 566972 190484 567028
rect 532812 565068 532868 565124
rect 532812 564844 532868 564900
rect 533260 564844 533316 564900
rect 532588 560364 532644 560420
rect 4396 558908 4452 558964
rect 533036 555660 533092 555716
rect 532924 550956 532980 551012
rect 184716 550732 184772 550788
rect 590828 549164 590884 549220
rect 532812 546252 532868 546308
rect 4172 544796 4228 544852
rect 184604 543564 184660 543620
rect 532700 541548 532756 541604
rect 529564 532140 529620 532196
rect 57932 530684 57988 530740
rect 186396 522060 186452 522116
rect 4508 516572 4564 516628
rect 590716 509516 590772 509572
rect 529452 508620 529508 508676
rect 180460 507724 180516 507780
rect 4284 502460 4340 502516
rect 180572 500556 180628 500612
rect 590604 496300 590660 496356
rect 529340 494508 529396 494564
rect 187292 493388 187348 493444
rect 529676 489804 529732 489860
rect 12572 488348 12628 488404
rect 188076 486220 188132 486276
rect 187180 479052 187236 479108
rect 4620 474236 4676 474292
rect 187964 471884 188020 471940
rect 590492 469868 590548 469924
rect 4396 469532 4452 469588
rect 167132 469532 167188 469588
rect 4508 467852 4564 467908
rect 168812 467852 168868 467908
rect 533148 466284 533204 466340
rect 4620 466172 4676 466228
rect 170492 466172 170548 466228
rect 187852 464716 187908 464772
rect 4508 460124 4564 460180
rect 187740 457548 187796 457604
rect 187404 450380 187460 450436
rect 187516 443212 187572 443268
rect 187628 436044 187684 436100
rect 162092 431900 162148 431956
rect 189084 428876 189140 428932
rect 532588 428652 532644 428708
rect 186284 421708 186340 421764
rect 4172 417788 4228 417844
rect 185612 414540 185668 414596
rect 62076 413420 62132 413476
rect 480508 410508 480564 410564
rect 359884 410396 359940 410452
rect 480620 410396 480676 410452
rect 479164 410172 479220 410228
rect 359548 410060 359604 410116
rect 478940 410060 478996 410116
rect 202300 409948 202356 410004
rect 83916 409836 83972 409892
rect 386204 409836 386260 409892
rect 404908 409836 404964 409892
rect 192668 409724 192724 409780
rect 202972 409724 203028 409780
rect 352828 409724 352884 409780
rect 359660 409724 359716 409780
rect 366268 409724 366324 409780
rect 188972 409612 189028 409668
rect 202860 409500 202916 409556
rect 203084 409388 203140 409444
rect 201180 409276 201236 409332
rect 240268 409276 240324 409332
rect 478828 409276 478884 409332
rect 496412 409276 496468 409332
rect 201068 409164 201124 409220
rect 479052 409164 479108 409220
rect 386092 409052 386148 409108
rect 199276 408940 199332 408996
rect 366044 408940 366100 408996
rect 369628 408940 369684 408996
rect 354508 408604 354564 408660
rect 374668 408604 374724 408660
rect 356188 408492 356244 408548
rect 384860 408492 384916 408548
rect 393484 408268 393540 408324
rect 366156 408156 366212 408212
rect 288092 408044 288148 408100
rect 479276 408044 479332 408100
rect 195916 407820 195972 407876
rect 278908 407820 278964 407876
rect 199388 407708 199444 407764
rect 342636 407708 342692 407764
rect 362796 407708 362852 407764
rect 328524 407596 328580 407652
rect 358540 407596 358596 407652
rect 197596 407484 197652 407540
rect 350476 407484 350532 407540
rect 362796 407484 362852 407540
rect 232316 407260 232372 407316
rect 192556 407148 192612 407204
rect 203196 407148 203252 407204
rect 196028 406700 196084 406756
rect 352156 406700 352212 406756
rect 383068 406700 383124 406756
rect 372764 406588 372820 406644
rect 434588 406588 434644 406644
rect 499324 406588 499380 406644
rect 501564 406588 501620 406644
rect 511868 406588 511924 406644
rect 514108 406588 514164 406644
rect 517020 406588 517076 406644
rect 522172 406588 522228 406644
rect 528892 406588 528948 406644
rect 543676 406588 543732 406644
rect 551068 406588 551124 406644
rect 558236 406588 558292 406644
rect 580636 406588 580692 406644
rect 196476 406476 196532 406532
rect 246876 406476 246932 406532
rect 362796 406476 362852 406532
rect 354620 406364 354676 406420
rect 340956 406140 341012 406196
rect 403228 406140 403284 406196
rect 338604 406028 338660 406084
rect 338828 405916 338884 405972
rect 202748 405804 202804 405860
rect 371308 405580 371364 405636
rect 347900 405356 347956 405412
rect 354732 405356 354788 405412
rect 357308 405356 357364 405412
rect 347788 405244 347844 405300
rect 393148 405244 393204 405300
rect 354508 405132 354564 405188
rect 367948 405132 368004 405188
rect 202748 405020 202804 405076
rect 356188 405020 356244 405076
rect 398188 405020 398244 405076
rect 202412 404908 202468 404964
rect 350588 404908 350644 404964
rect 350924 404908 350980 404964
rect 367612 404908 367668 404964
rect 367836 404908 367892 404964
rect 391468 404908 391524 404964
rect 199612 404796 199668 404852
rect 342524 404796 342580 404852
rect 342748 404796 342804 404852
rect 350700 404796 350756 404852
rect 362908 404796 362964 404852
rect 364812 404796 364868 404852
rect 527436 404796 527492 404852
rect 192780 404684 192836 404740
rect 439068 404684 439124 404740
rect 196140 404572 196196 404628
rect 383180 404460 383236 404516
rect 389676 404460 389732 404516
rect 389900 404460 389956 404516
rect 398300 404460 398356 404516
rect 197708 404348 197764 404404
rect 350812 404348 350868 404404
rect 363020 404348 363076 404404
rect 364700 404348 364756 404404
rect 366156 404348 366212 404404
rect 390572 404348 390628 404404
rect 395836 404348 395892 404404
rect 398412 404348 398468 404404
rect 398636 404348 398692 404404
rect 202524 404236 202580 404292
rect 351484 404236 351540 404292
rect 357868 404236 357924 404292
rect 367836 404236 367892 404292
rect 373660 404236 373716 404292
rect 447580 404236 447636 404292
rect 454972 404236 455028 404292
rect 565852 404236 565908 404292
rect 199500 404124 199556 404180
rect 389452 404124 389508 404180
rect 398412 404124 398468 404180
rect 196252 404012 196308 404068
rect 342524 404012 342580 404068
rect 374556 404012 374612 404068
rect 191324 403900 191380 403956
rect 346892 403900 346948 403956
rect 439068 403900 439124 403956
rect 367612 403788 367668 403844
rect 346892 403676 346948 403732
rect 364700 403676 364756 403732
rect 390572 403676 390628 403732
rect 398188 403676 398244 403732
rect 447580 403676 447636 403732
rect 356188 403564 356244 403620
rect 389788 403564 389844 403620
rect 352716 403452 352772 403508
rect 359772 403452 359828 403508
rect 374556 403452 374612 403508
rect 350476 403340 350532 403396
rect 359996 403340 360052 403396
rect 351036 403116 351092 403172
rect 357868 403116 357924 403172
rect 361228 403116 361284 403172
rect 384860 403116 384916 403172
rect 389900 403116 389956 403172
rect 393484 403116 393540 403172
rect 403228 403116 403284 403172
rect 347788 403004 347844 403060
rect 356636 403004 356692 403060
rect 363020 403004 363076 403060
rect 374668 403004 374724 403060
rect 383068 403004 383124 403060
rect 391468 403004 391524 403060
rect 393148 403004 393204 403060
rect 454972 403004 455028 403060
rect 342748 402892 342804 402948
rect 359884 402892 359940 402948
rect 373660 402892 373716 402948
rect 389676 402892 389732 402948
rect 434588 402892 434644 402948
rect 341180 402780 341236 402836
rect 395836 402780 395892 402836
rect 342636 402668 342692 402724
rect 367836 402668 367892 402724
rect 383180 402668 383236 402724
rect 389788 402668 389844 402724
rect 501564 402668 501620 402724
rect 189308 402556 189364 402612
rect 351484 402556 351540 402612
rect 366156 402556 366212 402612
rect 389452 402556 389508 402612
rect 350588 402444 350644 402500
rect 372764 402332 372820 402388
rect 527436 402332 527492 402388
rect 340172 402220 340228 402276
rect 336140 402108 336196 402164
rect 337596 402108 337652 402164
rect 197596 401548 197652 401604
rect 336140 401548 336196 401604
rect 196364 400988 196420 401044
rect 192892 400764 192948 400820
rect 201404 400652 201460 400708
rect 202636 400652 202692 400708
rect 201404 399868 201460 399924
rect 339612 399644 339668 399700
rect 197820 399308 197876 399364
rect 337596 399308 337652 399364
rect 189420 399196 189476 399252
rect 199276 399084 199332 399140
rect 184604 398972 184660 399028
rect 333564 398972 333620 399028
rect 199276 398188 199332 398244
rect 200956 398076 201012 398132
rect 202860 398076 202916 398132
rect 204764 398076 204820 398132
rect 193004 397852 193060 397908
rect 202860 397740 202916 397796
rect 201292 397628 201348 397684
rect 203532 397516 203588 397572
rect 339500 397516 339556 397572
rect 198044 396396 198100 396452
rect 337708 396284 337764 396340
rect 194908 395948 194964 396004
rect 197932 395948 197988 396004
rect 338828 395948 338884 396004
rect 198044 395836 198100 395892
rect 340620 395612 340676 395668
rect 194908 394828 194964 394884
rect 196252 394828 196308 394884
rect 333116 394828 333172 394884
rect 186284 394156 186340 394212
rect 333452 394156 333508 394212
rect 192444 393260 192500 393316
rect 334460 393260 334516 393316
rect 187180 393148 187236 393204
rect 334348 393148 334404 393204
rect 336924 392812 336980 392868
rect 337484 392812 337540 392868
rect 191548 392476 191604 392532
rect 193116 392476 193172 392532
rect 196476 391692 196532 391748
rect 186396 390908 186452 390964
rect 199612 390908 199668 390964
rect 201068 390796 201124 390852
rect 191436 390684 191492 390740
rect 201292 390460 201348 390516
rect 199500 390348 199556 390404
rect 590492 390348 590548 390404
rect 199388 390236 199444 390292
rect 330316 390236 330372 390292
rect 192556 389900 192612 389956
rect 330204 389900 330260 389956
rect 4284 389564 4340 389620
rect 201180 388780 201236 388836
rect 329756 388780 329812 388836
rect 196028 388332 196084 388388
rect 337820 388332 337876 388388
rect 317436 388220 317492 388276
rect 197484 387996 197540 388052
rect 331548 387996 331604 388052
rect 197484 386764 197540 386820
rect 197932 386764 197988 386820
rect 204540 386764 204596 386820
rect 339500 386764 339556 386820
rect 91532 386540 91588 386596
rect 204428 385196 204484 385252
rect 327404 385196 327460 385252
rect 91756 384972 91812 385028
rect 208348 384188 208404 384244
rect 199052 383740 199108 383796
rect 335916 383516 335972 383572
rect 197372 383180 197428 383236
rect 206668 382956 206724 383012
rect 237692 382956 237748 383012
rect 189532 382844 189588 382900
rect 202860 382620 202916 382676
rect 339052 382508 339108 382564
rect 201516 382396 201572 382452
rect 338604 382396 338660 382452
rect 199836 382284 199892 382340
rect 197708 382172 197764 382228
rect 198156 382172 198212 382228
rect 199724 382172 199780 382228
rect 199948 382172 200004 382228
rect 204092 382172 204148 382228
rect 237692 382060 237748 382116
rect 302316 382060 302372 382116
rect 303884 382060 303940 382116
rect 243516 381948 243572 382004
rect 263676 381948 263732 382004
rect 278796 381948 278852 382004
rect 297276 381948 297332 382004
rect 298956 381948 299012 382004
rect 300636 381948 300692 382004
rect 302204 381948 302260 382004
rect 303996 381948 304052 382004
rect 313404 381948 313460 382004
rect 261996 381612 262052 381668
rect 295596 381612 295652 381668
rect 305676 381612 305732 381668
rect 214508 381388 214564 381444
rect 216524 381388 216580 381444
rect 293916 381388 293972 381444
rect 197708 380604 197764 380660
rect 189532 380492 189588 380548
rect 209132 380492 209188 380548
rect 328636 380492 328692 380548
rect 209132 380044 209188 380100
rect 215852 379932 215908 379988
rect 218540 379596 218596 379652
rect 328636 379596 328692 379652
rect 329084 379596 329140 379652
rect 338492 379596 338548 379652
rect 190764 379484 190820 379540
rect 191324 379484 191380 379540
rect 192108 379484 192164 379540
rect 192668 379484 192724 379540
rect 193340 379484 193396 379540
rect 194684 379484 194740 379540
rect 195244 379484 195300 379540
rect 196364 379484 196420 379540
rect 193004 379260 193060 379316
rect 196140 379260 196196 379316
rect 213164 379260 213220 379316
rect 213836 379260 213892 379316
rect 215180 379260 215236 379316
rect 217196 379260 217252 379316
rect 204316 378700 204372 378756
rect 330092 378700 330148 378756
rect 587132 377356 587188 377412
rect 4284 377132 4340 377188
rect 165452 377132 165508 377188
rect 4172 375676 4228 375732
rect 330428 373100 330484 373156
rect 329420 372204 329476 372260
rect 340508 371308 340564 371364
rect 333340 370412 333396 370468
rect 340620 365932 340676 365988
rect 174748 363020 174804 363076
rect 338044 362348 338100 362404
rect 174860 361900 174916 361956
rect 176204 360780 176260 360836
rect 336364 360332 336420 360388
rect 174748 359772 174804 359828
rect 171388 359660 171444 359716
rect 177212 358540 177268 358596
rect 174860 356300 174916 356356
rect 330988 356076 331044 356132
rect 176204 353052 176260 353108
rect 590604 350700 590660 350756
rect 171388 349580 171444 349636
rect 4284 347228 4340 347284
rect 333452 344428 333508 344484
rect 332668 343532 332724 343588
rect 163772 338492 163828 338548
rect 177212 338492 177268 338548
rect 340620 335468 340676 335524
rect 332108 334572 332164 334628
rect 334572 334348 334628 334404
rect 329532 333676 329588 333732
rect 334572 332780 334628 332836
rect 329756 331884 329812 331940
rect 331100 330988 331156 331044
rect 337932 330092 337988 330148
rect 329756 329196 329812 329252
rect 334460 328300 334516 328356
rect 336812 327628 336868 327684
rect 338604 327404 338660 327460
rect 329308 326508 329364 326564
rect 163772 326060 163828 326116
rect 338492 325612 338548 325668
rect 338716 324716 338772 324772
rect 329308 323820 329364 323876
rect 335580 322924 335636 322980
rect 332332 322028 332388 322084
rect 329308 321132 329364 321188
rect 169596 320460 169652 320516
rect 331996 320236 332052 320292
rect 177100 319340 177156 319396
rect 334684 319340 334740 319396
rect 334460 318444 334516 318500
rect 336476 317548 336532 317604
rect 179564 317100 179620 317156
rect 333340 316988 333396 317044
rect 180124 315980 180180 316036
rect 332556 315980 332612 316036
rect 333788 315756 333844 315812
rect 336364 315756 336420 315812
rect 177548 314860 177604 314916
rect 334796 314860 334852 314916
rect 336364 314860 336420 314916
rect 329308 313964 329364 314020
rect 176204 313740 176260 313796
rect 4284 313292 4340 313348
rect 160412 313292 160468 313348
rect 329308 313068 329364 313124
rect 177884 312620 177940 312676
rect 340172 312172 340228 312228
rect 169484 311500 169540 311556
rect 338156 311276 338212 311332
rect 590716 311052 590772 311108
rect 174524 310380 174580 310436
rect 340284 310380 340340 310436
rect 339388 309484 339444 309540
rect 174300 309260 174356 309316
rect 330204 308812 330260 308868
rect 332220 308812 332276 308868
rect 333676 308588 333732 308644
rect 337596 308364 337652 308420
rect 333228 308252 333284 308308
rect 171276 308140 171332 308196
rect 333116 308028 333172 308084
rect 338044 307692 338100 307748
rect 180236 307020 180292 307076
rect 334012 306796 334068 306852
rect 179452 305900 179508 305956
rect 335020 305900 335076 305956
rect 332444 305676 332500 305732
rect 333788 305676 333844 305732
rect 333116 305004 333172 305060
rect 155372 304892 155428 304948
rect 167916 304780 167972 304836
rect 335468 304108 335524 304164
rect 334796 303996 334852 304052
rect 177772 303660 177828 303716
rect 334348 303212 334404 303268
rect 166236 302540 166292 302596
rect 333228 302316 333284 302372
rect 334012 302092 334068 302148
rect 336588 302092 336644 302148
rect 172956 301420 173012 301476
rect 331884 301420 331940 301476
rect 333676 300860 333732 300916
rect 337036 300748 337092 300804
rect 337820 300748 337876 300804
rect 331772 300524 331828 300580
rect 337820 300524 337876 300580
rect 174412 300300 174468 300356
rect 331324 299628 331380 299684
rect 330876 299292 330932 299348
rect 336476 299292 336532 299348
rect 177212 299180 177268 299236
rect 332556 299180 332612 299236
rect 332220 299068 332276 299124
rect 332668 299068 332724 299124
rect 331212 298732 331268 298788
rect 177324 298060 177380 298116
rect 329868 297836 329924 297892
rect 590828 297836 590884 297892
rect 332444 297388 332500 297444
rect 334684 297164 334740 297220
rect 177436 296940 177492 296996
rect 329644 296940 329700 296996
rect 335692 296492 335748 296548
rect 332780 296268 332836 296324
rect 333340 296268 333396 296324
rect 332780 296044 332836 296100
rect 177660 295820 177716 295876
rect 176092 294700 176148 294756
rect 335580 294700 335636 294756
rect 340396 294700 340452 294756
rect 72156 293916 72212 293972
rect 85596 293916 85652 293972
rect 334236 293916 334292 293972
rect 334460 293804 334516 293860
rect 333228 293692 333284 293748
rect 335244 293692 335300 293748
rect 108332 293132 108388 293188
rect 332780 293356 332836 293412
rect 334684 293356 334740 293412
rect 332780 293132 332836 293188
rect 333340 293132 333396 293188
rect 26012 292460 26068 292516
rect 333564 292460 333620 292516
rect 137788 292348 137844 292404
rect 333004 291564 333060 291620
rect 27692 291340 27748 291396
rect 335356 291004 335412 291060
rect 335020 290332 335076 290388
rect 338268 290332 338324 290388
rect 10892 290220 10948 290276
rect 332892 289772 332948 289828
rect 4284 289212 4340 289268
rect 96012 289212 96068 289268
rect 29372 289100 29428 289156
rect 336252 289100 336308 289156
rect 139244 288988 139300 289044
rect 162540 288876 162596 288932
rect 123452 287980 123508 288036
rect 337036 287980 337092 288036
rect 336700 287756 336756 287812
rect 332108 287420 332164 287476
rect 334796 287420 334852 287476
rect 332668 287084 332724 287140
rect 108332 286860 108388 286916
rect 335356 286748 335412 286804
rect 338156 286748 338212 286804
rect 336140 286188 336196 286244
rect 178892 285964 178948 286020
rect 180572 285964 180628 286020
rect 96012 285740 96068 285796
rect 330540 285740 330596 285796
rect 93660 285628 93716 285684
rect 163884 285628 163940 285684
rect 330876 285628 330932 285684
rect 335580 285516 335636 285572
rect 155372 285292 155428 285348
rect 330316 285292 330372 285348
rect 161868 284620 161924 284676
rect 333900 284396 333956 284452
rect 180460 283948 180516 284004
rect 336140 283836 336196 283892
rect 160412 283500 160468 283556
rect 334908 283500 334964 283556
rect 329308 282604 329364 282660
rect 165452 282380 165508 282436
rect 162540 282156 162596 282212
rect 163436 282156 163492 282212
rect 332108 282156 332164 282212
rect 333116 282156 333172 282212
rect 335356 282156 335412 282212
rect 178892 281932 178948 281988
rect 334460 281708 334516 281764
rect 332668 281372 332724 281428
rect 162092 281260 162148 281316
rect 334572 280812 334628 280868
rect 335020 280588 335076 280644
rect 161868 280476 161924 280532
rect 163996 280476 164052 280532
rect 93660 280364 93716 280420
rect 170492 280140 170548 280196
rect 179900 279916 179956 279972
rect 333116 279916 333172 279972
rect 330092 279580 330148 279636
rect 168812 279020 168868 279076
rect 339500 278124 339556 278180
rect 168924 278012 168980 278068
rect 167132 277900 167188 277956
rect 337708 277788 337764 277844
rect 335132 277340 335188 277396
rect 336700 277228 336756 277284
rect 332668 276332 332724 276388
rect 93996 276108 94052 276164
rect 164108 275884 164164 275940
rect 333116 275884 333172 275940
rect 334572 275884 334628 275940
rect 333452 275660 333508 275716
rect 163772 275548 163828 275604
rect 168476 275548 168532 275604
rect 330652 275548 330708 275604
rect 332108 275548 332164 275604
rect 334124 275548 334180 275604
rect 340396 275212 340452 275268
rect 169036 273868 169092 273924
rect 332556 273868 332612 273924
rect 334348 273868 334404 273924
rect 330764 272636 330820 272692
rect 332892 272636 332948 272692
rect 93436 271852 93492 271908
rect 165564 271852 165620 271908
rect 332892 271852 332948 271908
rect 590940 271404 590996 271460
rect 179676 271180 179732 271236
rect 167244 269836 167300 269892
rect 332108 268716 332164 268772
rect 332332 268044 332388 268100
rect 338156 268044 338212 268100
rect 163436 267820 163492 267876
rect 338940 267596 338996 267652
rect 174636 266700 174692 266756
rect 332668 266476 332724 266532
rect 334236 266252 334292 266308
rect 163996 265804 164052 265860
rect 176316 265580 176372 265636
rect 329308 265580 329364 265636
rect 330204 265468 330260 265524
rect 180572 265020 180628 265076
rect 340396 264684 340452 264740
rect 331660 264572 331716 264628
rect 337932 264572 337988 264628
rect 329868 264236 329924 264292
rect 333004 264236 333060 264292
rect 330540 264012 330596 264068
rect 331324 264012 331380 264068
rect 163884 263788 163940 263844
rect 336028 263900 336084 263956
rect 335132 263788 335188 263844
rect 334124 263676 334180 263732
rect 180012 263340 180068 263396
rect 333788 262892 333844 262948
rect 336924 262892 336980 262948
rect 337484 262892 337540 262948
rect 4284 262780 4340 262836
rect 180012 262220 180068 262276
rect 163772 261772 163828 261828
rect 138684 261660 138740 261716
rect 180684 261100 180740 261156
rect 333340 261100 333396 261156
rect 335916 260428 335972 260484
rect 330316 260316 330372 260372
rect 333228 260316 333284 260372
rect 334236 260316 334292 260372
rect 335468 260316 335524 260372
rect 180684 259980 180740 260036
rect 330092 259868 330148 259924
rect 334684 259868 334740 259924
rect 338380 259644 338436 259700
rect 336476 259308 336532 259364
rect 180684 258860 180740 258916
rect 329980 258636 330036 258692
rect 330876 258524 330932 258580
rect 331660 258524 331716 258580
rect 591052 258188 591108 258244
rect 336252 257516 336308 257572
rect 180572 257180 180628 257236
rect 336028 257180 336084 257236
rect 333676 257068 333732 257124
rect 334796 257068 334852 257124
rect 336140 257068 336196 257124
rect 339500 257068 339556 257124
rect 179676 256620 179732 256676
rect 333004 256172 333060 256228
rect 334348 256172 334404 256228
rect 333116 255724 333172 255780
rect 180348 255500 180404 255556
rect 334236 255276 334292 255332
rect 335692 255276 335748 255332
rect 338044 254940 338100 254996
rect 333228 254828 333284 254884
rect 337708 254604 337764 254660
rect 176988 254380 177044 254436
rect 336252 253932 336308 253988
rect 332220 253708 332276 253764
rect 334908 253708 334964 253764
rect 333788 253596 333844 253652
rect 334684 253596 334740 253652
rect 337820 253596 337876 253652
rect 336476 253484 336532 253540
rect 332668 253148 332724 253204
rect 180572 252700 180628 252756
rect 330092 252476 330148 252532
rect 329980 252364 330036 252420
rect 331212 252364 331268 252420
rect 180684 252140 180740 252196
rect 336028 252140 336084 252196
rect 333452 252028 333508 252084
rect 333788 251244 333844 251300
rect 333452 250572 333508 250628
rect 330764 250348 330820 250404
rect 332444 250348 332500 250404
rect 332780 250348 332836 250404
rect 336476 250236 336532 250292
rect 332332 249452 332388 249508
rect 333004 248892 333060 248948
rect 335916 248780 335972 248836
rect 331212 248668 331268 248724
rect 337932 248668 337988 248724
rect 338268 248668 338324 248724
rect 339948 248556 340004 248612
rect 4620 248444 4676 248500
rect 330988 246988 331044 247044
rect 336588 246988 336644 247044
rect 337372 246988 337428 247044
rect 339276 246988 339332 247044
rect 332444 246876 332500 246932
rect 334124 246876 334180 246932
rect 337260 246876 337316 246932
rect 339500 246876 339556 246932
rect 333228 245420 333284 245476
rect 329756 245308 329812 245364
rect 333676 245308 333732 245364
rect 334796 245308 334852 245364
rect 332108 245196 332164 245252
rect 336028 245196 336084 245252
rect 330540 244972 330596 245028
rect 332108 244972 332164 245028
rect 330876 244860 330932 244916
rect 334236 244860 334292 244916
rect 336476 244076 336532 244132
rect 334236 243740 334292 243796
rect 337708 243740 337764 243796
rect 333900 243516 333956 243572
rect 336028 243516 336084 243572
rect 337820 243516 337876 243572
rect 332668 243404 332724 243460
rect 333676 243404 333732 243460
rect 334124 243180 334180 243236
rect 336924 243180 336980 243236
rect 330988 242060 331044 242116
rect 332892 241948 332948 242004
rect 338940 241948 338996 242004
rect 332444 240716 332500 240772
rect 338156 240716 338212 240772
rect 326508 240604 326564 240660
rect 332220 240604 332276 240660
rect 197372 240492 197428 240548
rect 202524 240492 202580 240548
rect 199164 240380 199220 240436
rect 294812 240380 294868 240436
rect 327516 240380 327572 240436
rect 329980 240380 330036 240436
rect 328524 240268 328580 240324
rect 330204 240268 330260 240324
rect 336364 240268 336420 240324
rect 334572 240156 334628 240212
rect 335132 240156 335188 240212
rect 184828 240044 184884 240100
rect 202412 240044 202468 240100
rect 334460 240044 334516 240100
rect 335020 240044 335076 240100
rect 335356 240044 335412 240100
rect 204428 239932 204484 239988
rect 335580 239932 335636 239988
rect 321804 239820 321860 239876
rect 177548 239708 177604 239764
rect 268044 239708 268100 239764
rect 177212 239596 177268 239652
rect 275660 239596 275716 239652
rect 278124 239596 278180 239652
rect 278348 239484 278404 239540
rect 186284 239372 186340 239428
rect 204316 239372 204372 239428
rect 334460 239372 334516 239428
rect 186396 239260 186452 239316
rect 335356 239260 335412 239316
rect 335132 238812 335188 238868
rect 331548 238588 331604 238644
rect 332332 238588 332388 238644
rect 138572 238364 138628 238420
rect 204764 238364 204820 238420
rect 334684 238476 334740 238532
rect 187516 238252 187572 238308
rect 295260 238252 295316 238308
rect 324268 238252 324324 238308
rect 325836 238252 325892 238308
rect 330316 238252 330372 238308
rect 325724 238140 325780 238196
rect 330876 238140 330932 238196
rect 268828 238028 268884 238084
rect 298284 238028 298340 238084
rect 298284 237804 298340 237860
rect 68012 237692 68068 237748
rect 288876 237692 288932 237748
rect 71596 237580 71652 237636
rect 235116 237132 235172 237188
rect 234220 237020 234276 237076
rect 265244 237020 265300 237076
rect 268716 237020 268772 237076
rect 270396 237020 270452 237076
rect 275324 237020 275380 237076
rect 278796 237020 278852 237076
rect 293916 237020 293972 237076
rect 226716 236908 226772 236964
rect 231756 236908 231812 236964
rect 233436 236908 233492 236964
rect 265356 236908 265412 236964
rect 266812 236908 266868 236964
rect 267036 236908 267092 236964
rect 268604 236908 268660 236964
rect 270284 236908 270340 236964
rect 272076 236908 272132 236964
rect 275436 236908 275492 236964
rect 277116 236908 277172 236964
rect 278684 236908 278740 236964
rect 290556 236908 290612 236964
rect 293804 236908 293860 236964
rect 295372 236908 295428 236964
rect 298956 236908 299012 236964
rect 305676 236908 305732 236964
rect 178892 236796 178948 236852
rect 191548 236796 191604 236852
rect 325052 236796 325108 236852
rect 328636 236796 328692 236852
rect 197708 236684 197764 236740
rect 282604 236684 282660 236740
rect 289772 236684 289828 236740
rect 332668 236684 332724 236740
rect 187404 236572 187460 236628
rect 276556 236572 276612 236628
rect 288092 236572 288148 236628
rect 199388 236460 199444 236516
rect 308252 236460 308308 236516
rect 202972 236348 203028 236404
rect 191548 236236 191604 236292
rect 192556 236236 192612 236292
rect 330540 236236 330596 236292
rect 198940 236124 198996 236180
rect 330316 236124 330372 236180
rect 203308 236012 203364 236068
rect 204540 236012 204596 236068
rect 332668 236012 332724 236068
rect 204092 235900 204148 235956
rect 326508 235900 326564 235956
rect 327404 235900 327460 235956
rect 189420 235788 189476 235844
rect 333676 235788 333732 235844
rect 188076 235676 188132 235732
rect 203308 235676 203364 235732
rect 183932 235116 183988 235172
rect 202524 235116 202580 235172
rect 202748 235116 202804 235172
rect 267260 235116 267316 235172
rect 290108 235116 290164 235172
rect 326844 235116 326900 235172
rect 266924 235004 266980 235060
rect 280140 235004 280196 235060
rect 330092 235004 330148 235060
rect 189308 234892 189364 234948
rect 289660 234892 289716 234948
rect 289884 234892 289940 234948
rect 291452 234556 291508 234612
rect 336140 234556 336196 234612
rect 284732 234444 284788 234500
rect 333788 234444 333844 234500
rect 202524 234332 202580 234388
rect 308476 234332 308532 234388
rect 254492 234220 254548 234276
rect 42812 233436 42868 233492
rect 197820 233436 197876 233492
rect 198044 233436 198100 233492
rect 291564 233436 291620 233492
rect 199052 233324 199108 233380
rect 288428 233324 288484 233380
rect 328748 233324 328804 233380
rect 177884 233212 177940 233268
rect 269500 233212 269556 233268
rect 328412 233212 328468 233268
rect 325276 232876 325332 232932
rect 198044 232764 198100 232820
rect 279804 232764 279860 232820
rect 195692 232652 195748 232708
rect 335468 232652 335524 232708
rect 591164 231868 591220 231924
rect 267484 231756 267540 231812
rect 288204 231756 288260 231812
rect 328300 231756 328356 231812
rect 197596 231644 197652 231700
rect 286636 231644 286692 231700
rect 333228 231644 333284 231700
rect 167916 231532 167972 231588
rect 272300 231532 272356 231588
rect 201068 231084 201124 231140
rect 268940 230972 268996 231028
rect 284844 230972 284900 231028
rect 335804 230972 335860 231028
rect 289996 230860 290052 230916
rect 326620 230860 326676 230916
rect 166236 229852 166292 229908
rect 273308 229852 273364 229908
rect 196140 229404 196196 229460
rect 325164 229404 325220 229460
rect 284956 229292 285012 229348
rect 270508 227612 270564 227668
rect 279916 227612 279972 227668
rect 326732 227612 326788 227668
rect 269052 227500 269108 227556
rect 202860 226492 202916 226548
rect 271292 226492 271348 226548
rect 204652 226380 204708 226436
rect 278012 226380 278068 226436
rect 177772 226268 177828 226324
rect 273980 226268 274036 226324
rect 201180 226044 201236 226100
rect 333788 226044 333844 226100
rect 192892 225932 192948 225988
rect 330092 225932 330148 225988
rect 177324 224924 177380 224980
rect 270620 224924 270676 224980
rect 197932 224700 197988 224756
rect 41916 224364 41972 224420
rect 177436 223356 177492 223412
rect 275772 223356 275828 223412
rect 194684 222908 194740 222964
rect 274988 222908 275044 222964
rect 202300 222796 202356 222852
rect 293356 222796 293412 222852
rect 198156 221452 198212 221508
rect 199500 221340 199556 221396
rect 290668 221340 290724 221396
rect 177660 221228 177716 221284
rect 273868 221228 273924 221284
rect 200732 221004 200788 221060
rect 326732 221004 326788 221060
rect 108332 220220 108388 220276
rect 204876 219996 204932 220052
rect 276444 219996 276500 220052
rect 174300 219884 174356 219940
rect 272524 219884 272580 219940
rect 192444 219548 192500 219604
rect 323932 219548 323988 219604
rect 323372 219212 323428 219268
rect 591276 218540 591332 218596
rect 195804 218316 195860 218372
rect 293244 218316 293300 218372
rect 171276 218204 171332 218260
rect 273196 218204 273252 218260
rect 179676 218092 179732 218148
rect 283276 218092 283332 218148
rect 323148 217532 323204 217588
rect 193340 216524 193396 216580
rect 281708 216524 281764 216580
rect 179452 216412 179508 216468
rect 272636 216412 272692 216468
rect 177100 216300 177156 216356
rect 271516 216300 271572 216356
rect 169484 216188 169540 216244
rect 272860 216188 272916 216244
rect 288652 216076 288708 216132
rect 202636 214956 202692 215012
rect 285292 214956 285348 215012
rect 193004 214844 193060 214900
rect 278236 214844 278292 214900
rect 180348 214732 180404 214788
rect 271740 214732 271796 214788
rect 187292 214620 187348 214676
rect 280252 214620 280308 214676
rect 285068 214508 285124 214564
rect 196364 214396 196420 214452
rect 323372 214396 323428 214452
rect 337148 213948 337204 214004
rect 337148 213388 337204 213444
rect 177548 213276 177604 213332
rect 280028 212828 280084 212884
rect 180012 212716 180068 212772
rect 293132 212716 293188 212772
rect 199276 212604 199332 212660
rect 281596 212604 281652 212660
rect 283052 212380 283108 212436
rect 281372 211484 281428 211540
rect 267708 211372 267764 211428
rect 267932 211260 267988 211316
rect 180236 211036 180292 211092
rect 273420 211036 273476 211092
rect 267708 210924 267764 210980
rect 4284 210812 4340 210868
rect 123452 210812 123508 210868
rect 169596 210812 169652 210868
rect 327628 210812 327684 210868
rect 267932 210700 267988 210756
rect 176092 210588 176148 210644
rect 241388 210028 241444 210084
rect 189532 209916 189588 209972
rect 179564 209804 179620 209860
rect 272300 209804 272356 209860
rect 176204 209692 176260 209748
rect 272412 209692 272468 209748
rect 275548 209692 275604 209748
rect 174524 209580 174580 209636
rect 272748 209580 272804 209636
rect 174412 209468 174468 209524
rect 172956 209356 173012 209412
rect 273308 209132 273364 209188
rect 180124 209020 180180 209076
rect 269612 209020 269668 209076
rect 241388 208908 241444 208964
rect 4060 206332 4116 206388
rect 272972 206332 273028 206388
rect 269612 204764 269668 204820
rect 328636 204428 328692 204484
rect 270508 203308 270564 203364
rect 272188 203196 272244 203252
rect 272860 203196 272916 203252
rect 270732 203084 270788 203140
rect 295148 202748 295204 202804
rect 325388 202636 325444 202692
rect 308252 202524 308308 202580
rect 328412 202524 328468 202580
rect 308476 202412 308532 202468
rect 335804 202412 335860 202468
rect 269612 201404 269668 201460
rect 301196 199948 301252 200004
rect 301420 199948 301476 200004
rect 326956 199948 327012 200004
rect 328524 199948 328580 200004
rect 293692 199836 293748 199892
rect 308588 199388 308644 199444
rect 310828 199388 310884 199444
rect 311836 199388 311892 199444
rect 325276 199388 325332 199444
rect 273756 199164 273812 199220
rect 310268 199276 310324 199332
rect 290444 199052 290500 199108
rect 301420 199052 301476 199108
rect 310604 199052 310660 199108
rect 324044 199052 324100 199108
rect 310828 198940 310884 198996
rect 323260 198940 323316 198996
rect 292236 198828 292292 198884
rect 308588 198828 308644 198884
rect 311836 198828 311892 198884
rect 301196 198604 301252 198660
rect 326620 198604 326676 198660
rect 272412 198268 272468 198324
rect 337260 198268 337316 198324
rect 337708 198268 337764 198324
rect 332668 198156 332724 198212
rect 333900 198156 333956 198212
rect 336140 198044 336196 198100
rect 305676 197820 305732 197876
rect 321804 197708 321860 197764
rect 323372 197708 323428 197764
rect 289660 197596 289716 197652
rect 339388 197596 339444 197652
rect 332668 197484 332724 197540
rect 272748 197372 272804 197428
rect 273420 197372 273476 197428
rect 336140 197372 336196 197428
rect 339388 197260 339444 197316
rect 340060 197260 340116 197316
rect 339500 197148 339556 197204
rect 269500 195356 269556 195412
rect 272188 192444 272244 192500
rect 31052 191996 31108 192052
rect 590380 192108 590436 192164
rect 336028 191436 336084 191492
rect 272860 190652 272916 190708
rect 330764 189756 330820 189812
rect 334796 189756 334852 189812
rect 337932 189756 337988 189812
rect 272972 189532 273028 189588
rect 329084 188972 329140 189028
rect 338940 188972 338996 189028
rect 327068 188076 327124 188132
rect 334124 188076 334180 188132
rect 334460 188076 334516 188132
rect 272524 186620 272580 186676
rect 272412 186396 272468 186452
rect 334124 184940 334180 184996
rect 273196 183708 273252 183764
rect 337372 183708 337428 183764
rect 337372 182252 337428 182308
rect 272748 180796 272804 180852
rect 337260 179676 337316 179732
rect 337820 179676 337876 179732
rect 273644 178444 273700 178500
rect 333900 178444 333956 178500
rect 4284 177996 4340 178052
rect 272636 177884 272692 177940
rect 271852 176316 271908 176372
rect 328636 174636 328692 174692
rect 336028 174636 336084 174692
rect 273980 172060 274036 172116
rect 336140 171164 336196 171220
rect 336028 168252 336084 168308
rect 327628 166012 327684 166068
rect 39452 163772 39508 163828
rect 327628 161868 327684 161924
rect 422604 161084 422660 161140
rect 422828 160972 422884 161028
rect 467852 160860 467908 160916
rect 271740 160636 271796 160692
rect 590380 160636 590436 160692
rect 590716 160524 590772 160580
rect 275660 160412 275716 160468
rect 280252 160412 280308 160468
rect 297500 160300 297556 160356
rect 422604 159964 422660 160020
rect 422828 159964 422884 160020
rect 467852 159964 467908 160020
rect 591276 159628 591332 159684
rect 283276 159404 283332 159460
rect 591164 159404 591220 159460
rect 293244 159292 293300 159348
rect 590940 159292 590996 159348
rect 357868 159180 357924 159236
rect 341516 158844 341572 158900
rect 324268 158732 324324 158788
rect 281484 158620 281540 158676
rect 590604 158620 590660 158676
rect 558460 157612 558516 157668
rect 270620 157500 270676 157556
rect 514108 157500 514164 157556
rect 328860 156156 328916 156212
rect 337372 156044 337428 156100
rect 328076 155820 328132 155876
rect 278684 155708 278740 155764
rect 337260 155596 337316 155652
rect 578508 155596 578564 155652
rect 295148 155372 295204 155428
rect 574028 155372 574084 155428
rect 341180 155260 341236 155316
rect 341516 155260 341572 155316
rect 275772 154588 275828 154644
rect 293132 154476 293188 154532
rect 591276 154476 591332 154532
rect 293804 153916 293860 153972
rect 325388 153804 325444 153860
rect 281596 153692 281652 153748
rect 590828 153692 590884 153748
rect 574476 153020 574532 153076
rect 333676 152908 333732 152964
rect 338828 152796 338884 152852
rect 590044 152684 590100 152740
rect 333564 152124 333620 152180
rect 574700 152124 574756 152180
rect 292236 152012 292292 152068
rect 273868 151676 273924 151732
rect 331660 151116 331716 151172
rect 328524 150780 328580 150836
rect 578396 150780 578452 150836
rect 275324 150668 275380 150724
rect 278796 150556 278852 150612
rect 277116 150444 277172 150500
rect 275436 150332 275492 150388
rect 7532 149884 7588 149940
rect 462924 149660 462980 149716
rect 337484 149548 337540 149604
rect 272076 148988 272132 149044
rect 463708 148092 463764 148148
rect 575036 148092 575092 148148
rect 336028 147868 336084 147924
rect 337596 147868 337652 147924
rect 341404 147756 341460 147812
rect 288876 147308 288932 147364
rect 466396 146300 466452 146356
rect 462812 146188 462868 146244
rect 273644 146076 273700 146132
rect 327628 146076 327684 146132
rect 272636 145852 272692 145908
rect 273644 145852 273700 145908
rect 293916 145292 293972 145348
rect 341292 145180 341348 145236
rect 270284 145068 270340 145124
rect 520156 143948 520212 144004
rect 270620 143612 270676 143668
rect 520156 143612 520212 143668
rect 472892 143164 472948 143220
rect 576492 143164 576548 143220
rect 468636 143052 468692 143108
rect 578284 143052 578340 143108
rect 490028 142828 490084 142884
rect 497868 142828 497924 142884
rect 505708 142828 505764 142884
rect 507276 142828 507332 142884
rect 508844 142828 508900 142884
rect 511980 142828 512036 142884
rect 513548 142828 513604 142884
rect 335020 142604 335076 142660
rect 340620 142604 340676 142660
rect 463708 142604 463764 142660
rect 336028 142492 336084 142548
rect 335916 142268 335972 142324
rect 338940 142268 338996 142324
rect 578732 142268 578788 142324
rect 270396 142156 270452 142212
rect 479612 141708 479668 141764
rect 463036 141372 463092 141428
rect 466284 141260 466340 141316
rect 479612 141260 479668 141316
rect 466620 141148 466676 141204
rect 295372 141036 295428 141092
rect 330204 140924 330260 140980
rect 324044 140700 324100 140756
rect 323260 140476 323316 140532
rect 293692 140364 293748 140420
rect 290444 140252 290500 140308
rect 336140 140028 336196 140084
rect 480620 139692 480676 139748
rect 466172 139580 466228 139636
rect 482188 139580 482244 139636
rect 467068 139468 467124 139524
rect 501676 139468 501732 139524
rect 590156 139356 590212 139412
rect 337260 139132 337316 139188
rect 338492 139020 338548 139076
rect 578172 139020 578228 139076
rect 325276 138684 325332 138740
rect 323932 138572 323988 138628
rect 578620 138572 578676 138628
rect 290556 138460 290612 138516
rect 501676 138460 501732 138516
rect 272188 137116 272244 137172
rect 330428 135996 330484 136052
rect 457996 135996 458052 136052
rect 29372 135548 29428 135604
rect 339948 135436 340004 135492
rect 332668 134316 332724 134372
rect 333340 134316 333396 134372
rect 336812 134316 336868 134372
rect 327964 134092 328020 134148
rect 330652 132076 330708 132132
rect 273196 131292 273252 131348
rect 341516 130956 341572 131012
rect 335692 128716 335748 128772
rect 280140 128380 280196 128436
rect 337148 127596 337204 127652
rect 272972 125468 273028 125524
rect 332556 125356 332612 125412
rect 423276 122668 423332 122724
rect 335244 121996 335300 122052
rect 333900 121772 333956 121828
rect 331884 118636 331940 118692
rect 304892 116732 304948 116788
rect 331772 115276 331828 115332
rect 306572 113820 306628 113876
rect 575148 113820 575204 113876
rect 271628 113372 271684 113428
rect 590828 113036 590884 113092
rect 332108 111916 332164 111972
rect 293132 110908 293188 110964
rect 335804 110348 335860 110404
rect 458108 110348 458164 110404
rect 328412 110124 328468 110180
rect 457884 110124 457940 110180
rect 274876 110012 274932 110068
rect 327292 108556 327348 108612
rect 14252 107324 14308 107380
rect 334124 106988 334180 107044
rect 421820 106988 421876 107044
rect 335468 106652 335524 106708
rect 457772 106652 457828 106708
rect 269948 105308 270004 105364
rect 325724 105196 325780 105252
rect 270060 104972 270116 105028
rect 413308 104076 413364 104132
rect 414988 104076 415044 104132
rect 406700 103964 406756 104020
rect 403228 103852 403284 103908
rect 280252 102172 280308 102228
rect 329644 101836 329700 101892
rect 336924 101724 336980 101780
rect 458556 101724 458612 101780
rect 332220 101612 332276 101668
rect 456988 101612 457044 101668
rect 334012 100156 334068 100212
rect 421708 100156 421764 100212
rect 330540 100044 330596 100100
rect 458220 100044 458276 100100
rect 330316 99932 330372 99988
rect 458444 99932 458500 99988
rect 590716 99820 590772 99876
rect 274988 99260 275044 99316
rect 336812 99036 336868 99092
rect 337036 99036 337092 99092
rect 333452 98924 333508 98980
rect 458332 98924 458388 98980
rect 330092 98812 330148 98868
rect 326732 98700 326788 98756
rect 325836 98588 325892 98644
rect 457548 98588 457604 98644
rect 329868 98476 329924 98532
rect 295036 98364 295092 98420
rect 294812 98252 294868 98308
rect 457996 98252 458052 98308
rect 456988 97580 457044 97636
rect 421820 97020 421876 97076
rect 424172 97020 424228 97076
rect 366268 93996 366324 94052
rect 367052 93996 367108 94052
rect 10892 93436 10948 93492
rect 366268 91532 366324 91588
rect 421708 91532 421764 91588
rect 427532 91532 427588 91588
rect 578844 91084 578900 91140
rect 575036 89628 575092 89684
rect 458556 88396 458612 88452
rect 578508 87052 578564 87108
rect 457548 85036 457604 85092
rect 578732 85036 578788 85092
rect 276444 84812 276500 84868
rect 332668 83132 332724 83188
rect 574924 83020 574980 83076
rect 574812 81004 574868 81060
rect 4284 79100 4340 79156
rect 578396 78988 578452 79044
rect 578060 76972 578116 77028
rect 458332 74956 458388 75012
rect 574700 74956 574756 75012
rect 590604 73388 590660 73444
rect 578620 72940 578676 72996
rect 578284 70924 578340 70980
rect 458444 68236 458500 68292
rect 578172 66892 578228 66948
rect 32732 64988 32788 65044
rect 458220 64876 458276 64932
rect 574588 64876 574644 64932
rect 458108 61516 458164 61572
rect 574588 61068 574644 61124
rect 590492 60172 590548 60228
rect 577948 58828 578004 58884
rect 457884 58156 457940 58212
rect 576380 56812 576436 56868
rect 457772 54796 457828 54852
rect 576492 54796 576548 54852
rect 574476 52780 574532 52836
rect 209356 51772 209412 51828
rect 201740 51660 201796 51716
rect 196028 51548 196084 51604
rect 190428 51436 190484 51492
rect 327404 51436 327460 51492
rect 173180 51324 173236 51380
rect 267484 51324 267540 51380
rect 87500 51212 87556 51268
rect 89404 51212 89460 51268
rect 266924 51212 266980 51268
rect 27692 50876 27748 50932
rect 45612 50764 45668 50820
rect 577948 50764 578004 50820
rect 325052 50652 325108 50708
rect 87500 50540 87556 50596
rect 89404 50540 89460 50596
rect 173180 50540 173236 50596
rect 45612 50316 45668 50372
rect 190428 50316 190484 50372
rect 196028 50316 196084 50372
rect 201740 50316 201796 50372
rect 209356 50316 209412 50372
rect 267372 49756 267428 49812
rect 289996 49532 290052 49588
rect 288652 48524 288708 48580
rect 280028 48412 280084 48468
rect 275548 48300 275604 48356
rect 285068 48300 285124 48356
rect 288428 48188 288484 48244
rect 284844 48076 284900 48132
rect 457996 48076 458052 48132
rect 279804 47852 279860 47908
rect 335580 47852 335636 47908
rect 457660 47852 457716 47908
rect 278348 47740 278404 47796
rect 291564 47628 291620 47684
rect 267596 46172 267652 46228
rect 278124 45164 278180 45220
rect 289884 44940 289940 44996
rect 279916 44828 279972 44884
rect 290108 44716 290164 44772
rect 457660 44716 457716 44772
rect 578172 44716 578228 44772
rect 284956 44604 285012 44660
rect 291452 44492 291508 44548
rect 335356 44492 335412 44548
rect 456988 44492 457044 44548
rect 269052 43148 269108 43204
rect 268940 42924 268996 42980
rect 267260 42812 267316 42868
rect 335132 42812 335188 42868
rect 457100 42812 457156 42868
rect 286412 41692 286468 41748
rect 284732 41468 284788 41524
rect 286636 41356 286692 41412
rect 456988 41356 457044 41412
rect 288316 41244 288372 41300
rect 289772 41132 289828 41188
rect 576268 40684 576324 40740
rect 272860 39676 272916 39732
rect 270508 39452 270564 39508
rect 457100 37996 457156 38052
rect 279692 37884 279748 37940
rect 288204 37772 288260 37828
rect 424172 37772 424228 37828
rect 457660 37772 457716 37828
rect 272636 36764 272692 36820
rect 578060 36652 578116 36708
rect 273084 36316 273140 36372
rect 272300 36092 272356 36148
rect 457660 34636 457716 34692
rect 589932 33740 589988 33796
rect 578172 32620 578228 32676
rect 427532 31276 427588 31332
rect 288092 29372 288148 29428
rect 574588 29260 574644 29316
rect 271516 27916 271572 27972
rect 574588 26012 574644 26068
rect 4172 22876 4228 22932
rect 574588 22876 574644 22932
rect 340284 22764 340340 22820
rect 578172 22764 578228 22820
rect 340172 21532 340228 21588
rect 578060 21532 578116 21588
rect 340396 21420 340452 21476
rect 274764 20300 274820 20356
rect 327516 20076 327572 20132
rect 272412 19292 272468 19348
rect 4172 12572 4228 12628
rect 26012 12572 26068 12628
rect 268828 9212 268884 9268
rect 4172 8764 4228 8820
rect 278012 7644 278068 7700
rect 267148 7532 267204 7588
rect 271404 7532 271460 7588
rect 274652 7084 274708 7140
rect 271292 5852 271348 5908
rect 41804 4956 41860 5012
rect 41916 4396 41972 4452
rect 16716 4172 16772 4228
rect 18396 4172 18452 4228
rect 20076 4172 20132 4228
rect 35196 4172 35252 4228
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect 4396 558964 4452 558974
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect 4172 544852 4228 544862
rect 4172 418078 4228 544796
rect 4284 502516 4340 502526
rect 4284 420028 4340 502460
rect 4396 469588 4452 558908
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 4396 469522 4452 469532
rect 4508 516628 4564 516638
rect 4508 467908 4564 516572
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 4508 467842 4564 467852
rect 4620 474292 4676 474302
rect 4620 466228 4676 474236
rect 4620 466162 4676 466172
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect 4508 460180 4564 460190
rect 4284 419972 4452 420028
rect 4172 418022 4340 418078
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect 4172 417844 4228 417854
rect 4172 416818 4228 417788
rect 4172 416752 4228 416762
rect 4284 410698 4340 418022
rect 4284 410632 4340 410642
rect 4396 409438 4452 419972
rect 4396 409372 4452 409382
rect 4508 409258 4564 460124
rect 4508 409192 4564 409202
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect 4284 389620 4340 389630
rect 4060 380278 4116 380288
rect 4060 372988 4116 380222
rect 4284 377188 4340 389564
rect 4284 377122 4340 377132
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 4172 376318 4228 376328
rect 4172 375732 4228 376262
rect 4172 375666 4228 375676
rect 4060 372932 4228 372988
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect 4060 206578 4116 206588
rect 4060 206388 4116 206522
rect 4060 206322 4116 206332
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect 4172 22932 4228 372932
rect 5418 364350 6038 381922
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 36138 562350 36758 579922
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 36138 544350 36758 561922
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 36138 526350 36758 543922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 36138 490350 36758 507922
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 12572 488404 12628 488414
rect 12572 402418 12628 488348
rect 12572 402352 12628 402362
rect 36138 472350 36758 489922
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 36138 454350 36758 471922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 36138 418350 36758 435922
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 4284 347284 4340 347294
rect 4284 313348 4340 347228
rect 4284 313282 4340 313292
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5418 328350 6038 345922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 4284 289268 4340 289278
rect 4284 262836 4340 289212
rect 4284 262770 4340 262780
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 4620 248500 4676 248510
rect 4620 247078 4676 248444
rect 4620 247012 4676 247022
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 4284 210868 4340 210878
rect 4284 178052 4340 210812
rect 4284 177986 4340 177996
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 7532 378838 7588 378848
rect 7532 149940 7588 378782
rect 7532 149874 7588 149884
rect 9138 370350 9758 387922
rect 36138 400350 36758 417922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 20076 384778 20132 384788
rect 18396 383698 18452 383708
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 9138 334350 9758 351922
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 316350 9758 333922
rect 9138 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 9758 316350
rect 9138 316226 9758 316294
rect 9138 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 9758 316226
rect 9138 316102 9758 316170
rect 9138 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 9758 316102
rect 9138 315978 9758 316046
rect 9138 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 9758 315978
rect 9138 298350 9758 315922
rect 9138 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 9758 298350
rect 9138 298226 9758 298294
rect 9138 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 9758 298226
rect 9138 298102 9758 298170
rect 9138 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 9758 298102
rect 9138 297978 9758 298046
rect 9138 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 9758 297978
rect 9138 280350 9758 297922
rect 14252 383338 14308 383348
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 9138 262350 9758 279922
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 4284 79156 4340 79166
rect 4284 55378 4340 79100
rect 4284 55312 4340 55322
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 4172 22866 4228 22876
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 4172 12628 4228 12638
rect 4172 8820 4228 12572
rect 4172 8754 4228 8764
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 4350 6038 21922
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 136350 9758 153922
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 9138 118350 9758 135922
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 9138 100350 9758 117922
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 10892 290276 10948 290286
rect 10892 93492 10948 290220
rect 14252 107380 14308 383282
rect 14252 107314 14308 107324
rect 16716 372178 16772 372188
rect 10892 93426 10948 93436
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 9138 64350 9758 81922
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 9138 10350 9758 27922
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 16716 4228 16772 372122
rect 16716 4162 16772 4172
rect 18396 4228 18452 383642
rect 18396 4162 18452 4172
rect 20076 4228 20132 384722
rect 36138 382350 36758 399922
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 31052 379198 31108 379208
rect 26012 292516 26068 292526
rect 26012 12628 26068 292460
rect 27692 291396 27748 291406
rect 27692 50932 27748 291340
rect 29372 289156 29428 289166
rect 29372 135604 29428 289100
rect 31052 192052 31108 379142
rect 31052 191986 31108 191996
rect 32732 379018 32788 379028
rect 29372 135538 29428 135548
rect 32732 65044 32788 378962
rect 36138 364350 36758 381922
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 36138 346350 36758 363922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 36138 328350 36758 345922
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 36138 310350 36758 327922
rect 36138 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 36758 310350
rect 36138 310226 36758 310294
rect 36138 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 36758 310226
rect 36138 310102 36758 310170
rect 36138 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 36758 310102
rect 36138 309978 36758 310046
rect 36138 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 36758 309978
rect 36138 292350 36758 309922
rect 36138 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 36758 292350
rect 36138 292226 36758 292294
rect 36138 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 36758 292226
rect 36138 292102 36758 292170
rect 36138 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 36758 292102
rect 36138 291978 36758 292046
rect 36138 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 36758 291978
rect 36138 274350 36758 291922
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 36138 256350 36758 273922
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 36138 238350 36758 255922
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 32732 64978 32788 64988
rect 35196 229258 35252 229268
rect 27692 50866 27748 50876
rect 26012 12562 26068 12572
rect 20076 4162 20132 4172
rect 35196 4228 35252 229202
rect 35196 4162 35252 4172
rect 36138 220350 36758 237922
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 36138 202350 36758 219922
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568350 40478 585922
rect 39858 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 40478 568350
rect 39858 568226 40478 568294
rect 39858 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 40478 568226
rect 39858 568102 40478 568170
rect 39858 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 40478 568102
rect 39858 567978 40478 568046
rect 39858 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 40478 567978
rect 39858 550350 40478 567922
rect 39858 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 40478 550350
rect 39858 550226 40478 550294
rect 39858 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 40478 550226
rect 39858 550102 40478 550170
rect 39858 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 40478 550102
rect 39858 549978 40478 550046
rect 39858 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 40478 549978
rect 39858 532350 40478 549922
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 66858 535792 67478 543922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 539752 71198 549922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 562350 98198 579922
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 97578 549832 98198 561922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 568350 101918 585922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 130324 580063 130796 580120
rect 130324 580007 130346 580063
rect 130402 580007 130470 580063
rect 130526 580007 130594 580063
rect 130650 580007 130718 580063
rect 130774 580007 130796 580063
rect 130324 579939 130796 580007
rect 130324 579883 130346 579939
rect 130402 579883 130470 579939
rect 130526 579883 130594 579939
rect 130650 579883 130718 579939
rect 130774 579883 130796 579939
rect 130324 579826 130796 579883
rect 132018 578452 132638 585922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 101298 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 101918 568350
rect 101298 568226 101918 568294
rect 101298 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 101918 568226
rect 101298 568102 101918 568170
rect 101298 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 101918 568102
rect 101298 567978 101918 568046
rect 101298 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 101918 567978
rect 101298 550350 101918 567922
rect 159018 562350 159638 579922
rect 116160 562272 132720 562300
rect 116160 562216 116228 562272
rect 116284 562216 116352 562272
rect 116408 562216 116476 562272
rect 116532 562216 116600 562272
rect 116656 562216 116724 562272
rect 116780 562216 116848 562272
rect 116904 562216 116972 562272
rect 117028 562216 117096 562272
rect 117152 562216 117220 562272
rect 117276 562216 117344 562272
rect 117400 562216 117468 562272
rect 117524 562216 117592 562272
rect 117648 562216 117716 562272
rect 117772 562216 117840 562272
rect 117896 562216 117964 562272
rect 118020 562216 118088 562272
rect 118144 562216 118212 562272
rect 118268 562216 118336 562272
rect 118392 562216 118460 562272
rect 118516 562216 118584 562272
rect 118640 562216 118708 562272
rect 118764 562216 118832 562272
rect 118888 562216 118956 562272
rect 119012 562216 119080 562272
rect 119136 562216 119204 562272
rect 119260 562216 119328 562272
rect 119384 562216 119452 562272
rect 119508 562216 119576 562272
rect 119632 562216 119700 562272
rect 119756 562216 119824 562272
rect 119880 562216 119948 562272
rect 120004 562216 120072 562272
rect 120128 562216 120196 562272
rect 120252 562216 120320 562272
rect 120376 562216 120444 562272
rect 120500 562216 120568 562272
rect 120624 562216 120692 562272
rect 120748 562216 120816 562272
rect 120872 562216 120940 562272
rect 120996 562216 121064 562272
rect 121120 562216 121188 562272
rect 121244 562216 121312 562272
rect 121368 562216 121436 562272
rect 121492 562216 121560 562272
rect 121616 562216 121684 562272
rect 121740 562216 121808 562272
rect 121864 562216 121932 562272
rect 121988 562216 122056 562272
rect 122112 562216 122180 562272
rect 122236 562216 122304 562272
rect 122360 562216 122428 562272
rect 122484 562216 122552 562272
rect 122608 562216 122676 562272
rect 122732 562216 122800 562272
rect 122856 562216 122924 562272
rect 122980 562216 123048 562272
rect 123104 562216 123172 562272
rect 123228 562216 123296 562272
rect 123352 562216 123420 562272
rect 123476 562216 123544 562272
rect 123600 562216 123668 562272
rect 123724 562216 123792 562272
rect 123848 562216 123916 562272
rect 123972 562216 124040 562272
rect 124096 562216 124164 562272
rect 124220 562216 124288 562272
rect 124344 562216 124412 562272
rect 124468 562216 124536 562272
rect 124592 562216 124660 562272
rect 124716 562216 124784 562272
rect 124840 562216 124908 562272
rect 124964 562216 125032 562272
rect 125088 562216 125156 562272
rect 125212 562216 125280 562272
rect 125336 562216 125404 562272
rect 125460 562216 125528 562272
rect 125584 562216 125652 562272
rect 125708 562216 125776 562272
rect 125832 562216 125900 562272
rect 125956 562216 126024 562272
rect 126080 562216 126148 562272
rect 126204 562216 126272 562272
rect 126328 562216 126396 562272
rect 126452 562216 126520 562272
rect 126576 562216 126644 562272
rect 126700 562216 126768 562272
rect 126824 562216 126892 562272
rect 126948 562216 127016 562272
rect 127072 562216 127140 562272
rect 127196 562216 127264 562272
rect 127320 562216 127388 562272
rect 127444 562216 127512 562272
rect 127568 562216 127636 562272
rect 127692 562216 127760 562272
rect 127816 562216 127884 562272
rect 127940 562216 128008 562272
rect 128064 562216 128132 562272
rect 128188 562216 128256 562272
rect 128312 562216 128380 562272
rect 128436 562216 128504 562272
rect 128560 562216 128628 562272
rect 128684 562216 128752 562272
rect 128808 562216 128876 562272
rect 128932 562216 129000 562272
rect 129056 562216 129124 562272
rect 129180 562216 129248 562272
rect 129304 562216 129372 562272
rect 129428 562216 129496 562272
rect 129552 562216 129620 562272
rect 129676 562216 129744 562272
rect 129800 562216 129868 562272
rect 129924 562216 129992 562272
rect 130048 562216 130116 562272
rect 130172 562216 130240 562272
rect 130296 562216 130364 562272
rect 130420 562216 130488 562272
rect 130544 562216 130612 562272
rect 130668 562216 130736 562272
rect 130792 562216 130860 562272
rect 130916 562216 130984 562272
rect 131040 562216 131108 562272
rect 131164 562216 131232 562272
rect 131288 562216 131356 562272
rect 131412 562216 131480 562272
rect 131536 562216 131604 562272
rect 131660 562216 131728 562272
rect 131784 562216 131852 562272
rect 131908 562216 131976 562272
rect 132032 562216 132100 562272
rect 132156 562216 132224 562272
rect 132280 562216 132348 562272
rect 132404 562216 132472 562272
rect 132528 562216 132596 562272
rect 132652 562216 132720 562272
rect 116160 562148 132720 562216
rect 116160 562092 116228 562148
rect 116284 562092 116352 562148
rect 116408 562092 116476 562148
rect 116532 562092 116600 562148
rect 116656 562092 116724 562148
rect 116780 562092 116848 562148
rect 116904 562092 116972 562148
rect 117028 562092 117096 562148
rect 117152 562092 117220 562148
rect 117276 562092 117344 562148
rect 117400 562092 117468 562148
rect 117524 562092 117592 562148
rect 117648 562092 117716 562148
rect 117772 562092 117840 562148
rect 117896 562092 117964 562148
rect 118020 562092 118088 562148
rect 118144 562092 118212 562148
rect 118268 562092 118336 562148
rect 118392 562092 118460 562148
rect 118516 562092 118584 562148
rect 118640 562092 118708 562148
rect 118764 562092 118832 562148
rect 118888 562092 118956 562148
rect 119012 562092 119080 562148
rect 119136 562092 119204 562148
rect 119260 562092 119328 562148
rect 119384 562092 119452 562148
rect 119508 562092 119576 562148
rect 119632 562092 119700 562148
rect 119756 562092 119824 562148
rect 119880 562092 119948 562148
rect 120004 562092 120072 562148
rect 120128 562092 120196 562148
rect 120252 562092 120320 562148
rect 120376 562092 120444 562148
rect 120500 562092 120568 562148
rect 120624 562092 120692 562148
rect 120748 562092 120816 562148
rect 120872 562092 120940 562148
rect 120996 562092 121064 562148
rect 121120 562092 121188 562148
rect 121244 562092 121312 562148
rect 121368 562092 121436 562148
rect 121492 562092 121560 562148
rect 121616 562092 121684 562148
rect 121740 562092 121808 562148
rect 121864 562092 121932 562148
rect 121988 562092 122056 562148
rect 122112 562092 122180 562148
rect 122236 562092 122304 562148
rect 122360 562092 122428 562148
rect 122484 562092 122552 562148
rect 122608 562092 122676 562148
rect 122732 562092 122800 562148
rect 122856 562092 122924 562148
rect 122980 562092 123048 562148
rect 123104 562092 123172 562148
rect 123228 562092 123296 562148
rect 123352 562092 123420 562148
rect 123476 562092 123544 562148
rect 123600 562092 123668 562148
rect 123724 562092 123792 562148
rect 123848 562092 123916 562148
rect 123972 562092 124040 562148
rect 124096 562092 124164 562148
rect 124220 562092 124288 562148
rect 124344 562092 124412 562148
rect 124468 562092 124536 562148
rect 124592 562092 124660 562148
rect 124716 562092 124784 562148
rect 124840 562092 124908 562148
rect 124964 562092 125032 562148
rect 125088 562092 125156 562148
rect 125212 562092 125280 562148
rect 125336 562092 125404 562148
rect 125460 562092 125528 562148
rect 125584 562092 125652 562148
rect 125708 562092 125776 562148
rect 125832 562092 125900 562148
rect 125956 562092 126024 562148
rect 126080 562092 126148 562148
rect 126204 562092 126272 562148
rect 126328 562092 126396 562148
rect 126452 562092 126520 562148
rect 126576 562092 126644 562148
rect 126700 562092 126768 562148
rect 126824 562092 126892 562148
rect 126948 562092 127016 562148
rect 127072 562092 127140 562148
rect 127196 562092 127264 562148
rect 127320 562092 127388 562148
rect 127444 562092 127512 562148
rect 127568 562092 127636 562148
rect 127692 562092 127760 562148
rect 127816 562092 127884 562148
rect 127940 562092 128008 562148
rect 128064 562092 128132 562148
rect 128188 562092 128256 562148
rect 128312 562092 128380 562148
rect 128436 562092 128504 562148
rect 128560 562092 128628 562148
rect 128684 562092 128752 562148
rect 128808 562092 128876 562148
rect 128932 562092 129000 562148
rect 129056 562092 129124 562148
rect 129180 562092 129248 562148
rect 129304 562092 129372 562148
rect 129428 562092 129496 562148
rect 129552 562092 129620 562148
rect 129676 562092 129744 562148
rect 129800 562092 129868 562148
rect 129924 562092 129992 562148
rect 130048 562092 130116 562148
rect 130172 562092 130240 562148
rect 130296 562092 130364 562148
rect 130420 562092 130488 562148
rect 130544 562092 130612 562148
rect 130668 562092 130736 562148
rect 130792 562092 130860 562148
rect 130916 562092 130984 562148
rect 131040 562092 131108 562148
rect 131164 562092 131232 562148
rect 131288 562092 131356 562148
rect 131412 562092 131480 562148
rect 131536 562092 131604 562148
rect 131660 562092 131728 562148
rect 131784 562092 131852 562148
rect 131908 562092 131976 562148
rect 132032 562092 132100 562148
rect 132156 562092 132224 562148
rect 132280 562092 132348 562148
rect 132404 562092 132472 562148
rect 132528 562092 132596 562148
rect 132652 562092 132720 562148
rect 116160 562024 132720 562092
rect 116160 561968 116228 562024
rect 116284 561968 116352 562024
rect 116408 561968 116476 562024
rect 116532 561968 116600 562024
rect 116656 561968 116724 562024
rect 116780 561968 116848 562024
rect 116904 561968 116972 562024
rect 117028 561968 117096 562024
rect 117152 561968 117220 562024
rect 117276 561968 117344 562024
rect 117400 561968 117468 562024
rect 117524 561968 117592 562024
rect 117648 561968 117716 562024
rect 117772 561968 117840 562024
rect 117896 561968 117964 562024
rect 118020 561968 118088 562024
rect 118144 561968 118212 562024
rect 118268 561968 118336 562024
rect 118392 561968 118460 562024
rect 118516 561968 118584 562024
rect 118640 561968 118708 562024
rect 118764 561968 118832 562024
rect 118888 561968 118956 562024
rect 119012 561968 119080 562024
rect 119136 561968 119204 562024
rect 119260 561968 119328 562024
rect 119384 561968 119452 562024
rect 119508 561968 119576 562024
rect 119632 561968 119700 562024
rect 119756 561968 119824 562024
rect 119880 561968 119948 562024
rect 120004 561968 120072 562024
rect 120128 561968 120196 562024
rect 120252 561968 120320 562024
rect 120376 561968 120444 562024
rect 120500 561968 120568 562024
rect 120624 561968 120692 562024
rect 120748 561968 120816 562024
rect 120872 561968 120940 562024
rect 120996 561968 121064 562024
rect 121120 561968 121188 562024
rect 121244 561968 121312 562024
rect 121368 561968 121436 562024
rect 121492 561968 121560 562024
rect 121616 561968 121684 562024
rect 121740 561968 121808 562024
rect 121864 561968 121932 562024
rect 121988 561968 122056 562024
rect 122112 561968 122180 562024
rect 122236 561968 122304 562024
rect 122360 561968 122428 562024
rect 122484 561968 122552 562024
rect 122608 561968 122676 562024
rect 122732 561968 122800 562024
rect 122856 561968 122924 562024
rect 122980 561968 123048 562024
rect 123104 561968 123172 562024
rect 123228 561968 123296 562024
rect 123352 561968 123420 562024
rect 123476 561968 123544 562024
rect 123600 561968 123668 562024
rect 123724 561968 123792 562024
rect 123848 561968 123916 562024
rect 123972 561968 124040 562024
rect 124096 561968 124164 562024
rect 124220 561968 124288 562024
rect 124344 561968 124412 562024
rect 124468 561968 124536 562024
rect 124592 561968 124660 562024
rect 124716 561968 124784 562024
rect 124840 561968 124908 562024
rect 124964 561968 125032 562024
rect 125088 561968 125156 562024
rect 125212 561968 125280 562024
rect 125336 561968 125404 562024
rect 125460 561968 125528 562024
rect 125584 561968 125652 562024
rect 125708 561968 125776 562024
rect 125832 561968 125900 562024
rect 125956 561968 126024 562024
rect 126080 561968 126148 562024
rect 126204 561968 126272 562024
rect 126328 561968 126396 562024
rect 126452 561968 126520 562024
rect 126576 561968 126644 562024
rect 126700 561968 126768 562024
rect 126824 561968 126892 562024
rect 126948 561968 127016 562024
rect 127072 561968 127140 562024
rect 127196 561968 127264 562024
rect 127320 561968 127388 562024
rect 127444 561968 127512 562024
rect 127568 561968 127636 562024
rect 127692 561968 127760 562024
rect 127816 561968 127884 562024
rect 127940 561968 128008 562024
rect 128064 561968 128132 562024
rect 128188 561968 128256 562024
rect 128312 561968 128380 562024
rect 128436 561968 128504 562024
rect 128560 561968 128628 562024
rect 128684 561968 128752 562024
rect 128808 561968 128876 562024
rect 128932 561968 129000 562024
rect 129056 561968 129124 562024
rect 129180 561968 129248 562024
rect 129304 561968 129372 562024
rect 129428 561968 129496 562024
rect 129552 561968 129620 562024
rect 129676 561968 129744 562024
rect 129800 561968 129868 562024
rect 129924 561968 129992 562024
rect 130048 561968 130116 562024
rect 130172 561968 130240 562024
rect 130296 561968 130364 562024
rect 130420 561968 130488 562024
rect 130544 561968 130612 562024
rect 130668 561968 130736 562024
rect 130792 561968 130860 562024
rect 130916 561968 130984 562024
rect 131040 561968 131108 562024
rect 131164 561968 131232 562024
rect 131288 561968 131356 562024
rect 131412 561968 131480 562024
rect 131536 561968 131604 562024
rect 131660 561968 131728 562024
rect 131784 561968 131852 562024
rect 131908 561968 131976 562024
rect 132032 561968 132100 562024
rect 132156 561968 132224 562024
rect 132280 561968 132348 562024
rect 132404 561968 132472 562024
rect 132528 561968 132596 562024
rect 132652 561968 132720 562024
rect 116160 561940 132720 561968
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 101298 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 101918 550350
rect 101298 550226 101918 550294
rect 101298 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 101918 550226
rect 101298 550102 101918 550170
rect 101298 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 101918 550102
rect 101298 549978 101918 550046
rect 101298 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 101918 549978
rect 101298 549472 101918 549922
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 159018 544350 159638 561922
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 104280 544058 126420 544120
rect 104280 544002 104348 544058
rect 104404 544002 104472 544058
rect 104528 544002 104596 544058
rect 104652 544002 104720 544058
rect 104776 544002 104844 544058
rect 104900 544002 104968 544058
rect 105024 544002 105092 544058
rect 105148 544002 105216 544058
rect 105272 544002 105340 544058
rect 105396 544002 105464 544058
rect 105520 544002 105588 544058
rect 105644 544002 105712 544058
rect 105768 544002 105836 544058
rect 105892 544002 105960 544058
rect 106016 544002 106084 544058
rect 106140 544002 106208 544058
rect 106264 544002 106332 544058
rect 106388 544002 106456 544058
rect 106512 544002 106580 544058
rect 106636 544002 106704 544058
rect 106760 544002 106828 544058
rect 106884 544002 106952 544058
rect 107008 544002 107076 544058
rect 107132 544002 107200 544058
rect 107256 544002 107324 544058
rect 107380 544002 107448 544058
rect 107504 544002 107572 544058
rect 107628 544002 107696 544058
rect 107752 544002 107820 544058
rect 107876 544002 107944 544058
rect 108000 544002 108068 544058
rect 108124 544002 108192 544058
rect 108248 544002 108316 544058
rect 108372 544002 108440 544058
rect 108496 544002 108564 544058
rect 108620 544002 108688 544058
rect 108744 544002 108812 544058
rect 108868 544002 108936 544058
rect 108992 544002 109060 544058
rect 109116 544002 109184 544058
rect 109240 544002 109308 544058
rect 109364 544002 109432 544058
rect 109488 544002 109556 544058
rect 109612 544002 109680 544058
rect 109736 544002 109804 544058
rect 109860 544002 109928 544058
rect 109984 544002 110052 544058
rect 110108 544002 110176 544058
rect 110232 544002 110300 544058
rect 110356 544002 110424 544058
rect 110480 544002 110548 544058
rect 110604 544002 110672 544058
rect 110728 544002 110796 544058
rect 110852 544002 110920 544058
rect 110976 544002 111044 544058
rect 111100 544002 111168 544058
rect 111224 544002 111292 544058
rect 111348 544002 111416 544058
rect 111472 544002 111540 544058
rect 111596 544002 111664 544058
rect 111720 544002 111788 544058
rect 111844 544002 111912 544058
rect 111968 544002 112036 544058
rect 112092 544002 112160 544058
rect 112216 544002 112284 544058
rect 112340 544002 112408 544058
rect 112464 544002 112532 544058
rect 112588 544002 112656 544058
rect 112712 544002 112780 544058
rect 112836 544002 112904 544058
rect 112960 544002 113028 544058
rect 113084 544002 113152 544058
rect 113208 544002 113276 544058
rect 113332 544002 113400 544058
rect 113456 544002 113524 544058
rect 113580 544002 113648 544058
rect 113704 544002 113772 544058
rect 113828 544002 113896 544058
rect 113952 544002 114020 544058
rect 114076 544002 114144 544058
rect 114200 544002 114268 544058
rect 114324 544002 114392 544058
rect 114448 544002 114516 544058
rect 114572 544002 114640 544058
rect 114696 544002 114764 544058
rect 114820 544002 114888 544058
rect 114944 544002 115012 544058
rect 115068 544002 115136 544058
rect 115192 544002 115260 544058
rect 115316 544002 115384 544058
rect 115440 544002 115508 544058
rect 115564 544002 115632 544058
rect 115688 544002 115756 544058
rect 115812 544002 115880 544058
rect 115936 544002 116004 544058
rect 116060 544002 116128 544058
rect 116184 544002 116252 544058
rect 116308 544002 116376 544058
rect 116432 544002 116500 544058
rect 116556 544002 116624 544058
rect 116680 544002 116748 544058
rect 116804 544002 116872 544058
rect 116928 544002 116996 544058
rect 117052 544002 117120 544058
rect 117176 544002 117244 544058
rect 117300 544002 117368 544058
rect 117424 544002 117492 544058
rect 117548 544002 117616 544058
rect 117672 544002 117740 544058
rect 117796 544002 117864 544058
rect 117920 544002 117988 544058
rect 118044 544002 118112 544058
rect 118168 544002 118236 544058
rect 118292 544002 118360 544058
rect 118416 544002 118484 544058
rect 118540 544002 118608 544058
rect 118664 544002 118732 544058
rect 118788 544002 118856 544058
rect 118912 544002 118980 544058
rect 119036 544002 119104 544058
rect 119160 544002 119228 544058
rect 119284 544002 119352 544058
rect 119408 544002 119476 544058
rect 119532 544002 119600 544058
rect 119656 544002 119724 544058
rect 119780 544002 119848 544058
rect 119904 544002 119972 544058
rect 120028 544002 120096 544058
rect 120152 544002 120220 544058
rect 120276 544002 120344 544058
rect 120400 544002 120468 544058
rect 120524 544002 120592 544058
rect 120648 544002 120716 544058
rect 120772 544002 120840 544058
rect 120896 544002 120964 544058
rect 121020 544002 121088 544058
rect 121144 544002 121212 544058
rect 121268 544002 121336 544058
rect 121392 544002 121460 544058
rect 121516 544002 121584 544058
rect 121640 544002 121708 544058
rect 121764 544002 121832 544058
rect 121888 544002 121956 544058
rect 122012 544002 122080 544058
rect 122136 544002 122204 544058
rect 122260 544002 122328 544058
rect 122384 544002 122452 544058
rect 122508 544002 122576 544058
rect 122632 544002 122700 544058
rect 122756 544002 122824 544058
rect 122880 544002 122948 544058
rect 123004 544002 123072 544058
rect 123128 544002 123196 544058
rect 123252 544002 123320 544058
rect 123376 544002 123444 544058
rect 123500 544002 123568 544058
rect 123624 544002 123692 544058
rect 123748 544002 123816 544058
rect 123872 544002 123940 544058
rect 123996 544002 124064 544058
rect 124120 544002 124188 544058
rect 124244 544002 124312 544058
rect 124368 544002 124436 544058
rect 124492 544002 124560 544058
rect 124616 544002 124684 544058
rect 124740 544002 124808 544058
rect 124864 544002 124932 544058
rect 124988 544002 125056 544058
rect 125112 544002 125180 544058
rect 125236 544002 125304 544058
rect 125360 544002 125428 544058
rect 125484 544002 125552 544058
rect 125608 544002 125676 544058
rect 125732 544002 125800 544058
rect 125856 544002 125924 544058
rect 125980 544002 126048 544058
rect 126104 544002 126172 544058
rect 126228 544002 126296 544058
rect 126352 544002 126420 544058
rect 104280 543940 126420 544002
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 39858 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 40478 532350
rect 39858 532226 40478 532294
rect 66660 532358 74760 532420
rect 66660 532302 66714 532358
rect 66770 532302 66838 532358
rect 66894 532302 66962 532358
rect 67018 532302 67086 532358
rect 67142 532302 67210 532358
rect 67266 532302 67334 532358
rect 67390 532302 67458 532358
rect 67514 532302 67582 532358
rect 67638 532302 67706 532358
rect 67762 532302 67830 532358
rect 67886 532302 67954 532358
rect 68010 532302 68078 532358
rect 68134 532302 68202 532358
rect 68258 532302 68326 532358
rect 68382 532302 68450 532358
rect 68506 532302 68574 532358
rect 68630 532302 68698 532358
rect 68754 532302 68822 532358
rect 68878 532302 68946 532358
rect 69002 532302 69070 532358
rect 69126 532302 69194 532358
rect 69250 532302 69318 532358
rect 69374 532302 69442 532358
rect 69498 532302 69566 532358
rect 69622 532302 69690 532358
rect 69746 532302 69814 532358
rect 69870 532302 69938 532358
rect 69994 532302 70062 532358
rect 70118 532302 70186 532358
rect 70242 532302 70310 532358
rect 70366 532302 70434 532358
rect 70490 532302 70558 532358
rect 70614 532302 70682 532358
rect 70738 532302 70806 532358
rect 70862 532302 70930 532358
rect 70986 532302 71054 532358
rect 71110 532302 71178 532358
rect 71234 532302 71302 532358
rect 71358 532302 71426 532358
rect 71482 532302 71550 532358
rect 71606 532302 71674 532358
rect 71730 532302 71798 532358
rect 71854 532302 71922 532358
rect 71978 532302 72046 532358
rect 72102 532302 72170 532358
rect 72226 532302 72294 532358
rect 72350 532302 72418 532358
rect 72474 532302 72542 532358
rect 72598 532302 72666 532358
rect 72722 532302 72790 532358
rect 72846 532302 72914 532358
rect 72970 532302 73038 532358
rect 73094 532302 73162 532358
rect 73218 532302 73286 532358
rect 73342 532302 73410 532358
rect 73466 532302 73534 532358
rect 73590 532302 73658 532358
rect 73714 532302 73782 532358
rect 73838 532302 73906 532358
rect 73962 532302 74030 532358
rect 74086 532302 74154 532358
rect 74210 532302 74278 532358
rect 74334 532302 74402 532358
rect 74458 532302 74526 532358
rect 74582 532302 74650 532358
rect 74706 532302 74760 532358
rect 66660 532240 74760 532302
rect 39858 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 40478 532226
rect 39858 532102 40478 532170
rect 39858 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 40478 532102
rect 39858 531978 40478 532046
rect 39858 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 40478 531978
rect 39858 514350 40478 531922
rect 66480 531998 66960 532060
rect 66480 531942 66506 531998
rect 66562 531942 66630 531998
rect 66686 531942 66754 531998
rect 66810 531942 66878 531998
rect 66934 531942 66960 531998
rect 66480 531880 66960 531942
rect 66976 531998 67456 532060
rect 66976 531942 67002 531998
rect 67058 531942 67126 531998
rect 67182 531942 67250 531998
rect 67306 531942 67374 531998
rect 67430 531942 67456 531998
rect 66976 531880 67456 531942
rect 67472 531998 67952 532060
rect 67472 531942 67498 531998
rect 67554 531942 67622 531998
rect 67678 531942 67746 531998
rect 67802 531942 67870 531998
rect 67926 531942 67952 531998
rect 67472 531880 67952 531942
rect 67968 531998 68448 532060
rect 67968 531942 67994 531998
rect 68050 531942 68118 531998
rect 68174 531942 68242 531998
rect 68298 531942 68366 531998
rect 68422 531942 68448 531998
rect 67968 531880 68448 531942
rect 68464 531998 68944 532060
rect 68464 531942 68490 531998
rect 68546 531942 68614 531998
rect 68670 531942 68738 531998
rect 68794 531942 68862 531998
rect 68918 531942 68944 531998
rect 68464 531880 68944 531942
rect 68960 531998 69440 532060
rect 68960 531942 68986 531998
rect 69042 531942 69110 531998
rect 69166 531942 69234 531998
rect 69290 531942 69358 531998
rect 69414 531942 69440 531998
rect 68960 531880 69440 531942
rect 69456 531998 69936 532060
rect 69456 531942 69482 531998
rect 69538 531942 69606 531998
rect 69662 531942 69730 531998
rect 69786 531942 69854 531998
rect 69910 531942 69936 531998
rect 69456 531880 69936 531942
rect 69952 531998 70432 532060
rect 69952 531942 69978 531998
rect 70034 531942 70102 531998
rect 70158 531942 70226 531998
rect 70282 531942 70350 531998
rect 70406 531942 70432 531998
rect 69952 531880 70432 531942
rect 70448 531998 70928 532060
rect 70448 531942 70474 531998
rect 70530 531942 70598 531998
rect 70654 531942 70722 531998
rect 70778 531942 70846 531998
rect 70902 531942 70928 531998
rect 70448 531880 70928 531942
rect 70944 531998 71424 532060
rect 70944 531942 70970 531998
rect 71026 531942 71094 531998
rect 71150 531942 71218 531998
rect 71274 531942 71342 531998
rect 71398 531942 71424 531998
rect 70944 531880 71424 531942
rect 71440 531998 71920 532060
rect 71440 531942 71466 531998
rect 71522 531942 71590 531998
rect 71646 531942 71714 531998
rect 71770 531942 71838 531998
rect 71894 531942 71920 531998
rect 71440 531880 71920 531942
rect 71936 531998 72416 532060
rect 71936 531942 71962 531998
rect 72018 531942 72086 531998
rect 72142 531942 72210 531998
rect 72266 531942 72334 531998
rect 72390 531942 72416 531998
rect 71936 531880 72416 531942
rect 72432 531998 72912 532060
rect 72432 531942 72458 531998
rect 72514 531942 72582 531998
rect 72638 531942 72706 531998
rect 72762 531942 72830 531998
rect 72886 531942 72912 531998
rect 72432 531880 72912 531942
rect 72928 531998 73408 532060
rect 72928 531942 72954 531998
rect 73010 531942 73078 531998
rect 73134 531942 73202 531998
rect 73258 531942 73326 531998
rect 73382 531942 73408 531998
rect 72928 531880 73408 531942
rect 73424 531998 73904 532060
rect 73424 531942 73450 531998
rect 73506 531942 73574 531998
rect 73630 531942 73698 531998
rect 73754 531942 73822 531998
rect 73878 531942 73904 531998
rect 73424 531880 73904 531942
rect 73920 531998 74400 532060
rect 73920 531942 73946 531998
rect 74002 531942 74070 531998
rect 74126 531942 74194 531998
rect 74250 531942 74318 531998
rect 74374 531942 74400 531998
rect 73920 531880 74400 531942
rect 39858 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 40478 514350
rect 39858 514226 40478 514294
rect 39858 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 40478 514226
rect 39858 514102 40478 514170
rect 39858 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 40478 514102
rect 39858 513978 40478 514046
rect 39858 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 40478 513978
rect 39858 496350 40478 513922
rect 39858 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 40478 496350
rect 39858 496226 40478 496294
rect 39858 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 40478 496226
rect 39858 496102 40478 496170
rect 39858 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 40478 496102
rect 39858 495978 40478 496046
rect 39858 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 40478 495978
rect 39858 478350 40478 495922
rect 39858 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 40478 478350
rect 39858 478226 40478 478294
rect 39858 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 40478 478226
rect 39858 478102 40478 478170
rect 39858 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 40478 478102
rect 39858 477978 40478 478046
rect 39858 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 40478 477978
rect 39858 460350 40478 477922
rect 39858 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 40478 460350
rect 39858 460226 40478 460294
rect 39858 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 40478 460226
rect 39858 460102 40478 460170
rect 39858 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 40478 460102
rect 39858 459978 40478 460046
rect 39858 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 40478 459978
rect 39858 442350 40478 459922
rect 39858 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 40478 442350
rect 39858 442226 40478 442294
rect 39858 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 40478 442226
rect 39858 442102 40478 442170
rect 39858 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 40478 442102
rect 39858 441978 40478 442046
rect 39858 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 40478 441978
rect 39858 424350 40478 441922
rect 39858 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 40478 424350
rect 39858 424226 40478 424294
rect 39858 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 40478 424226
rect 39858 424102 40478 424170
rect 39858 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 40478 424102
rect 39858 423978 40478 424046
rect 39858 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 40478 423978
rect 39858 406350 40478 423922
rect 39858 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 40478 406350
rect 39858 406226 40478 406294
rect 39858 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 40478 406226
rect 39858 406102 40478 406170
rect 39858 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 40478 406102
rect 39858 405978 40478 406046
rect 39858 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 40478 405978
rect 39858 388350 40478 405922
rect 57932 530740 57988 530750
rect 57932 404038 57988 530684
rect 159018 526350 159638 543922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 95820 526058 96052 526120
rect 95820 526002 95846 526058
rect 95902 526002 95970 526058
rect 96026 526002 96052 526058
rect 95820 525940 96052 526002
rect 96068 526058 96548 526120
rect 96068 526002 96094 526058
rect 96150 526002 96218 526058
rect 96274 526002 96342 526058
rect 96398 526002 96466 526058
rect 96522 526002 96548 526058
rect 96068 525940 96548 526002
rect 96564 526058 97044 526120
rect 96564 526002 96590 526058
rect 96646 526002 96714 526058
rect 96770 526002 96838 526058
rect 96894 526002 96962 526058
rect 97018 526002 97044 526058
rect 96564 525940 97044 526002
rect 97060 526058 97540 526120
rect 97060 526002 97086 526058
rect 97142 526002 97210 526058
rect 97266 526002 97334 526058
rect 97390 526002 97458 526058
rect 97514 526002 97540 526058
rect 97060 525940 97540 526002
rect 97556 526058 98036 526120
rect 97556 526002 97582 526058
rect 97638 526002 97706 526058
rect 97762 526002 97830 526058
rect 97886 526002 97954 526058
rect 98010 526002 98036 526058
rect 97556 525940 98036 526002
rect 98052 526058 98532 526120
rect 98052 526002 98078 526058
rect 98134 526002 98202 526058
rect 98258 526002 98326 526058
rect 98382 526002 98450 526058
rect 98506 526002 98532 526058
rect 98052 525940 98532 526002
rect 98548 526058 99028 526120
rect 98548 526002 98574 526058
rect 98630 526002 98698 526058
rect 98754 526002 98822 526058
rect 98878 526002 98946 526058
rect 99002 526002 99028 526058
rect 98548 525940 99028 526002
rect 99044 526058 99524 526120
rect 99044 526002 99070 526058
rect 99126 526002 99194 526058
rect 99250 526002 99318 526058
rect 99374 526002 99442 526058
rect 99498 526002 99524 526058
rect 99044 525940 99524 526002
rect 99540 526058 100020 526120
rect 99540 526002 99566 526058
rect 99622 526002 99690 526058
rect 99746 526002 99814 526058
rect 99870 526002 99938 526058
rect 99994 526002 100020 526058
rect 99540 525940 100020 526002
rect 100036 526058 100516 526120
rect 100036 526002 100062 526058
rect 100118 526002 100186 526058
rect 100242 526002 100310 526058
rect 100366 526002 100434 526058
rect 100490 526002 100516 526058
rect 100036 525940 100516 526002
rect 100532 526058 101012 526120
rect 100532 526002 100558 526058
rect 100614 526002 100682 526058
rect 100738 526002 100806 526058
rect 100862 526002 100930 526058
rect 100986 526002 101012 526058
rect 100532 525940 101012 526002
rect 101028 526058 101508 526120
rect 101028 526002 101054 526058
rect 101110 526002 101178 526058
rect 101234 526002 101302 526058
rect 101358 526002 101426 526058
rect 101482 526002 101508 526058
rect 101028 525940 101508 526002
rect 101524 526058 102004 526120
rect 101524 526002 101550 526058
rect 101606 526002 101674 526058
rect 101730 526002 101798 526058
rect 101854 526002 101922 526058
rect 101978 526002 102004 526058
rect 101524 525940 102004 526002
rect 102020 526058 102500 526120
rect 102020 526002 102046 526058
rect 102102 526002 102170 526058
rect 102226 526002 102294 526058
rect 102350 526002 102418 526058
rect 102474 526002 102500 526058
rect 102020 525940 102500 526002
rect 102516 526058 102996 526120
rect 102516 526002 102542 526058
rect 102598 526002 102666 526058
rect 102722 526002 102790 526058
rect 102846 526002 102914 526058
rect 102970 526002 102996 526058
rect 102516 525940 102996 526002
rect 103012 526058 103492 526120
rect 103012 526002 103038 526058
rect 103094 526002 103162 526058
rect 103218 526002 103286 526058
rect 103342 526002 103410 526058
rect 103466 526002 103492 526058
rect 103012 525940 103492 526002
rect 103508 526058 103988 526120
rect 103508 526002 103534 526058
rect 103590 526002 103658 526058
rect 103714 526002 103782 526058
rect 103838 526002 103906 526058
rect 103962 526002 103988 526058
rect 103508 525940 103988 526002
rect 104004 526058 104484 526120
rect 104004 526002 104030 526058
rect 104086 526002 104154 526058
rect 104210 526002 104278 526058
rect 104334 526002 104402 526058
rect 104458 526002 104484 526058
rect 104004 525940 104484 526002
rect 104500 526058 104980 526120
rect 104500 526002 104526 526058
rect 104582 526002 104650 526058
rect 104706 526002 104774 526058
rect 104830 526002 104898 526058
rect 104954 526002 104980 526058
rect 104500 525940 104980 526002
rect 104996 526058 105476 526120
rect 104996 526002 105022 526058
rect 105078 526002 105146 526058
rect 105202 526002 105270 526058
rect 105326 526002 105394 526058
rect 105450 526002 105476 526058
rect 104996 525940 105476 526002
rect 105492 526058 105972 526120
rect 105492 526002 105518 526058
rect 105574 526002 105642 526058
rect 105698 526002 105766 526058
rect 105822 526002 105890 526058
rect 105946 526002 105972 526058
rect 105492 525940 105972 526002
rect 105988 526058 106468 526120
rect 105988 526002 106014 526058
rect 106070 526002 106138 526058
rect 106194 526002 106262 526058
rect 106318 526002 106386 526058
rect 106442 526002 106468 526058
rect 105988 525940 106468 526002
rect 106484 526058 106964 526120
rect 106484 526002 106510 526058
rect 106566 526002 106634 526058
rect 106690 526002 106758 526058
rect 106814 526002 106882 526058
rect 106938 526002 106964 526058
rect 106484 525940 106964 526002
rect 106980 526058 107460 526120
rect 106980 526002 107006 526058
rect 107062 526002 107130 526058
rect 107186 526002 107254 526058
rect 107310 526002 107378 526058
rect 107434 526002 107460 526058
rect 106980 525940 107460 526002
rect 107476 526058 107956 526120
rect 107476 526002 107502 526058
rect 107558 526002 107626 526058
rect 107682 526002 107750 526058
rect 107806 526002 107874 526058
rect 107930 526002 107956 526058
rect 107476 525940 107956 526002
rect 107972 526058 108452 526120
rect 107972 526002 107998 526058
rect 108054 526002 108122 526058
rect 108178 526002 108246 526058
rect 108302 526002 108370 526058
rect 108426 526002 108452 526058
rect 107972 525940 108452 526002
rect 108468 526058 108948 526120
rect 108468 526002 108494 526058
rect 108550 526002 108618 526058
rect 108674 526002 108742 526058
rect 108798 526002 108866 526058
rect 108922 526002 108948 526058
rect 108468 525940 108948 526002
rect 108964 526058 109444 526120
rect 108964 526002 108990 526058
rect 109046 526002 109114 526058
rect 109170 526002 109238 526058
rect 109294 526002 109362 526058
rect 109418 526002 109444 526058
rect 108964 525940 109444 526002
rect 109460 526058 109940 526120
rect 109460 526002 109486 526058
rect 109542 526002 109610 526058
rect 109666 526002 109734 526058
rect 109790 526002 109858 526058
rect 109914 526002 109940 526058
rect 109460 525940 109940 526002
rect 109956 526058 110436 526120
rect 109956 526002 109982 526058
rect 110038 526002 110106 526058
rect 110162 526002 110230 526058
rect 110286 526002 110354 526058
rect 110410 526002 110436 526058
rect 109956 525940 110436 526002
rect 110452 526058 110932 526120
rect 110452 526002 110478 526058
rect 110534 526002 110602 526058
rect 110658 526002 110726 526058
rect 110782 526002 110850 526058
rect 110906 526002 110932 526058
rect 110452 525940 110932 526002
rect 110948 526058 111428 526120
rect 110948 526002 110974 526058
rect 111030 526002 111098 526058
rect 111154 526002 111222 526058
rect 111278 526002 111346 526058
rect 111402 526002 111428 526058
rect 110948 525940 111428 526002
rect 111444 526058 111924 526120
rect 111444 526002 111470 526058
rect 111526 526002 111594 526058
rect 111650 526002 111718 526058
rect 111774 526002 111842 526058
rect 111898 526002 111924 526058
rect 111444 525940 111924 526002
rect 111940 526058 112420 526120
rect 111940 526002 111966 526058
rect 112022 526002 112090 526058
rect 112146 526002 112214 526058
rect 112270 526002 112338 526058
rect 112394 526002 112420 526058
rect 111940 525940 112420 526002
rect 112436 526058 112916 526120
rect 112436 526002 112462 526058
rect 112518 526002 112586 526058
rect 112642 526002 112710 526058
rect 112766 526002 112834 526058
rect 112890 526002 112916 526058
rect 112436 525940 112916 526002
rect 112932 526058 113412 526120
rect 112932 526002 112958 526058
rect 113014 526002 113082 526058
rect 113138 526002 113206 526058
rect 113262 526002 113330 526058
rect 113386 526002 113412 526058
rect 112932 525940 113412 526002
rect 113428 526058 113908 526120
rect 113428 526002 113454 526058
rect 113510 526002 113578 526058
rect 113634 526002 113702 526058
rect 113758 526002 113826 526058
rect 113882 526002 113908 526058
rect 113428 525940 113908 526002
rect 113924 526058 114404 526120
rect 113924 526002 113950 526058
rect 114006 526002 114074 526058
rect 114130 526002 114198 526058
rect 114254 526002 114322 526058
rect 114378 526002 114404 526058
rect 113924 525940 114404 526002
rect 114420 526058 114900 526120
rect 114420 526002 114446 526058
rect 114502 526002 114570 526058
rect 114626 526002 114694 526058
rect 114750 526002 114818 526058
rect 114874 526002 114900 526058
rect 114420 525940 114900 526002
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 60180 514412 60528 514446
rect 60180 514356 60202 514412
rect 60258 514356 60326 514412
rect 60382 514356 60450 514412
rect 60506 514356 60528 514412
rect 60180 514288 60528 514356
rect 60180 514232 60202 514288
rect 60258 514232 60326 514288
rect 60382 514232 60450 514288
rect 60506 514232 60528 514288
rect 60180 514164 60528 514232
rect 60180 514108 60202 514164
rect 60258 514108 60326 514164
rect 60382 514108 60450 514164
rect 60506 514108 60528 514164
rect 60180 514040 60528 514108
rect 60180 513984 60202 514040
rect 60258 513984 60326 514040
rect 60382 513984 60450 514040
rect 60506 513984 60528 514040
rect 60180 513916 60528 513984
rect 60180 513860 60202 513916
rect 60258 513860 60326 513916
rect 60382 513860 60450 513916
rect 60506 513860 60528 513916
rect 60180 513826 60528 513860
rect 60552 514412 61024 514446
rect 60552 514356 60574 514412
rect 60630 514356 60698 514412
rect 60754 514356 60822 514412
rect 60878 514356 60946 514412
rect 61002 514356 61024 514412
rect 60552 514288 61024 514356
rect 60552 514232 60574 514288
rect 60630 514232 60698 514288
rect 60754 514232 60822 514288
rect 60878 514232 60946 514288
rect 61002 514232 61024 514288
rect 60552 514164 61024 514232
rect 60552 514108 60574 514164
rect 60630 514108 60698 514164
rect 60754 514108 60822 514164
rect 60878 514108 60946 514164
rect 61002 514108 61024 514164
rect 60552 514040 61024 514108
rect 60552 513984 60574 514040
rect 60630 513984 60698 514040
rect 60754 513984 60822 514040
rect 60878 513984 60946 514040
rect 61002 513984 61024 514040
rect 60552 513916 61024 513984
rect 60552 513860 60574 513916
rect 60630 513860 60698 513916
rect 60754 513860 60822 513916
rect 60878 513860 60946 513916
rect 61002 513860 61024 513916
rect 60552 513826 61024 513860
rect 61048 514412 61520 514446
rect 61048 514356 61070 514412
rect 61126 514356 61194 514412
rect 61250 514356 61318 514412
rect 61374 514356 61442 514412
rect 61498 514356 61520 514412
rect 61048 514288 61520 514356
rect 61048 514232 61070 514288
rect 61126 514232 61194 514288
rect 61250 514232 61318 514288
rect 61374 514232 61442 514288
rect 61498 514232 61520 514288
rect 61048 514164 61520 514232
rect 61048 514108 61070 514164
rect 61126 514108 61194 514164
rect 61250 514108 61318 514164
rect 61374 514108 61442 514164
rect 61498 514108 61520 514164
rect 61048 514040 61520 514108
rect 61048 513984 61070 514040
rect 61126 513984 61194 514040
rect 61250 513984 61318 514040
rect 61374 513984 61442 514040
rect 61498 513984 61520 514040
rect 61048 513916 61520 513984
rect 61048 513860 61070 513916
rect 61126 513860 61194 513916
rect 61250 513860 61318 513916
rect 61374 513860 61442 513916
rect 61498 513860 61520 513916
rect 61048 513826 61520 513860
rect 61544 514412 62016 514446
rect 61544 514356 61566 514412
rect 61622 514356 61690 514412
rect 61746 514356 61814 514412
rect 61870 514356 61938 514412
rect 61994 514356 62016 514412
rect 61544 514288 62016 514356
rect 61544 514232 61566 514288
rect 61622 514232 61690 514288
rect 61746 514232 61814 514288
rect 61870 514232 61938 514288
rect 61994 514232 62016 514288
rect 61544 514164 62016 514232
rect 61544 514108 61566 514164
rect 61622 514108 61690 514164
rect 61746 514108 61814 514164
rect 61870 514108 61938 514164
rect 61994 514108 62016 514164
rect 61544 514040 62016 514108
rect 61544 513984 61566 514040
rect 61622 513984 61690 514040
rect 61746 513984 61814 514040
rect 61870 513984 61938 514040
rect 61994 513984 62016 514040
rect 61544 513916 62016 513984
rect 61544 513860 61566 513916
rect 61622 513860 61690 513916
rect 61746 513860 61814 513916
rect 61870 513860 61938 513916
rect 61994 513860 62016 513916
rect 61544 513826 62016 513860
rect 62040 514412 62512 514446
rect 62040 514356 62062 514412
rect 62118 514356 62186 514412
rect 62242 514356 62310 514412
rect 62366 514356 62434 514412
rect 62490 514356 62512 514412
rect 62040 514288 62512 514356
rect 62040 514232 62062 514288
rect 62118 514232 62186 514288
rect 62242 514232 62310 514288
rect 62366 514232 62434 514288
rect 62490 514232 62512 514288
rect 62040 514164 62512 514232
rect 62040 514108 62062 514164
rect 62118 514108 62186 514164
rect 62242 514108 62310 514164
rect 62366 514108 62434 514164
rect 62490 514108 62512 514164
rect 62040 514040 62512 514108
rect 62040 513984 62062 514040
rect 62118 513984 62186 514040
rect 62242 513984 62310 514040
rect 62366 513984 62434 514040
rect 62490 513984 62512 514040
rect 62040 513916 62512 513984
rect 62040 513860 62062 513916
rect 62118 513860 62186 513916
rect 62242 513860 62310 513916
rect 62366 513860 62434 513916
rect 62490 513860 62512 513916
rect 62040 513826 62512 513860
rect 62536 514412 63008 514446
rect 62536 514356 62558 514412
rect 62614 514356 62682 514412
rect 62738 514356 62806 514412
rect 62862 514356 62930 514412
rect 62986 514356 63008 514412
rect 62536 514288 63008 514356
rect 62536 514232 62558 514288
rect 62614 514232 62682 514288
rect 62738 514232 62806 514288
rect 62862 514232 62930 514288
rect 62986 514232 63008 514288
rect 62536 514164 63008 514232
rect 62536 514108 62558 514164
rect 62614 514108 62682 514164
rect 62738 514108 62806 514164
rect 62862 514108 62930 514164
rect 62986 514108 63008 514164
rect 62536 514040 63008 514108
rect 62536 513984 62558 514040
rect 62614 513984 62682 514040
rect 62738 513984 62806 514040
rect 62862 513984 62930 514040
rect 62986 513984 63008 514040
rect 62536 513916 63008 513984
rect 62536 513860 62558 513916
rect 62614 513860 62682 513916
rect 62738 513860 62806 513916
rect 62862 513860 62930 513916
rect 62986 513860 63008 513916
rect 62536 513826 63008 513860
rect 63032 514412 63504 514446
rect 63032 514356 63054 514412
rect 63110 514356 63178 514412
rect 63234 514356 63302 514412
rect 63358 514356 63426 514412
rect 63482 514356 63504 514412
rect 63032 514288 63504 514356
rect 63032 514232 63054 514288
rect 63110 514232 63178 514288
rect 63234 514232 63302 514288
rect 63358 514232 63426 514288
rect 63482 514232 63504 514288
rect 63032 514164 63504 514232
rect 63032 514108 63054 514164
rect 63110 514108 63178 514164
rect 63234 514108 63302 514164
rect 63358 514108 63426 514164
rect 63482 514108 63504 514164
rect 63032 514040 63504 514108
rect 63032 513984 63054 514040
rect 63110 513984 63178 514040
rect 63234 513984 63302 514040
rect 63358 513984 63426 514040
rect 63482 513984 63504 514040
rect 63032 513916 63504 513984
rect 63032 513860 63054 513916
rect 63110 513860 63178 513916
rect 63234 513860 63302 513916
rect 63358 513860 63426 513916
rect 63482 513860 63504 513916
rect 63032 513826 63504 513860
rect 63528 514412 64000 514446
rect 63528 514356 63550 514412
rect 63606 514356 63674 514412
rect 63730 514356 63798 514412
rect 63854 514356 63922 514412
rect 63978 514356 64000 514412
rect 63528 514288 64000 514356
rect 63528 514232 63550 514288
rect 63606 514232 63674 514288
rect 63730 514232 63798 514288
rect 63854 514232 63922 514288
rect 63978 514232 64000 514288
rect 63528 514164 64000 514232
rect 63528 514108 63550 514164
rect 63606 514108 63674 514164
rect 63730 514108 63798 514164
rect 63854 514108 63922 514164
rect 63978 514108 64000 514164
rect 63528 514040 64000 514108
rect 63528 513984 63550 514040
rect 63606 513984 63674 514040
rect 63730 513984 63798 514040
rect 63854 513984 63922 514040
rect 63978 513984 64000 514040
rect 63528 513916 64000 513984
rect 63528 513860 63550 513916
rect 63606 513860 63674 513916
rect 63730 513860 63798 513916
rect 63854 513860 63922 513916
rect 63978 513860 64000 513916
rect 63528 513826 64000 513860
rect 64024 514412 64496 514446
rect 64024 514356 64046 514412
rect 64102 514356 64170 514412
rect 64226 514356 64294 514412
rect 64350 514356 64418 514412
rect 64474 514356 64496 514412
rect 64024 514288 64496 514356
rect 64024 514232 64046 514288
rect 64102 514232 64170 514288
rect 64226 514232 64294 514288
rect 64350 514232 64418 514288
rect 64474 514232 64496 514288
rect 64024 514164 64496 514232
rect 64024 514108 64046 514164
rect 64102 514108 64170 514164
rect 64226 514108 64294 514164
rect 64350 514108 64418 514164
rect 64474 514108 64496 514164
rect 64024 514040 64496 514108
rect 64024 513984 64046 514040
rect 64102 513984 64170 514040
rect 64226 513984 64294 514040
rect 64350 513984 64418 514040
rect 64474 513984 64496 514040
rect 64024 513916 64496 513984
rect 64024 513860 64046 513916
rect 64102 513860 64170 513916
rect 64226 513860 64294 513916
rect 64350 513860 64418 513916
rect 64474 513860 64496 513916
rect 64024 513826 64496 513860
rect 64520 514412 64992 514446
rect 64520 514356 64542 514412
rect 64598 514356 64666 514412
rect 64722 514356 64790 514412
rect 64846 514356 64914 514412
rect 64970 514356 64992 514412
rect 64520 514288 64992 514356
rect 64520 514232 64542 514288
rect 64598 514232 64666 514288
rect 64722 514232 64790 514288
rect 64846 514232 64914 514288
rect 64970 514232 64992 514288
rect 64520 514164 64992 514232
rect 64520 514108 64542 514164
rect 64598 514108 64666 514164
rect 64722 514108 64790 514164
rect 64846 514108 64914 514164
rect 64970 514108 64992 514164
rect 64520 514040 64992 514108
rect 64520 513984 64542 514040
rect 64598 513984 64666 514040
rect 64722 513984 64790 514040
rect 64846 513984 64914 514040
rect 64970 513984 64992 514040
rect 64520 513916 64992 513984
rect 64520 513860 64542 513916
rect 64598 513860 64666 513916
rect 64722 513860 64790 513916
rect 64846 513860 64914 513916
rect 64970 513860 64992 513916
rect 64520 513826 64992 513860
rect 65016 514412 65488 514446
rect 65016 514356 65038 514412
rect 65094 514356 65162 514412
rect 65218 514356 65286 514412
rect 65342 514356 65410 514412
rect 65466 514356 65488 514412
rect 65016 514288 65488 514356
rect 65016 514232 65038 514288
rect 65094 514232 65162 514288
rect 65218 514232 65286 514288
rect 65342 514232 65410 514288
rect 65466 514232 65488 514288
rect 65016 514164 65488 514232
rect 65016 514108 65038 514164
rect 65094 514108 65162 514164
rect 65218 514108 65286 514164
rect 65342 514108 65410 514164
rect 65466 514108 65488 514164
rect 65016 514040 65488 514108
rect 65016 513984 65038 514040
rect 65094 513984 65162 514040
rect 65218 513984 65286 514040
rect 65342 513984 65410 514040
rect 65466 513984 65488 514040
rect 65016 513916 65488 513984
rect 65016 513860 65038 513916
rect 65094 513860 65162 513916
rect 65218 513860 65286 513916
rect 65342 513860 65410 513916
rect 65466 513860 65488 513916
rect 65016 513826 65488 513860
rect 65512 514412 65984 514446
rect 65512 514356 65534 514412
rect 65590 514356 65658 514412
rect 65714 514356 65782 514412
rect 65838 514356 65906 514412
rect 65962 514356 65984 514412
rect 65512 514288 65984 514356
rect 65512 514232 65534 514288
rect 65590 514232 65658 514288
rect 65714 514232 65782 514288
rect 65838 514232 65906 514288
rect 65962 514232 65984 514288
rect 65512 514164 65984 514232
rect 65512 514108 65534 514164
rect 65590 514108 65658 514164
rect 65714 514108 65782 514164
rect 65838 514108 65906 514164
rect 65962 514108 65984 514164
rect 65512 514040 65984 514108
rect 65512 513984 65534 514040
rect 65590 513984 65658 514040
rect 65714 513984 65782 514040
rect 65838 513984 65906 514040
rect 65962 513984 65984 514040
rect 65512 513916 65984 513984
rect 65512 513860 65534 513916
rect 65590 513860 65658 513916
rect 65714 513860 65782 513916
rect 65838 513860 65906 513916
rect 65962 513860 65984 513916
rect 65512 513826 65984 513860
rect 66008 514412 66480 514446
rect 66008 514356 66030 514412
rect 66086 514356 66154 514412
rect 66210 514356 66278 514412
rect 66334 514356 66402 514412
rect 66458 514356 66480 514412
rect 66008 514288 66480 514356
rect 66008 514232 66030 514288
rect 66086 514232 66154 514288
rect 66210 514232 66278 514288
rect 66334 514232 66402 514288
rect 66458 514232 66480 514288
rect 66008 514164 66480 514232
rect 66008 514108 66030 514164
rect 66086 514108 66154 514164
rect 66210 514108 66278 514164
rect 66334 514108 66402 514164
rect 66458 514108 66480 514164
rect 66008 514040 66480 514108
rect 66008 513984 66030 514040
rect 66086 513984 66154 514040
rect 66210 513984 66278 514040
rect 66334 513984 66402 514040
rect 66458 513984 66480 514040
rect 66008 513916 66480 513984
rect 66008 513860 66030 513916
rect 66086 513860 66154 513916
rect 66210 513860 66278 513916
rect 66334 513860 66402 513916
rect 66458 513860 66480 513916
rect 66008 513826 66480 513860
rect 90060 508435 100140 508446
rect 90060 508379 90112 508435
rect 90168 508379 90236 508435
rect 90292 508379 90360 508435
rect 90416 508379 90484 508435
rect 90540 508379 90608 508435
rect 90664 508379 90732 508435
rect 90788 508379 90856 508435
rect 90912 508379 90980 508435
rect 91036 508379 91104 508435
rect 91160 508379 91228 508435
rect 91284 508379 91352 508435
rect 91408 508379 91476 508435
rect 91532 508379 91600 508435
rect 91656 508379 91724 508435
rect 91780 508379 91848 508435
rect 91904 508379 91972 508435
rect 92028 508379 92096 508435
rect 92152 508379 92220 508435
rect 92276 508379 92344 508435
rect 92400 508379 92468 508435
rect 92524 508379 92592 508435
rect 92648 508379 92716 508435
rect 92772 508379 92840 508435
rect 92896 508379 92964 508435
rect 93020 508379 93088 508435
rect 93144 508379 93212 508435
rect 93268 508379 93336 508435
rect 93392 508379 93460 508435
rect 93516 508379 93584 508435
rect 93640 508379 93708 508435
rect 93764 508379 93832 508435
rect 93888 508379 93956 508435
rect 94012 508379 94080 508435
rect 94136 508379 94204 508435
rect 94260 508379 94328 508435
rect 94384 508379 94452 508435
rect 94508 508379 94576 508435
rect 94632 508379 94700 508435
rect 94756 508379 94824 508435
rect 94880 508379 94948 508435
rect 95004 508379 95072 508435
rect 95128 508379 95196 508435
rect 95252 508379 95320 508435
rect 95376 508379 95444 508435
rect 95500 508379 95568 508435
rect 95624 508379 95692 508435
rect 95748 508379 95816 508435
rect 95872 508379 95940 508435
rect 95996 508379 96064 508435
rect 96120 508379 96188 508435
rect 96244 508379 96312 508435
rect 96368 508379 96436 508435
rect 96492 508379 96560 508435
rect 96616 508379 96684 508435
rect 96740 508379 96808 508435
rect 96864 508379 96932 508435
rect 96988 508379 97056 508435
rect 97112 508379 97180 508435
rect 97236 508379 97304 508435
rect 97360 508379 97428 508435
rect 97484 508379 97552 508435
rect 97608 508379 97676 508435
rect 97732 508379 97800 508435
rect 97856 508379 97924 508435
rect 97980 508379 98048 508435
rect 98104 508379 98172 508435
rect 98228 508379 98296 508435
rect 98352 508379 98420 508435
rect 98476 508379 98544 508435
rect 98600 508379 98668 508435
rect 98724 508379 98792 508435
rect 98848 508379 98916 508435
rect 98972 508379 99040 508435
rect 99096 508379 99164 508435
rect 99220 508379 99288 508435
rect 99344 508379 99412 508435
rect 99468 508379 99536 508435
rect 99592 508379 99660 508435
rect 99716 508379 99784 508435
rect 99840 508379 99908 508435
rect 99964 508379 100032 508435
rect 100088 508379 100140 508435
rect 90060 508311 100140 508379
rect 90060 508255 90112 508311
rect 90168 508255 90236 508311
rect 90292 508255 90360 508311
rect 90416 508255 90484 508311
rect 90540 508255 90608 508311
rect 90664 508255 90732 508311
rect 90788 508255 90856 508311
rect 90912 508255 90980 508311
rect 91036 508255 91104 508311
rect 91160 508255 91228 508311
rect 91284 508255 91352 508311
rect 91408 508255 91476 508311
rect 91532 508255 91600 508311
rect 91656 508255 91724 508311
rect 91780 508255 91848 508311
rect 91904 508255 91972 508311
rect 92028 508255 92096 508311
rect 92152 508255 92220 508311
rect 92276 508255 92344 508311
rect 92400 508255 92468 508311
rect 92524 508255 92592 508311
rect 92648 508255 92716 508311
rect 92772 508255 92840 508311
rect 92896 508255 92964 508311
rect 93020 508255 93088 508311
rect 93144 508255 93212 508311
rect 93268 508255 93336 508311
rect 93392 508255 93460 508311
rect 93516 508255 93584 508311
rect 93640 508255 93708 508311
rect 93764 508255 93832 508311
rect 93888 508255 93956 508311
rect 94012 508255 94080 508311
rect 94136 508255 94204 508311
rect 94260 508255 94328 508311
rect 94384 508255 94452 508311
rect 94508 508255 94576 508311
rect 94632 508255 94700 508311
rect 94756 508255 94824 508311
rect 94880 508255 94948 508311
rect 95004 508255 95072 508311
rect 95128 508255 95196 508311
rect 95252 508255 95320 508311
rect 95376 508255 95444 508311
rect 95500 508255 95568 508311
rect 95624 508255 95692 508311
rect 95748 508255 95816 508311
rect 95872 508255 95940 508311
rect 95996 508255 96064 508311
rect 96120 508255 96188 508311
rect 96244 508255 96312 508311
rect 96368 508255 96436 508311
rect 96492 508255 96560 508311
rect 96616 508255 96684 508311
rect 96740 508255 96808 508311
rect 96864 508255 96932 508311
rect 96988 508255 97056 508311
rect 97112 508255 97180 508311
rect 97236 508255 97304 508311
rect 97360 508255 97428 508311
rect 97484 508255 97552 508311
rect 97608 508255 97676 508311
rect 97732 508255 97800 508311
rect 97856 508255 97924 508311
rect 97980 508255 98048 508311
rect 98104 508255 98172 508311
rect 98228 508255 98296 508311
rect 98352 508255 98420 508311
rect 98476 508255 98544 508311
rect 98600 508255 98668 508311
rect 98724 508255 98792 508311
rect 98848 508255 98916 508311
rect 98972 508255 99040 508311
rect 99096 508255 99164 508311
rect 99220 508255 99288 508311
rect 99344 508255 99412 508311
rect 99468 508255 99536 508311
rect 99592 508255 99660 508311
rect 99716 508255 99784 508311
rect 99840 508255 99908 508311
rect 99964 508255 100032 508311
rect 100088 508255 100140 508311
rect 90060 508187 100140 508255
rect 90060 508131 90112 508187
rect 90168 508131 90236 508187
rect 90292 508131 90360 508187
rect 90416 508131 90484 508187
rect 90540 508131 90608 508187
rect 90664 508131 90732 508187
rect 90788 508131 90856 508187
rect 90912 508131 90980 508187
rect 91036 508131 91104 508187
rect 91160 508131 91228 508187
rect 91284 508131 91352 508187
rect 91408 508131 91476 508187
rect 91532 508131 91600 508187
rect 91656 508131 91724 508187
rect 91780 508131 91848 508187
rect 91904 508131 91972 508187
rect 92028 508131 92096 508187
rect 92152 508131 92220 508187
rect 92276 508131 92344 508187
rect 92400 508131 92468 508187
rect 92524 508131 92592 508187
rect 92648 508131 92716 508187
rect 92772 508131 92840 508187
rect 92896 508131 92964 508187
rect 93020 508131 93088 508187
rect 93144 508131 93212 508187
rect 93268 508131 93336 508187
rect 93392 508131 93460 508187
rect 93516 508131 93584 508187
rect 93640 508131 93708 508187
rect 93764 508131 93832 508187
rect 93888 508131 93956 508187
rect 94012 508131 94080 508187
rect 94136 508131 94204 508187
rect 94260 508131 94328 508187
rect 94384 508131 94452 508187
rect 94508 508131 94576 508187
rect 94632 508131 94700 508187
rect 94756 508131 94824 508187
rect 94880 508131 94948 508187
rect 95004 508131 95072 508187
rect 95128 508131 95196 508187
rect 95252 508131 95320 508187
rect 95376 508131 95444 508187
rect 95500 508131 95568 508187
rect 95624 508131 95692 508187
rect 95748 508131 95816 508187
rect 95872 508131 95940 508187
rect 95996 508131 96064 508187
rect 96120 508131 96188 508187
rect 96244 508131 96312 508187
rect 96368 508131 96436 508187
rect 96492 508131 96560 508187
rect 96616 508131 96684 508187
rect 96740 508131 96808 508187
rect 96864 508131 96932 508187
rect 96988 508131 97056 508187
rect 97112 508131 97180 508187
rect 97236 508131 97304 508187
rect 97360 508131 97428 508187
rect 97484 508131 97552 508187
rect 97608 508131 97676 508187
rect 97732 508131 97800 508187
rect 97856 508131 97924 508187
rect 97980 508131 98048 508187
rect 98104 508131 98172 508187
rect 98228 508131 98296 508187
rect 98352 508131 98420 508187
rect 98476 508131 98544 508187
rect 98600 508131 98668 508187
rect 98724 508131 98792 508187
rect 98848 508131 98916 508187
rect 98972 508131 99040 508187
rect 99096 508131 99164 508187
rect 99220 508131 99288 508187
rect 99344 508131 99412 508187
rect 99468 508131 99536 508187
rect 99592 508131 99660 508187
rect 99716 508131 99784 508187
rect 99840 508131 99908 508187
rect 99964 508131 100032 508187
rect 100088 508131 100140 508187
rect 90060 508120 100140 508131
rect 159018 508350 159638 525922
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 89880 507911 90356 507940
rect 89880 507855 89904 507911
rect 89960 507855 90028 507911
rect 90084 507855 90152 507911
rect 90208 507855 90276 507911
rect 90332 507855 90356 507911
rect 89880 507826 90356 507855
rect 90376 507911 90852 507940
rect 90376 507855 90400 507911
rect 90456 507855 90524 507911
rect 90580 507855 90648 507911
rect 90704 507855 90772 507911
rect 90828 507855 90852 507911
rect 90376 507826 90852 507855
rect 90872 507911 91348 507940
rect 90872 507855 90896 507911
rect 90952 507855 91020 507911
rect 91076 507855 91144 507911
rect 91200 507855 91268 507911
rect 91324 507855 91348 507911
rect 90872 507826 91348 507855
rect 91368 507911 91844 507940
rect 91368 507855 91392 507911
rect 91448 507855 91516 507911
rect 91572 507855 91640 507911
rect 91696 507855 91764 507911
rect 91820 507855 91844 507911
rect 91368 507826 91844 507855
rect 91864 507911 92340 507940
rect 91864 507855 91888 507911
rect 91944 507855 92012 507911
rect 92068 507855 92136 507911
rect 92192 507855 92260 507911
rect 92316 507855 92340 507911
rect 91864 507826 92340 507855
rect 92360 507911 92836 507940
rect 92360 507855 92384 507911
rect 92440 507855 92508 507911
rect 92564 507855 92632 507911
rect 92688 507855 92756 507911
rect 92812 507855 92836 507911
rect 92360 507826 92836 507855
rect 92856 507911 93332 507940
rect 92856 507855 92880 507911
rect 92936 507855 93004 507911
rect 93060 507855 93128 507911
rect 93184 507855 93252 507911
rect 93308 507855 93332 507911
rect 92856 507826 93332 507855
rect 93352 507911 93828 507940
rect 93352 507855 93376 507911
rect 93432 507855 93500 507911
rect 93556 507855 93624 507911
rect 93680 507855 93748 507911
rect 93804 507855 93828 507911
rect 93352 507826 93828 507855
rect 93848 507911 94324 507940
rect 93848 507855 93872 507911
rect 93928 507855 93996 507911
rect 94052 507855 94120 507911
rect 94176 507855 94244 507911
rect 94300 507855 94324 507911
rect 93848 507826 94324 507855
rect 94344 507911 94820 507940
rect 94344 507855 94368 507911
rect 94424 507855 94492 507911
rect 94548 507855 94616 507911
rect 94672 507855 94740 507911
rect 94796 507855 94820 507911
rect 94344 507826 94820 507855
rect 94840 507911 95316 507940
rect 94840 507855 94864 507911
rect 94920 507855 94988 507911
rect 95044 507855 95112 507911
rect 95168 507855 95236 507911
rect 95292 507855 95316 507911
rect 94840 507826 95316 507855
rect 95336 507911 95812 507940
rect 95336 507855 95360 507911
rect 95416 507855 95484 507911
rect 95540 507855 95608 507911
rect 95664 507855 95732 507911
rect 95788 507855 95812 507911
rect 95336 507826 95812 507855
rect 95832 507911 96308 507940
rect 95832 507855 95856 507911
rect 95912 507855 95980 507911
rect 96036 507855 96104 507911
rect 96160 507855 96228 507911
rect 96284 507855 96308 507911
rect 95832 507826 96308 507855
rect 96328 507911 96804 507940
rect 96328 507855 96352 507911
rect 96408 507855 96476 507911
rect 96532 507855 96600 507911
rect 96656 507855 96724 507911
rect 96780 507855 96804 507911
rect 96328 507826 96804 507855
rect 96824 507911 97300 507940
rect 96824 507855 96848 507911
rect 96904 507855 96972 507911
rect 97028 507855 97096 507911
rect 97152 507855 97220 507911
rect 97276 507855 97300 507911
rect 96824 507826 97300 507855
rect 97320 507911 97796 507940
rect 97320 507855 97344 507911
rect 97400 507855 97468 507911
rect 97524 507855 97592 507911
rect 97648 507855 97716 507911
rect 97772 507855 97796 507911
rect 97320 507826 97796 507855
rect 97816 507911 98292 507940
rect 97816 507855 97840 507911
rect 97896 507855 97964 507911
rect 98020 507855 98088 507911
rect 98144 507855 98212 507911
rect 98268 507855 98292 507911
rect 97816 507826 98292 507855
rect 98312 507911 98788 507940
rect 98312 507855 98336 507911
rect 98392 507855 98460 507911
rect 98516 507855 98584 507911
rect 98640 507855 98708 507911
rect 98764 507855 98788 507911
rect 98312 507826 98788 507855
rect 98808 507911 99284 507940
rect 98808 507855 98832 507911
rect 98888 507855 98956 507911
rect 99012 507855 99080 507911
rect 99136 507855 99204 507911
rect 99260 507855 99284 507911
rect 98808 507826 99284 507855
rect 99304 507911 99780 507940
rect 99304 507855 99328 507911
rect 99384 507855 99452 507911
rect 99508 507855 99576 507911
rect 99632 507855 99700 507911
rect 99756 507855 99780 507911
rect 99304 507826 99780 507855
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 63420 496212 63496 496240
rect 63420 496156 63430 496212
rect 63486 496156 63496 496212
rect 63420 496088 63496 496156
rect 63420 496032 63430 496088
rect 63486 496032 63496 496088
rect 63420 495964 63496 496032
rect 63420 495908 63430 495964
rect 63486 495908 63496 495964
rect 63420 495880 63496 495908
rect 63544 496212 63992 496240
rect 63544 496156 63554 496212
rect 63610 496156 63678 496212
rect 63734 496156 63802 496212
rect 63858 496156 63926 496212
rect 63982 496156 63992 496212
rect 63544 496088 63992 496156
rect 63544 496032 63554 496088
rect 63610 496032 63678 496088
rect 63734 496032 63802 496088
rect 63858 496032 63926 496088
rect 63982 496032 63992 496088
rect 63544 495964 63992 496032
rect 63544 495908 63554 495964
rect 63610 495908 63678 495964
rect 63734 495908 63802 495964
rect 63858 495908 63926 495964
rect 63982 495908 63992 495964
rect 63544 495880 63992 495908
rect 64040 496212 64488 496240
rect 64040 496156 64050 496212
rect 64106 496156 64174 496212
rect 64230 496156 64298 496212
rect 64354 496156 64422 496212
rect 64478 496156 64488 496212
rect 64040 496088 64488 496156
rect 64040 496032 64050 496088
rect 64106 496032 64174 496088
rect 64230 496032 64298 496088
rect 64354 496032 64422 496088
rect 64478 496032 64488 496088
rect 64040 495964 64488 496032
rect 64040 495908 64050 495964
rect 64106 495908 64174 495964
rect 64230 495908 64298 495964
rect 64354 495908 64422 495964
rect 64478 495908 64488 495964
rect 64040 495880 64488 495908
rect 64536 496212 64984 496240
rect 64536 496156 64546 496212
rect 64602 496156 64670 496212
rect 64726 496156 64794 496212
rect 64850 496156 64918 496212
rect 64974 496156 64984 496212
rect 64536 496088 64984 496156
rect 64536 496032 64546 496088
rect 64602 496032 64670 496088
rect 64726 496032 64794 496088
rect 64850 496032 64918 496088
rect 64974 496032 64984 496088
rect 64536 495964 64984 496032
rect 64536 495908 64546 495964
rect 64602 495908 64670 495964
rect 64726 495908 64794 495964
rect 64850 495908 64918 495964
rect 64974 495908 64984 495964
rect 64536 495880 64984 495908
rect 65032 496212 65480 496240
rect 65032 496156 65042 496212
rect 65098 496156 65166 496212
rect 65222 496156 65290 496212
rect 65346 496156 65414 496212
rect 65470 496156 65480 496212
rect 65032 496088 65480 496156
rect 65032 496032 65042 496088
rect 65098 496032 65166 496088
rect 65222 496032 65290 496088
rect 65346 496032 65414 496088
rect 65470 496032 65480 496088
rect 65032 495964 65480 496032
rect 65032 495908 65042 495964
rect 65098 495908 65166 495964
rect 65222 495908 65290 495964
rect 65346 495908 65414 495964
rect 65470 495908 65480 495964
rect 65032 495880 65480 495908
rect 65528 496212 65976 496240
rect 65528 496156 65538 496212
rect 65594 496156 65662 496212
rect 65718 496156 65786 496212
rect 65842 496156 65910 496212
rect 65966 496156 65976 496212
rect 65528 496088 65976 496156
rect 65528 496032 65538 496088
rect 65594 496032 65662 496088
rect 65718 496032 65786 496088
rect 65842 496032 65910 496088
rect 65966 496032 65976 496088
rect 65528 495964 65976 496032
rect 65528 495908 65538 495964
rect 65594 495908 65662 495964
rect 65718 495908 65786 495964
rect 65842 495908 65910 495964
rect 65966 495908 65976 495964
rect 65528 495880 65976 495908
rect 66024 496212 66472 496240
rect 66024 496156 66034 496212
rect 66090 496156 66158 496212
rect 66214 496156 66282 496212
rect 66338 496156 66406 496212
rect 66462 496156 66472 496212
rect 66024 496088 66472 496156
rect 66024 496032 66034 496088
rect 66090 496032 66158 496088
rect 66214 496032 66282 496088
rect 66338 496032 66406 496088
rect 66462 496032 66472 496088
rect 66024 495964 66472 496032
rect 66024 495908 66034 495964
rect 66090 495908 66158 495964
rect 66214 495908 66282 495964
rect 66338 495908 66406 495964
rect 66462 495908 66472 495964
rect 66024 495880 66472 495908
rect 66520 496212 66968 496240
rect 66520 496156 66530 496212
rect 66586 496156 66654 496212
rect 66710 496156 66778 496212
rect 66834 496156 66902 496212
rect 66958 496156 66968 496212
rect 66520 496088 66968 496156
rect 66520 496032 66530 496088
rect 66586 496032 66654 496088
rect 66710 496032 66778 496088
rect 66834 496032 66902 496088
rect 66958 496032 66968 496088
rect 66520 495964 66968 496032
rect 66520 495908 66530 495964
rect 66586 495908 66654 495964
rect 66710 495908 66778 495964
rect 66834 495908 66902 495964
rect 66958 495908 66968 495964
rect 66520 495880 66968 495908
rect 67016 496212 67464 496240
rect 67016 496156 67026 496212
rect 67082 496156 67150 496212
rect 67206 496156 67274 496212
rect 67330 496156 67398 496212
rect 67454 496156 67464 496212
rect 67016 496088 67464 496156
rect 67016 496032 67026 496088
rect 67082 496032 67150 496088
rect 67206 496032 67274 496088
rect 67330 496032 67398 496088
rect 67454 496032 67464 496088
rect 67016 495964 67464 496032
rect 67016 495908 67026 495964
rect 67082 495908 67150 495964
rect 67206 495908 67274 495964
rect 67330 495908 67398 495964
rect 67454 495908 67464 495964
rect 67016 495880 67464 495908
rect 67512 496212 67960 496240
rect 67512 496156 67522 496212
rect 67578 496156 67646 496212
rect 67702 496156 67770 496212
rect 67826 496156 67894 496212
rect 67950 496156 67960 496212
rect 67512 496088 67960 496156
rect 67512 496032 67522 496088
rect 67578 496032 67646 496088
rect 67702 496032 67770 496088
rect 67826 496032 67894 496088
rect 67950 496032 67960 496088
rect 67512 495964 67960 496032
rect 67512 495908 67522 495964
rect 67578 495908 67646 495964
rect 67702 495908 67770 495964
rect 67826 495908 67894 495964
rect 67950 495908 67960 495964
rect 67512 495880 67960 495908
rect 68008 496212 68456 496240
rect 68008 496156 68018 496212
rect 68074 496156 68142 496212
rect 68198 496156 68266 496212
rect 68322 496156 68390 496212
rect 68446 496156 68456 496212
rect 68008 496088 68456 496156
rect 68008 496032 68018 496088
rect 68074 496032 68142 496088
rect 68198 496032 68266 496088
rect 68322 496032 68390 496088
rect 68446 496032 68456 496088
rect 68008 495964 68456 496032
rect 68008 495908 68018 495964
rect 68074 495908 68142 495964
rect 68198 495908 68266 495964
rect 68322 495908 68390 495964
rect 68446 495908 68456 495964
rect 68008 495880 68456 495908
rect 68504 496212 68952 496240
rect 68504 496156 68514 496212
rect 68570 496156 68638 496212
rect 68694 496156 68762 496212
rect 68818 496156 68886 496212
rect 68942 496156 68952 496212
rect 68504 496088 68952 496156
rect 68504 496032 68514 496088
rect 68570 496032 68638 496088
rect 68694 496032 68762 496088
rect 68818 496032 68886 496088
rect 68942 496032 68952 496088
rect 68504 495964 68952 496032
rect 68504 495908 68514 495964
rect 68570 495908 68638 495964
rect 68694 495908 68762 495964
rect 68818 495908 68886 495964
rect 68942 495908 68952 495964
rect 68504 495880 68952 495908
rect 69000 496212 69448 496240
rect 69000 496156 69010 496212
rect 69066 496156 69134 496212
rect 69190 496156 69258 496212
rect 69314 496156 69382 496212
rect 69438 496156 69448 496212
rect 69000 496088 69448 496156
rect 69000 496032 69010 496088
rect 69066 496032 69134 496088
rect 69190 496032 69258 496088
rect 69314 496032 69382 496088
rect 69438 496032 69448 496088
rect 69000 495964 69448 496032
rect 69000 495908 69010 495964
rect 69066 495908 69134 495964
rect 69190 495908 69258 495964
rect 69314 495908 69382 495964
rect 69438 495908 69448 495964
rect 69000 495880 69448 495908
rect 69496 496212 69944 496240
rect 69496 496156 69506 496212
rect 69562 496156 69630 496212
rect 69686 496156 69754 496212
rect 69810 496156 69878 496212
rect 69934 496156 69944 496212
rect 69496 496088 69944 496156
rect 69496 496032 69506 496088
rect 69562 496032 69630 496088
rect 69686 496032 69754 496088
rect 69810 496032 69878 496088
rect 69934 496032 69944 496088
rect 69496 495964 69944 496032
rect 69496 495908 69506 495964
rect 69562 495908 69630 495964
rect 69686 495908 69754 495964
rect 69810 495908 69878 495964
rect 69934 495908 69944 495964
rect 69496 495880 69944 495908
rect 69992 496212 70440 496240
rect 69992 496156 70002 496212
rect 70058 496156 70126 496212
rect 70182 496156 70250 496212
rect 70306 496156 70374 496212
rect 70430 496156 70440 496212
rect 69992 496088 70440 496156
rect 69992 496032 70002 496088
rect 70058 496032 70126 496088
rect 70182 496032 70250 496088
rect 70306 496032 70374 496088
rect 70430 496032 70440 496088
rect 69992 495964 70440 496032
rect 69992 495908 70002 495964
rect 70058 495908 70126 495964
rect 70182 495908 70250 495964
rect 70306 495908 70374 495964
rect 70430 495908 70440 495964
rect 69992 495880 70440 495908
rect 85200 490272 88800 490300
rect 85200 490216 85236 490272
rect 85292 490216 85360 490272
rect 85416 490216 85484 490272
rect 85540 490216 85608 490272
rect 85664 490216 85732 490272
rect 85788 490216 85856 490272
rect 85912 490216 85980 490272
rect 86036 490216 86104 490272
rect 86160 490216 86228 490272
rect 86284 490216 86352 490272
rect 86408 490216 86476 490272
rect 86532 490216 86600 490272
rect 86656 490216 86724 490272
rect 86780 490216 86848 490272
rect 86904 490216 86972 490272
rect 87028 490216 87096 490272
rect 87152 490216 87220 490272
rect 87276 490216 87344 490272
rect 87400 490216 87468 490272
rect 87524 490216 87592 490272
rect 87648 490216 87716 490272
rect 87772 490216 87840 490272
rect 87896 490216 87964 490272
rect 88020 490216 88088 490272
rect 88144 490216 88212 490272
rect 88268 490216 88336 490272
rect 88392 490216 88460 490272
rect 88516 490216 88584 490272
rect 88640 490216 88708 490272
rect 88764 490216 88800 490272
rect 85200 490148 88800 490216
rect 85200 490092 85236 490148
rect 85292 490092 85360 490148
rect 85416 490092 85484 490148
rect 85540 490092 85608 490148
rect 85664 490092 85732 490148
rect 85788 490092 85856 490148
rect 85912 490092 85980 490148
rect 86036 490092 86104 490148
rect 86160 490092 86228 490148
rect 86284 490092 86352 490148
rect 86408 490092 86476 490148
rect 86532 490092 86600 490148
rect 86656 490092 86724 490148
rect 86780 490092 86848 490148
rect 86904 490092 86972 490148
rect 87028 490092 87096 490148
rect 87152 490092 87220 490148
rect 87276 490092 87344 490148
rect 87400 490092 87468 490148
rect 87524 490092 87592 490148
rect 87648 490092 87716 490148
rect 87772 490092 87840 490148
rect 87896 490092 87964 490148
rect 88020 490092 88088 490148
rect 88144 490092 88212 490148
rect 88268 490092 88336 490148
rect 88392 490092 88460 490148
rect 88516 490092 88584 490148
rect 88640 490092 88708 490148
rect 88764 490092 88800 490148
rect 85200 490024 88800 490092
rect 85200 489968 85236 490024
rect 85292 489968 85360 490024
rect 85416 489968 85484 490024
rect 85540 489968 85608 490024
rect 85664 489968 85732 490024
rect 85788 489968 85856 490024
rect 85912 489968 85980 490024
rect 86036 489968 86104 490024
rect 86160 489968 86228 490024
rect 86284 489968 86352 490024
rect 86408 489968 86476 490024
rect 86532 489968 86600 490024
rect 86656 489968 86724 490024
rect 86780 489968 86848 490024
rect 86904 489968 86972 490024
rect 87028 489968 87096 490024
rect 87152 489968 87220 490024
rect 87276 489968 87344 490024
rect 87400 489968 87468 490024
rect 87524 489968 87592 490024
rect 87648 489968 87716 490024
rect 87772 489968 87840 490024
rect 87896 489968 87964 490024
rect 88020 489968 88088 490024
rect 88144 489968 88212 490024
rect 88268 489968 88336 490024
rect 88392 489968 88460 490024
rect 88516 489968 88584 490024
rect 88640 489968 88708 490024
rect 88764 489968 88800 490024
rect 85200 489940 88800 489968
rect 66858 472350 67478 486928
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 66858 436350 67478 453922
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 66858 418350 67478 435922
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 57932 403972 57988 403982
rect 62076 413476 62132 413486
rect 62076 395578 62132 413420
rect 66858 412556 67478 417922
rect 70578 478350 71198 482968
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 70578 478226 71198 478294
rect 80880 478358 81420 478420
rect 80880 478302 80936 478358
rect 80992 478302 81060 478358
rect 81116 478302 81184 478358
rect 81240 478302 81308 478358
rect 81364 478302 81420 478358
rect 80880 478240 81420 478302
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 70578 460350 71198 477922
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 70578 424350 71198 441922
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 66504 406350 66824 406384
rect 66504 406294 66574 406350
rect 66630 406294 66698 406350
rect 66754 406294 66824 406350
rect 66504 406226 66824 406294
rect 66504 406170 66574 406226
rect 66630 406170 66698 406226
rect 66754 406170 66824 406226
rect 66504 406102 66824 406170
rect 66504 406046 66574 406102
rect 66630 406046 66698 406102
rect 66754 406046 66824 406102
rect 66504 405978 66824 406046
rect 66504 405922 66574 405978
rect 66630 405922 66698 405978
rect 66754 405922 66824 405978
rect 66504 405888 66824 405922
rect 70578 406350 71198 423922
rect 97578 472350 98198 472944
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 97578 454350 98198 471922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 97578 436350 98198 453922
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 97578 418350 98198 435922
rect 97578 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 98198 418350
rect 97578 418226 98198 418294
rect 97578 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 98198 418226
rect 97578 418102 98198 418170
rect 97578 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 98198 418102
rect 97578 417978 98198 418046
rect 97578 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 98198 417978
rect 83916 416818 83972 416828
rect 83916 409892 83972 416762
rect 83916 409826 83972 409836
rect 70578 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71198 406350
rect 70578 406226 71198 406294
rect 70578 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71198 406226
rect 70578 406102 71198 406170
rect 70578 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71198 406102
rect 70578 405978 71198 406046
rect 70578 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71198 405978
rect 70578 405142 71198 405922
rect 71824 406350 72144 406384
rect 71824 406294 71894 406350
rect 71950 406294 72018 406350
rect 72074 406294 72144 406350
rect 71824 406226 72144 406294
rect 71824 406170 71894 406226
rect 71950 406170 72018 406226
rect 72074 406170 72144 406226
rect 71824 406102 72144 406170
rect 71824 406046 71894 406102
rect 71950 406046 72018 406102
rect 72074 406046 72144 406102
rect 71824 405978 72144 406046
rect 71824 405922 71894 405978
rect 71950 405922 72018 405978
rect 72074 405922 72144 405978
rect 71824 405888 72144 405922
rect 77144 406350 77464 406384
rect 77144 406294 77214 406350
rect 77270 406294 77338 406350
rect 77394 406294 77464 406350
rect 77144 406226 77464 406294
rect 77144 406170 77214 406226
rect 77270 406170 77338 406226
rect 77394 406170 77464 406226
rect 77144 406102 77464 406170
rect 77144 406046 77214 406102
rect 77270 406046 77338 406102
rect 77394 406046 77464 406102
rect 77144 405978 77464 406046
rect 77144 405922 77214 405978
rect 77270 405922 77338 405978
rect 77394 405922 77464 405978
rect 77144 405888 77464 405922
rect 82464 406350 82784 406384
rect 82464 406294 82534 406350
rect 82590 406294 82658 406350
rect 82714 406294 82784 406350
rect 82464 406226 82784 406294
rect 82464 406170 82534 406226
rect 82590 406170 82658 406226
rect 82714 406170 82784 406226
rect 82464 406102 82784 406170
rect 82464 406046 82534 406102
rect 82590 406046 82658 406102
rect 82714 406046 82784 406102
rect 82464 405978 82784 406046
rect 82464 405922 82534 405978
rect 82590 405922 82658 405978
rect 82714 405922 82784 405978
rect 82464 405888 82784 405922
rect 63844 400350 64164 400384
rect 63844 400294 63914 400350
rect 63970 400294 64038 400350
rect 64094 400294 64164 400350
rect 63844 400226 64164 400294
rect 63844 400170 63914 400226
rect 63970 400170 64038 400226
rect 64094 400170 64164 400226
rect 63844 400102 64164 400170
rect 63844 400046 63914 400102
rect 63970 400046 64038 400102
rect 64094 400046 64164 400102
rect 63844 399978 64164 400046
rect 63844 399922 63914 399978
rect 63970 399922 64038 399978
rect 64094 399922 64164 399978
rect 63844 399888 64164 399922
rect 69164 400350 69484 400384
rect 69164 400294 69234 400350
rect 69290 400294 69358 400350
rect 69414 400294 69484 400350
rect 69164 400226 69484 400294
rect 69164 400170 69234 400226
rect 69290 400170 69358 400226
rect 69414 400170 69484 400226
rect 74484 400350 74804 400384
rect 74484 400294 74554 400350
rect 74610 400294 74678 400350
rect 74734 400294 74804 400350
rect 74484 400226 74804 400294
rect 74484 400170 74554 400226
rect 74610 400170 74678 400226
rect 74734 400170 74804 400226
rect 69164 400102 69484 400170
rect 69164 400046 69234 400102
rect 69290 400046 69358 400102
rect 69414 400046 69484 400102
rect 69164 399978 69484 400046
rect 69164 399922 69234 399978
rect 69290 399922 69358 399978
rect 69414 399922 69484 399978
rect 69164 399888 69484 399922
rect 62076 395512 62132 395522
rect 39858 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 40478 388350
rect 39858 388226 40478 388294
rect 39858 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 40478 388226
rect 39858 388102 40478 388170
rect 39858 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 40478 388102
rect 39858 387978 40478 388046
rect 39858 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 40478 387978
rect 39858 370350 40478 387922
rect 39858 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 40478 370350
rect 39858 370226 40478 370294
rect 39858 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 40478 370226
rect 39858 370102 40478 370170
rect 39858 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 40478 370102
rect 39858 369978 40478 370046
rect 39858 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 40478 369978
rect 39858 352350 40478 369922
rect 66858 382350 67478 390964
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 66858 364350 67478 381922
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 39858 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 40478 352350
rect 39858 352226 40478 352294
rect 39858 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 40478 352226
rect 39858 352102 40478 352170
rect 39858 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 40478 352102
rect 39858 351978 40478 352046
rect 39858 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 40478 351978
rect 39858 334350 40478 351922
rect 64808 352350 65128 352384
rect 64808 352294 64878 352350
rect 64934 352294 65002 352350
rect 65058 352294 65128 352350
rect 64808 352226 65128 352294
rect 64808 352170 64878 352226
rect 64934 352170 65002 352226
rect 65058 352170 65128 352226
rect 64808 352102 65128 352170
rect 64808 352046 64878 352102
rect 64934 352046 65002 352102
rect 65058 352046 65128 352102
rect 64808 351978 65128 352046
rect 64808 351922 64878 351978
rect 64934 351922 65002 351978
rect 65058 351922 65128 351978
rect 64808 351888 65128 351922
rect 66858 351422 67478 363922
rect 70578 388350 71198 400170
rect 74484 400102 74804 400170
rect 74484 400046 74554 400102
rect 74610 400046 74678 400102
rect 74734 400046 74804 400102
rect 74484 399978 74804 400046
rect 74484 399922 74554 399978
rect 74610 399922 74678 399978
rect 74734 399922 74804 399978
rect 74484 399888 74804 399922
rect 79804 400350 80124 400384
rect 79804 400294 79874 400350
rect 79930 400294 79998 400350
rect 80054 400294 80124 400350
rect 79804 400226 80124 400294
rect 79804 400170 79874 400226
rect 79930 400170 79998 400226
rect 80054 400170 80124 400226
rect 79804 400102 80124 400170
rect 79804 400046 79874 400102
rect 79930 400046 79998 400102
rect 80054 400046 80124 400102
rect 79804 399978 80124 400046
rect 79804 399922 79874 399978
rect 79930 399922 79998 399978
rect 80054 399922 80124 399978
rect 79804 399888 80124 399922
rect 97578 400350 98198 417922
rect 97578 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 98198 400350
rect 97578 400226 98198 400294
rect 97578 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 98198 400226
rect 97578 400102 98198 400170
rect 97578 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 98198 400102
rect 97578 399978 98198 400046
rect 97578 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 98198 399978
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 70578 370350 71198 387922
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 352350 71198 369922
rect 70578 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 71198 352350
rect 70578 352226 71198 352294
rect 70578 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 71198 352226
rect 70578 352102 71198 352170
rect 70578 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 71198 352102
rect 70578 351978 71198 352046
rect 70578 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 71198 351978
rect 70578 351422 71198 351922
rect 91532 386596 91588 386606
rect 49448 346350 49768 346384
rect 49448 346294 49518 346350
rect 49574 346294 49642 346350
rect 49698 346294 49768 346350
rect 49448 346226 49768 346294
rect 49448 346170 49518 346226
rect 49574 346170 49642 346226
rect 49698 346170 49768 346226
rect 49448 346102 49768 346170
rect 49448 346046 49518 346102
rect 49574 346046 49642 346102
rect 49698 346046 49768 346102
rect 49448 345978 49768 346046
rect 49448 345922 49518 345978
rect 49574 345922 49642 345978
rect 49698 345922 49768 345978
rect 49448 345888 49768 345922
rect 80168 346350 80488 346384
rect 80168 346294 80238 346350
rect 80294 346294 80362 346350
rect 80418 346294 80488 346350
rect 80168 346226 80488 346294
rect 80168 346170 80238 346226
rect 80294 346170 80362 346226
rect 80418 346170 80488 346226
rect 80168 346102 80488 346170
rect 80168 346046 80238 346102
rect 80294 346046 80362 346102
rect 80418 346046 80488 346102
rect 80168 345978 80488 346046
rect 80168 345922 80238 345978
rect 80294 345922 80362 345978
rect 80418 345922 80488 345978
rect 80168 345888 80488 345922
rect 39858 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 40478 334350
rect 39858 334226 40478 334294
rect 39858 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 40478 334226
rect 39858 334102 40478 334170
rect 39858 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 40478 334102
rect 39858 333978 40478 334046
rect 39858 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 40478 333978
rect 39858 316350 40478 333922
rect 64808 334350 65128 334384
rect 64808 334294 64878 334350
rect 64934 334294 65002 334350
rect 65058 334294 65128 334350
rect 64808 334226 65128 334294
rect 64808 334170 64878 334226
rect 64934 334170 65002 334226
rect 65058 334170 65128 334226
rect 64808 334102 65128 334170
rect 64808 334046 64878 334102
rect 64934 334046 65002 334102
rect 65058 334046 65128 334102
rect 64808 333978 65128 334046
rect 64808 333922 64878 333978
rect 64934 333922 65002 333978
rect 65058 333922 65128 333978
rect 64808 333888 65128 333922
rect 49448 328350 49768 328384
rect 49448 328294 49518 328350
rect 49574 328294 49642 328350
rect 49698 328294 49768 328350
rect 49448 328226 49768 328294
rect 49448 328170 49518 328226
rect 49574 328170 49642 328226
rect 49698 328170 49768 328226
rect 49448 328102 49768 328170
rect 49448 328046 49518 328102
rect 49574 328046 49642 328102
rect 49698 328046 49768 328102
rect 49448 327978 49768 328046
rect 49448 327922 49518 327978
rect 49574 327922 49642 327978
rect 49698 327922 49768 327978
rect 49448 327888 49768 327922
rect 66858 328350 67478 337490
rect 66858 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 67478 328350
rect 66858 328226 67478 328294
rect 66858 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 67478 328226
rect 66858 328102 67478 328170
rect 66858 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 67478 328102
rect 66858 327978 67478 328046
rect 66858 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 67478 327978
rect 39858 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 40478 316350
rect 39858 316226 40478 316294
rect 39858 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 40478 316226
rect 39858 316102 40478 316170
rect 39858 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 40478 316102
rect 39858 315978 40478 316046
rect 39858 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 40478 315978
rect 39858 298350 40478 315922
rect 39858 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 40478 298350
rect 39858 298226 40478 298294
rect 39858 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 40478 298226
rect 39858 298102 40478 298170
rect 39858 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 40478 298102
rect 39858 297978 40478 298046
rect 39858 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 40478 297978
rect 39858 280350 40478 297922
rect 66858 310350 67478 327922
rect 66858 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 67478 310350
rect 66858 310226 67478 310294
rect 66858 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 67478 310226
rect 66858 310102 67478 310170
rect 66858 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 67478 310102
rect 66858 309978 67478 310046
rect 66858 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 67478 309978
rect 66858 292350 67478 309922
rect 66858 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 67478 292350
rect 66858 292226 67478 292294
rect 66858 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 67478 292226
rect 66858 292102 67478 292170
rect 66858 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 67478 292102
rect 66858 291978 67478 292046
rect 66858 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 67478 291978
rect 66858 289526 67478 291922
rect 70578 334350 71198 337490
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 70578 316350 71198 333922
rect 80168 328350 80488 328384
rect 80168 328294 80238 328350
rect 80294 328294 80362 328350
rect 80418 328294 80488 328350
rect 80168 328226 80488 328294
rect 80168 328170 80238 328226
rect 80294 328170 80362 328226
rect 80418 328170 80488 328226
rect 80168 328102 80488 328170
rect 80168 328046 80238 328102
rect 80294 328046 80362 328102
rect 80418 328046 80488 328102
rect 80168 327978 80488 328046
rect 80168 327922 80238 327978
rect 80294 327922 80362 327978
rect 80418 327922 80488 327978
rect 80168 327888 80488 327922
rect 70578 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 71198 316350
rect 70578 316226 71198 316294
rect 70578 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 71198 316226
rect 70578 316102 71198 316170
rect 70578 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 71198 316102
rect 70578 315978 71198 316046
rect 70578 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 71198 315978
rect 70578 298350 71198 315922
rect 85596 305938 85652 305948
rect 70578 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 71198 298350
rect 70578 298226 71198 298294
rect 70578 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 71198 298226
rect 70578 298102 71198 298170
rect 70578 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 71198 298102
rect 70578 297978 71198 298046
rect 70578 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 71198 297978
rect 70578 289526 71198 297922
rect 72156 302518 72212 302528
rect 72156 293972 72212 302462
rect 72156 293906 72212 293916
rect 85596 293972 85652 305882
rect 85596 293906 85652 293916
rect 39858 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 40478 280350
rect 39858 280226 40478 280294
rect 39858 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 40478 280226
rect 39858 280102 40478 280170
rect 39858 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 40478 280102
rect 39858 279978 40478 280046
rect 39858 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 40478 279978
rect 39858 262350 40478 279922
rect 59808 280350 60128 280384
rect 59808 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 60128 280350
rect 59808 280226 60128 280294
rect 59808 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 60128 280226
rect 59808 280102 60128 280170
rect 59808 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 60128 280102
rect 59808 279978 60128 280046
rect 59808 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 60128 279978
rect 59808 279888 60128 279922
rect 44448 274350 44768 274384
rect 44448 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 44768 274350
rect 44448 274226 44768 274294
rect 44448 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 44768 274226
rect 44448 274102 44768 274170
rect 44448 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 44768 274102
rect 44448 273978 44768 274046
rect 44448 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 44768 273978
rect 44448 273888 44768 273922
rect 75168 274350 75488 274384
rect 75168 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 75488 274350
rect 75168 274226 75488 274294
rect 75168 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 75488 274226
rect 75168 274102 75488 274170
rect 75168 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 75488 274102
rect 75168 273978 75488 274046
rect 75168 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 75488 273978
rect 75168 273888 75488 273922
rect 39858 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 40478 262350
rect 39858 262226 40478 262294
rect 39858 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 40478 262226
rect 39858 262102 40478 262170
rect 39858 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 40478 262102
rect 39858 261978 40478 262046
rect 39858 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 40478 261978
rect 39858 244350 40478 261922
rect 59808 262350 60128 262384
rect 59808 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 60128 262350
rect 59808 262226 60128 262294
rect 59808 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 60128 262226
rect 59808 262102 60128 262170
rect 59808 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 60128 262102
rect 59808 261978 60128 262046
rect 59808 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 60128 261978
rect 59808 261888 60128 261922
rect 44448 256350 44768 256384
rect 44448 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 44768 256350
rect 44448 256226 44768 256294
rect 44448 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 44768 256226
rect 44448 256102 44768 256170
rect 44448 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 44768 256102
rect 44448 255978 44768 256046
rect 44448 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 44768 255978
rect 44448 255888 44768 255922
rect 75168 256350 75488 256384
rect 75168 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 75488 256350
rect 75168 256226 75488 256294
rect 75168 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 75488 256226
rect 75168 256102 75488 256170
rect 75168 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 75488 256102
rect 75168 255978 75488 256046
rect 75168 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 75488 255978
rect 75168 255888 75488 255922
rect 39858 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 40478 244350
rect 39858 244226 40478 244294
rect 39858 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 40478 244226
rect 39858 244102 40478 244170
rect 39858 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 40478 244102
rect 39858 243978 40478 244046
rect 39858 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 40478 243978
rect 39858 226350 40478 243922
rect 42812 247078 42868 247088
rect 42812 233492 42868 247022
rect 59808 244350 60128 244384
rect 59808 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 60128 244350
rect 59808 244226 60128 244294
rect 59808 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 60128 244226
rect 59808 244102 60128 244170
rect 59808 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 60128 244102
rect 59808 243978 60128 244046
rect 59808 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 60128 243978
rect 59808 243888 60128 243922
rect 42812 233426 42868 233436
rect 66858 238350 67478 241770
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 39858 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 40478 226350
rect 39858 226226 40478 226294
rect 39858 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 40478 226226
rect 39858 226102 40478 226170
rect 39858 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 40478 226102
rect 39858 225978 40478 226046
rect 39858 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 40478 225978
rect 39858 208350 40478 225922
rect 41916 224420 41972 224430
rect 39858 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 40478 208350
rect 39858 208226 40478 208294
rect 39858 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 40478 208226
rect 39858 208102 40478 208170
rect 39858 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 40478 208102
rect 39858 207978 40478 208046
rect 39858 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 40478 207978
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 36138 184350 36758 201922
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 36138 166350 36758 183922
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 36138 148350 36758 165922
rect 39452 205858 39508 205868
rect 39452 163828 39508 205802
rect 39452 163762 39508 163772
rect 39858 190350 40478 207922
rect 39858 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 40478 190350
rect 39858 190226 40478 190294
rect 39858 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 40478 190226
rect 39858 190102 40478 190170
rect 39858 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 40478 190102
rect 39858 189978 40478 190046
rect 39858 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 40478 189978
rect 39858 172350 40478 189922
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 36138 130350 36758 147922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 36138 112350 36758 129922
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 36138 94350 36758 111922
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 36138 58350 36758 75922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 36138 40350 36758 57922
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 36138 22350 36758 39922
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 36138 4350 36758 21922
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 154350 40478 171922
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 136350 40478 153922
rect 39858 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 40478 136350
rect 39858 136226 40478 136294
rect 39858 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 40478 136226
rect 39858 136102 40478 136170
rect 39858 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 40478 136102
rect 39858 135978 40478 136046
rect 39858 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 40478 135978
rect 39858 118350 40478 135922
rect 39858 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 40478 118350
rect 39858 118226 40478 118294
rect 39858 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 40478 118226
rect 39858 118102 40478 118170
rect 39858 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 40478 118102
rect 39858 117978 40478 118046
rect 39858 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 40478 117978
rect 39858 100350 40478 117922
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 64350 40478 81922
rect 39858 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 40478 64350
rect 39858 64226 40478 64294
rect 39858 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 40478 64226
rect 39858 64102 40478 64170
rect 39858 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 40478 64102
rect 39858 63978 40478 64046
rect 39858 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 40478 63978
rect 39858 46350 40478 63922
rect 39858 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 40478 46350
rect 39858 46226 40478 46294
rect 39858 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 40478 46226
rect 39858 46102 40478 46170
rect 39858 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 40478 46102
rect 39858 45978 40478 46046
rect 39858 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 40478 45978
rect 39858 28350 40478 45922
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 41804 210898 41860 210908
rect 41804 5012 41860 210842
rect 41804 4946 41860 4956
rect 41916 4452 41972 224364
rect 66858 220350 67478 237922
rect 68012 237748 68068 237758
rect 68012 237652 68068 237662
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 66858 205590 67478 219922
rect 70578 226350 71198 241770
rect 71596 237636 71652 237646
rect 71596 237538 71652 237580
rect 71596 237472 71652 237482
rect 91532 237538 91588 386540
rect 91756 385028 91812 385038
rect 91756 237718 91812 384972
rect 97578 382350 98198 399922
rect 97578 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 98198 382350
rect 97578 382226 98198 382294
rect 97578 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 98198 382226
rect 97578 382102 98198 382170
rect 97578 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 98198 382102
rect 97578 381978 98198 382046
rect 97578 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 98198 381978
rect 97578 364350 98198 381922
rect 97578 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 98198 364350
rect 97578 364226 98198 364294
rect 97578 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 98198 364226
rect 97578 364102 98198 364170
rect 97578 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 98198 364102
rect 97578 363978 98198 364046
rect 97578 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 98198 363978
rect 97578 346350 98198 363922
rect 97578 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 98198 346350
rect 97578 346226 98198 346294
rect 97578 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 98198 346226
rect 97578 346102 98198 346170
rect 97578 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 98198 346102
rect 97578 345978 98198 346046
rect 97578 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 98198 345978
rect 97578 328350 98198 345922
rect 97578 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 98198 328350
rect 97578 328226 98198 328294
rect 97578 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 98198 328226
rect 97578 328102 98198 328170
rect 97578 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 98198 328102
rect 97578 327978 98198 328046
rect 97578 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 98198 327978
rect 97578 310350 98198 327922
rect 97578 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 98198 310350
rect 97578 310226 98198 310294
rect 97578 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 98198 310226
rect 97578 310102 98198 310170
rect 97578 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 98198 310102
rect 97578 309978 98198 310046
rect 97578 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 98198 309978
rect 97578 292350 98198 309922
rect 97578 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 98198 292350
rect 97578 292226 98198 292294
rect 97578 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 98198 292226
rect 97578 292102 98198 292170
rect 97578 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 98198 292102
rect 97578 291978 98198 292046
rect 97578 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 98198 291978
rect 96012 289268 96068 289278
rect 96012 285796 96068 289212
rect 96012 285730 96068 285740
rect 93660 285684 93716 285694
rect 93660 280420 93716 285628
rect 93660 280354 93716 280364
rect 93996 276164 94052 276174
rect 93996 275698 94052 276108
rect 93996 275632 94052 275642
rect 97578 274350 98198 291922
rect 97578 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 98198 274350
rect 97578 274226 98198 274294
rect 97578 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 98198 274226
rect 97578 274102 98198 274170
rect 97578 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 98198 274102
rect 97578 273978 98198 274046
rect 97578 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 98198 273978
rect 93436 271908 93492 271918
rect 93436 270658 93492 271852
rect 93436 270592 93492 270602
rect 91756 237652 91812 237662
rect 97578 256350 98198 273922
rect 97578 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 98198 256350
rect 97578 256226 98198 256294
rect 97578 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 98198 256226
rect 97578 256102 98198 256170
rect 97578 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 98198 256102
rect 97578 255978 98198 256046
rect 97578 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 98198 255978
rect 97578 238350 98198 255922
rect 97578 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 98198 238350
rect 97578 238226 98198 238294
rect 97578 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 98198 238226
rect 97578 238102 98198 238170
rect 97578 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 98198 238102
rect 97578 237978 98198 238046
rect 97578 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 98198 237978
rect 91532 237472 91588 237482
rect 70578 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 71198 226350
rect 70578 226226 71198 226294
rect 70578 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 71198 226226
rect 70578 226102 71198 226170
rect 70578 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 71198 226102
rect 70578 225978 71198 226046
rect 70578 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 71198 225978
rect 70578 208350 71198 225922
rect 70578 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 71198 208350
rect 70578 208226 71198 208294
rect 70578 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 71198 208226
rect 70578 208102 71198 208170
rect 70578 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 71198 208102
rect 70578 207978 71198 208046
rect 70578 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 71198 207978
rect 70578 205590 71198 207922
rect 97578 220350 98198 237922
rect 97578 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 98198 220350
rect 97578 220226 98198 220294
rect 97578 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 98198 220226
rect 97578 220102 98198 220170
rect 97578 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 98198 220102
rect 97578 219978 98198 220046
rect 97578 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 98198 219978
rect 97578 205590 98198 219922
rect 101298 460350 101918 473124
rect 101298 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 101918 460350
rect 101298 460226 101918 460294
rect 101298 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 101918 460226
rect 101298 460102 101918 460170
rect 101298 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 101918 460102
rect 101298 459978 101918 460046
rect 101298 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 101918 459978
rect 101298 442350 101918 459922
rect 101298 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 101918 442350
rect 101298 442226 101918 442294
rect 101298 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 101918 442226
rect 101298 442102 101918 442170
rect 101298 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 101918 442102
rect 101298 441978 101918 442046
rect 101298 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 101918 441978
rect 101298 424350 101918 441922
rect 101298 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 101918 424350
rect 101298 424226 101918 424294
rect 101298 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 101918 424226
rect 101298 424102 101918 424170
rect 101298 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 101918 424102
rect 101298 423978 101918 424046
rect 101298 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 101918 423978
rect 101298 406350 101918 423922
rect 101298 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 101918 406350
rect 101298 406226 101918 406294
rect 101298 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 101918 406226
rect 101298 406102 101918 406170
rect 101298 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 101918 406102
rect 101298 405978 101918 406046
rect 101298 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 101918 405978
rect 101298 388350 101918 405922
rect 101298 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 101918 388350
rect 101298 388226 101918 388294
rect 101298 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 101918 388226
rect 101298 388102 101918 388170
rect 101298 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 101918 388102
rect 101298 387978 101918 388046
rect 101298 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 101918 387978
rect 101298 370350 101918 387922
rect 128298 472350 128918 488604
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 128298 418350 128918 435922
rect 128298 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 128918 418350
rect 128298 418226 128918 418294
rect 128298 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 128918 418226
rect 128298 418102 128918 418170
rect 128298 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 128918 418102
rect 128298 417978 128918 418046
rect 128298 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 128918 417978
rect 128298 400350 128918 417922
rect 128298 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 128918 400350
rect 128298 400226 128918 400294
rect 128298 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 128918 400226
rect 128298 400102 128918 400170
rect 128298 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 128918 400102
rect 128298 399978 128918 400046
rect 128298 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 128918 399978
rect 128298 382350 128918 399922
rect 128298 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 128918 382350
rect 128298 382226 128918 382294
rect 128298 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 128918 382226
rect 128298 382102 128918 382170
rect 128298 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 128918 382102
rect 128298 381978 128918 382046
rect 128298 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 128918 381978
rect 101298 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 101918 370350
rect 101298 370226 101918 370294
rect 101298 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 101918 370226
rect 101298 370102 101918 370170
rect 101298 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 101918 370102
rect 101298 369978 101918 370046
rect 101298 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 101918 369978
rect 101298 352350 101918 369922
rect 101298 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 101918 352350
rect 101298 352226 101918 352294
rect 101298 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 101918 352226
rect 101298 352102 101918 352170
rect 101298 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 101918 352102
rect 101298 351978 101918 352046
rect 101298 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 101918 351978
rect 101298 334350 101918 351922
rect 101298 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 101918 334350
rect 101298 334226 101918 334294
rect 101298 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 101918 334226
rect 101298 334102 101918 334170
rect 101298 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 101918 334102
rect 101298 333978 101918 334046
rect 101298 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 101918 333978
rect 101298 316350 101918 333922
rect 101298 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 101918 316350
rect 101298 316226 101918 316294
rect 101298 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 101918 316226
rect 101298 316102 101918 316170
rect 101298 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 101918 316102
rect 101298 315978 101918 316046
rect 101298 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 101918 315978
rect 101298 298350 101918 315922
rect 101298 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 101918 298350
rect 101298 298226 101918 298294
rect 101298 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 101918 298226
rect 101298 298102 101918 298170
rect 101298 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 101918 298102
rect 101298 297978 101918 298046
rect 101298 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 101918 297978
rect 101298 280350 101918 297922
rect 108332 376498 108388 376508
rect 108332 293188 108388 376442
rect 128298 364350 128918 381922
rect 128298 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 128918 364350
rect 128298 364226 128918 364294
rect 128298 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 128918 364226
rect 128298 364102 128918 364170
rect 128298 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 128918 364102
rect 128298 363978 128918 364046
rect 128298 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 128918 363978
rect 119448 346350 119768 346384
rect 119448 346294 119518 346350
rect 119574 346294 119642 346350
rect 119698 346294 119768 346350
rect 119448 346226 119768 346294
rect 119448 346170 119518 346226
rect 119574 346170 119642 346226
rect 119698 346170 119768 346226
rect 119448 346102 119768 346170
rect 119448 346046 119518 346102
rect 119574 346046 119642 346102
rect 119698 346046 119768 346102
rect 119448 345978 119768 346046
rect 119448 345922 119518 345978
rect 119574 345922 119642 345978
rect 119698 345922 119768 345978
rect 119448 345888 119768 345922
rect 128298 346350 128918 363922
rect 132018 478350 132638 490764
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 132018 442350 132638 459922
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 424350 132638 441922
rect 132018 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 132638 424350
rect 132018 424226 132638 424294
rect 132018 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 132638 424226
rect 132018 424102 132638 424170
rect 132018 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 132638 424102
rect 132018 423978 132638 424046
rect 132018 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 132638 423978
rect 132018 406350 132638 423922
rect 132018 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 132638 406350
rect 132018 406226 132638 406294
rect 132018 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 132638 406226
rect 132018 406102 132638 406170
rect 132018 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 132638 406102
rect 132018 405978 132638 406046
rect 132018 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 132638 405978
rect 132018 388350 132638 405922
rect 132018 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 132638 388350
rect 132018 388226 132638 388294
rect 132018 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 132638 388226
rect 132018 388102 132638 388170
rect 132018 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 132638 388102
rect 132018 387978 132638 388046
rect 132018 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 132638 387978
rect 132018 370350 132638 387922
rect 132018 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 132638 370350
rect 132018 370226 132638 370294
rect 132018 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 132638 370226
rect 132018 370102 132638 370170
rect 132018 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 132638 370102
rect 132018 369978 132638 370046
rect 132018 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 132638 369978
rect 132018 359670 132638 369922
rect 159018 490350 159638 507922
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 159018 454350 159638 471922
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 159018 418350 159638 435922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 188972 590212 189028 590222
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 550350 163358 567922
rect 162738 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 163358 550350
rect 162738 550226 163358 550294
rect 162738 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 163358 550226
rect 162738 550102 163358 550170
rect 162738 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 163358 550102
rect 162738 549978 163358 550046
rect 162738 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 163358 549978
rect 162738 532350 163358 549922
rect 162738 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163358 532350
rect 162738 532226 163358 532294
rect 162738 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163358 532226
rect 162738 532102 163358 532170
rect 162738 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163358 532102
rect 162738 531978 163358 532046
rect 162738 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163358 531978
rect 162738 514350 163358 531922
rect 162738 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 163358 514350
rect 162738 514226 163358 514294
rect 162738 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 163358 514226
rect 162738 514102 163358 514170
rect 162738 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 163358 514102
rect 162738 513978 163358 514046
rect 162738 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 163358 513978
rect 162738 496350 163358 513922
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 162738 460350 163358 477922
rect 174636 573778 174692 573788
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 162738 442350 163358 459922
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 159018 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 159638 418350
rect 159018 418226 159638 418294
rect 159018 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 159638 418226
rect 159018 418102 159638 418170
rect 159018 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 159638 418102
rect 159018 417978 159638 418046
rect 159018 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 159638 417978
rect 159018 400350 159638 417922
rect 159018 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 159638 400350
rect 159018 400226 159638 400294
rect 159018 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 159638 400226
rect 159018 400102 159638 400170
rect 159018 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 159638 400102
rect 159018 399978 159638 400046
rect 159018 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 159638 399978
rect 159018 382350 159638 399922
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 159018 364350 159638 381922
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 159018 359670 159638 363922
rect 162092 431956 162148 431966
rect 134808 352350 135128 352384
rect 134808 352294 134878 352350
rect 134934 352294 135002 352350
rect 135058 352294 135128 352350
rect 134808 352226 135128 352294
rect 134808 352170 134878 352226
rect 134934 352170 135002 352226
rect 135058 352170 135128 352226
rect 134808 352102 135128 352170
rect 134808 352046 134878 352102
rect 134934 352046 135002 352102
rect 135058 352046 135128 352102
rect 134808 351978 135128 352046
rect 134808 351922 134878 351978
rect 134934 351922 135002 351978
rect 135058 351922 135128 351978
rect 134808 351888 135128 351922
rect 128298 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 128918 346350
rect 128298 346226 128918 346294
rect 128298 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 128918 346226
rect 128298 346102 128918 346170
rect 128298 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 128918 346102
rect 128298 345978 128918 346046
rect 128298 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 128918 345978
rect 119448 328350 119768 328384
rect 119448 328294 119518 328350
rect 119574 328294 119642 328350
rect 119698 328294 119768 328350
rect 119448 328226 119768 328294
rect 119448 328170 119518 328226
rect 119574 328170 119642 328226
rect 119698 328170 119768 328226
rect 119448 328102 119768 328170
rect 119448 328046 119518 328102
rect 119574 328046 119642 328102
rect 119698 328046 119768 328102
rect 119448 327978 119768 328046
rect 119448 327922 119518 327978
rect 119574 327922 119642 327978
rect 119698 327922 119768 327978
rect 119448 327888 119768 327922
rect 128298 328350 128918 345922
rect 150168 346350 150488 346384
rect 150168 346294 150238 346350
rect 150294 346294 150362 346350
rect 150418 346294 150488 346350
rect 150168 346226 150488 346294
rect 150168 346170 150238 346226
rect 150294 346170 150362 346226
rect 150418 346170 150488 346226
rect 150168 346102 150488 346170
rect 150168 346046 150238 346102
rect 150294 346046 150362 346102
rect 150418 346046 150488 346102
rect 150168 345978 150488 346046
rect 150168 345922 150238 345978
rect 150294 345922 150362 345978
rect 150418 345922 150488 345978
rect 150168 345888 150488 345922
rect 134808 334350 135128 334384
rect 134808 334294 134878 334350
rect 134934 334294 135002 334350
rect 135058 334294 135128 334350
rect 134808 334226 135128 334294
rect 134808 334170 134878 334226
rect 134934 334170 135002 334226
rect 135058 334170 135128 334226
rect 134808 334102 135128 334170
rect 134808 334046 134878 334102
rect 134934 334046 135002 334102
rect 135058 334046 135128 334102
rect 134808 333978 135128 334046
rect 134808 333922 134878 333978
rect 134934 333922 135002 333978
rect 135058 333922 135128 333978
rect 134808 333888 135128 333922
rect 128298 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 128918 328350
rect 128298 328226 128918 328294
rect 128298 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 128918 328226
rect 128298 328102 128918 328170
rect 128298 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 128918 328102
rect 128298 327978 128918 328046
rect 128298 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 128918 327978
rect 108332 293122 108388 293132
rect 128298 310350 128918 327922
rect 150168 328350 150488 328384
rect 150168 328294 150238 328350
rect 150294 328294 150362 328350
rect 150418 328294 150488 328350
rect 150168 328226 150488 328294
rect 150168 328170 150238 328226
rect 150294 328170 150362 328226
rect 150418 328170 150488 328226
rect 150168 328102 150488 328170
rect 150168 328046 150238 328102
rect 150294 328046 150362 328102
rect 150418 328046 150488 328102
rect 150168 327978 150488 328046
rect 150168 327922 150238 327978
rect 150294 327922 150362 327978
rect 150418 327922 150488 327978
rect 150168 327888 150488 327922
rect 128298 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 128918 310350
rect 128298 310226 128918 310294
rect 128298 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 128918 310226
rect 128298 310102 128918 310170
rect 128298 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 128918 310102
rect 128298 309978 128918 310046
rect 128298 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 128918 309978
rect 128298 292350 128918 309922
rect 128298 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 128918 292350
rect 128298 292226 128918 292294
rect 128298 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 128918 292226
rect 128298 292102 128918 292170
rect 128298 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 128918 292102
rect 128298 291978 128918 292046
rect 128298 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 128918 291978
rect 123452 288036 123508 288046
rect 101298 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 101918 280350
rect 101298 280226 101918 280294
rect 101298 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 101918 280226
rect 101298 280102 101918 280170
rect 101298 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 101918 280102
rect 101298 279978 101918 280046
rect 101298 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 101918 279978
rect 101298 262350 101918 279922
rect 101298 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 101918 262350
rect 101298 262226 101918 262294
rect 101298 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 101918 262226
rect 101298 262102 101918 262170
rect 101298 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 101918 262102
rect 101298 261978 101918 262046
rect 101298 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 101918 261978
rect 101298 244350 101918 261922
rect 101298 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 101918 244350
rect 101298 244226 101918 244294
rect 101298 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 101918 244226
rect 101298 244102 101918 244170
rect 101298 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 101918 244102
rect 101298 243978 101918 244046
rect 101298 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 101918 243978
rect 101298 226350 101918 243922
rect 101298 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 101918 226350
rect 101298 226226 101918 226294
rect 101298 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 101918 226226
rect 101298 226102 101918 226170
rect 101298 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 101918 226102
rect 101298 225978 101918 226046
rect 101298 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 101918 225978
rect 101298 208350 101918 225922
rect 108332 286916 108388 286926
rect 108332 220276 108388 286860
rect 108332 220210 108388 220220
rect 123452 210868 123508 287980
rect 123452 210802 123508 210812
rect 128298 274350 128918 291922
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 128298 256350 128918 273922
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 128298 238350 128918 255922
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 128298 220350 128918 237922
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 101298 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 101918 208350
rect 101298 208226 101918 208294
rect 101298 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 101918 208226
rect 101298 208102 101918 208170
rect 101298 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 101918 208102
rect 101298 207978 101918 208046
rect 101298 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 101918 207978
rect 101298 205590 101918 207922
rect 128298 205590 128918 219922
rect 132018 316350 132638 322218
rect 132018 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 132638 316350
rect 132018 316226 132638 316294
rect 132018 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 132638 316226
rect 132018 316102 132638 316170
rect 132018 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 132638 316102
rect 132018 315978 132638 316046
rect 132018 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 132638 315978
rect 132018 298350 132638 315922
rect 159018 310350 159638 322218
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 132018 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 132638 298350
rect 132018 298226 132638 298294
rect 132018 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 132638 298226
rect 132018 298102 132638 298170
rect 132018 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 132638 298102
rect 132018 297978 132638 298046
rect 132018 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 132638 297978
rect 132018 280350 132638 297922
rect 155372 304948 155428 304958
rect 137788 292404 137844 292414
rect 137788 290638 137844 292348
rect 137788 290572 137844 290582
rect 139244 290638 139300 290648
rect 139244 289044 139300 290582
rect 139244 288978 139300 288988
rect 155372 285348 155428 304892
rect 155372 285282 155428 285292
rect 159018 292350 159638 309922
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 159018 284908 159638 291922
rect 160412 313348 160468 313358
rect 160412 283556 160468 313292
rect 160412 283490 160468 283500
rect 161868 284676 161924 284686
rect 161868 280532 161924 284620
rect 162092 281316 162148 431900
rect 162738 424350 163358 441922
rect 162738 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 163358 424350
rect 162738 424226 163358 424294
rect 162738 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 163358 424226
rect 162738 424102 163358 424170
rect 162738 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 163358 424102
rect 162738 423978 163358 424046
rect 162738 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 163358 423978
rect 162738 406350 163358 423922
rect 162738 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163358 406350
rect 162738 406226 163358 406294
rect 162738 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163358 406226
rect 162738 406102 163358 406170
rect 162738 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163358 406102
rect 162738 405978 163358 406046
rect 162738 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163358 405978
rect 162738 388350 163358 405922
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 167132 469588 167188 469598
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162738 352350 163358 369922
rect 162738 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163358 352350
rect 162738 352226 163358 352294
rect 162738 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163358 352226
rect 162738 352102 163358 352170
rect 162738 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163358 352102
rect 162738 351978 163358 352046
rect 162738 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163358 351978
rect 162738 334350 163358 351922
rect 165452 377188 165508 377198
rect 162738 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 163358 334350
rect 162738 334226 163358 334294
rect 162738 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 163358 334226
rect 162738 334102 163358 334170
rect 162738 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 163358 334102
rect 162738 333978 163358 334046
rect 162738 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 163358 333978
rect 162738 316350 163358 333922
rect 163772 338548 163828 338558
rect 163772 326116 163828 338492
rect 163772 326050 163828 326060
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 162738 298350 163358 315922
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 162540 288932 162596 288942
rect 162540 282212 162596 288876
rect 162540 282146 162596 282156
rect 162092 281250 162148 281260
rect 161868 280466 161924 280476
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 132018 262350 132638 279922
rect 142008 280350 142328 280384
rect 142008 280294 142078 280350
rect 142134 280294 142202 280350
rect 142258 280294 142328 280350
rect 142008 280226 142328 280294
rect 142008 280170 142078 280226
rect 142134 280170 142202 280226
rect 142258 280170 142328 280226
rect 142008 280102 142328 280170
rect 142008 280046 142078 280102
rect 142134 280046 142202 280102
rect 142258 280046 142328 280102
rect 142008 279978 142328 280046
rect 142008 279922 142078 279978
rect 142134 279922 142202 279978
rect 142258 279922 142328 279978
rect 142008 279888 142328 279922
rect 147832 280350 148152 280384
rect 147832 280294 147902 280350
rect 147958 280294 148026 280350
rect 148082 280294 148152 280350
rect 147832 280226 148152 280294
rect 147832 280170 147902 280226
rect 147958 280170 148026 280226
rect 148082 280170 148152 280226
rect 147832 280102 148152 280170
rect 147832 280046 147902 280102
rect 147958 280046 148026 280102
rect 148082 280046 148152 280102
rect 147832 279978 148152 280046
rect 147832 279922 147902 279978
rect 147958 279922 148026 279978
rect 148082 279922 148152 279978
rect 147832 279888 148152 279922
rect 153656 280350 153976 280384
rect 153656 280294 153726 280350
rect 153782 280294 153850 280350
rect 153906 280294 153976 280350
rect 153656 280226 153976 280294
rect 153656 280170 153726 280226
rect 153782 280170 153850 280226
rect 153906 280170 153976 280226
rect 153656 280102 153976 280170
rect 153656 280046 153726 280102
rect 153782 280046 153850 280102
rect 153906 280046 153976 280102
rect 153656 279978 153976 280046
rect 153656 279922 153726 279978
rect 153782 279922 153850 279978
rect 153906 279922 153976 279978
rect 153656 279888 153976 279922
rect 159480 280350 159800 280384
rect 159480 280294 159550 280350
rect 159606 280294 159674 280350
rect 159730 280294 159800 280350
rect 159480 280226 159800 280294
rect 159480 280170 159550 280226
rect 159606 280170 159674 280226
rect 159730 280170 159800 280226
rect 159480 280102 159800 280170
rect 159480 280046 159550 280102
rect 159606 280046 159674 280102
rect 159730 280046 159800 280102
rect 159480 279978 159800 280046
rect 159480 279922 159550 279978
rect 159606 279922 159674 279978
rect 159730 279922 159800 279978
rect 159480 279888 159800 279922
rect 162738 280350 163358 297922
rect 163884 285684 163940 285694
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 138684 275698 138740 275708
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 132018 244350 132638 261922
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 138572 270658 138628 270668
rect 138572 238420 138628 270602
rect 138684 261716 138740 275642
rect 139096 274350 139416 274384
rect 139096 274294 139166 274350
rect 139222 274294 139290 274350
rect 139346 274294 139416 274350
rect 139096 274226 139416 274294
rect 139096 274170 139166 274226
rect 139222 274170 139290 274226
rect 139346 274170 139416 274226
rect 139096 274102 139416 274170
rect 139096 274046 139166 274102
rect 139222 274046 139290 274102
rect 139346 274046 139416 274102
rect 139096 273978 139416 274046
rect 139096 273922 139166 273978
rect 139222 273922 139290 273978
rect 139346 273922 139416 273978
rect 139096 273888 139416 273922
rect 144920 274350 145240 274384
rect 144920 274294 144990 274350
rect 145046 274294 145114 274350
rect 145170 274294 145240 274350
rect 144920 274226 145240 274294
rect 144920 274170 144990 274226
rect 145046 274170 145114 274226
rect 145170 274170 145240 274226
rect 144920 274102 145240 274170
rect 144920 274046 144990 274102
rect 145046 274046 145114 274102
rect 145170 274046 145240 274102
rect 144920 273978 145240 274046
rect 144920 273922 144990 273978
rect 145046 273922 145114 273978
rect 145170 273922 145240 273978
rect 144920 273888 145240 273922
rect 150744 274350 151064 274384
rect 150744 274294 150814 274350
rect 150870 274294 150938 274350
rect 150994 274294 151064 274350
rect 150744 274226 151064 274294
rect 150744 274170 150814 274226
rect 150870 274170 150938 274226
rect 150994 274170 151064 274226
rect 150744 274102 151064 274170
rect 150744 274046 150814 274102
rect 150870 274046 150938 274102
rect 150994 274046 151064 274102
rect 150744 273978 151064 274046
rect 150744 273922 150814 273978
rect 150870 273922 150938 273978
rect 150994 273922 151064 273978
rect 150744 273888 151064 273922
rect 156568 274350 156888 274384
rect 156568 274294 156638 274350
rect 156694 274294 156762 274350
rect 156818 274294 156888 274350
rect 156568 274226 156888 274294
rect 156568 274170 156638 274226
rect 156694 274170 156762 274226
rect 156818 274170 156888 274226
rect 156568 274102 156888 274170
rect 156568 274046 156638 274102
rect 156694 274046 156762 274102
rect 156818 274046 156888 274102
rect 156568 273978 156888 274046
rect 156568 273922 156638 273978
rect 156694 273922 156762 273978
rect 156818 273922 156888 273978
rect 156568 273888 156888 273922
rect 138684 261650 138740 261660
rect 162738 262350 163358 279922
rect 163436 282212 163492 282222
rect 163436 280738 163492 282156
rect 163436 267876 163492 280682
rect 163884 278938 163940 285628
rect 164108 284698 164164 284708
rect 163436 267810 163492 267820
rect 163772 275604 163828 275614
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 138572 238354 138628 238364
rect 159018 256350 159638 260964
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 132018 208350 132638 225922
rect 132018 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 132638 208350
rect 132018 208226 132638 208294
rect 132018 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 132638 208226
rect 132018 208102 132638 208170
rect 132018 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 132638 208102
rect 132018 207978 132638 208046
rect 132018 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 132638 207978
rect 132018 205590 132638 207922
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 205590 159638 219922
rect 162738 244350 163358 261922
rect 163772 261828 163828 275548
rect 163884 263844 163940 278882
rect 163996 280532 164052 280542
rect 163996 278038 164052 280476
rect 163996 265860 164052 277982
rect 164108 275940 164164 284642
rect 165452 282436 165508 377132
rect 166236 302596 166292 302606
rect 165452 282370 165508 282380
rect 165564 283078 165620 283088
rect 164108 275874 164164 275884
rect 165564 271908 165620 283022
rect 165564 271842 165620 271852
rect 163996 265794 164052 265804
rect 163884 263778 163940 263788
rect 163772 261762 163828 261772
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 166236 229908 166292 302540
rect 167132 277956 167188 469532
rect 168812 467908 168868 467918
rect 167916 304836 167972 304846
rect 167132 277890 167188 277900
rect 167244 281458 167300 281468
rect 167244 269892 167300 281402
rect 167244 269826 167300 269836
rect 167916 231588 167972 304780
rect 168812 279076 168868 467852
rect 170492 466228 170548 466238
rect 169596 320516 169652 320526
rect 169484 311556 169540 311566
rect 168812 279010 168868 279020
rect 168924 286498 168980 286508
rect 168924 278068 168980 286442
rect 168924 278002 168980 278012
rect 169036 283258 169092 283268
rect 168476 277318 168532 277328
rect 168476 275604 168532 277262
rect 168476 275538 168532 275548
rect 169036 273924 169092 283202
rect 169036 273858 169092 273868
rect 167916 231522 167972 231532
rect 166236 229842 166292 229852
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 208350 163358 225922
rect 169484 216244 169540 311500
rect 169484 216178 169540 216188
rect 169596 210868 169652 320460
rect 170492 280196 170548 466172
rect 171388 359716 171444 359726
rect 171388 349636 171444 359660
rect 171388 349570 171444 349580
rect 174524 310436 174580 310446
rect 174300 309316 174356 309326
rect 170492 280130 170548 280140
rect 171276 308196 171332 308206
rect 171276 218260 171332 308140
rect 171276 218194 171332 218204
rect 172956 301476 173012 301486
rect 169596 210802 169652 210812
rect 172956 209412 173012 301420
rect 174300 219940 174356 309260
rect 174300 219874 174356 219884
rect 174412 300356 174468 300366
rect 174412 209524 174468 300300
rect 174524 209636 174580 310380
rect 174636 266756 174692 573722
rect 179676 571978 179732 571988
rect 176316 569638 176372 569648
rect 174748 363076 174804 363086
rect 174748 359828 174804 363020
rect 174748 359762 174804 359772
rect 174860 361956 174916 361966
rect 174860 356356 174916 361900
rect 174860 356290 174916 356300
rect 176204 360836 176260 360846
rect 176204 353108 176260 360780
rect 176204 353042 176260 353052
rect 176204 313796 176260 313806
rect 174636 266690 174692 266700
rect 176092 294756 176148 294766
rect 176092 210644 176148 294700
rect 176092 210578 176148 210588
rect 176204 209748 176260 313740
rect 176316 265636 176372 569582
rect 177212 358596 177268 358606
rect 177212 338548 177268 358540
rect 177212 338482 177268 338492
rect 176316 265570 176372 265580
rect 177100 319396 177156 319406
rect 176988 254436 177044 254446
rect 176988 234298 177044 254380
rect 176988 234232 177044 234242
rect 177100 216356 177156 319340
rect 179564 317156 179620 317166
rect 177548 314916 177604 314926
rect 177212 299236 177268 299246
rect 177212 239652 177268 299180
rect 177212 239586 177268 239596
rect 177324 298116 177380 298126
rect 177324 224980 177380 298060
rect 177324 224914 177380 224924
rect 177436 296996 177492 297006
rect 177436 223412 177492 296940
rect 177548 239764 177604 314860
rect 177884 312676 177940 312686
rect 177772 303716 177828 303726
rect 177548 239698 177604 239708
rect 177660 295876 177716 295886
rect 177436 223346 177492 223356
rect 177660 221284 177716 295820
rect 177772 226324 177828 303660
rect 177884 233268 177940 312620
rect 179452 305956 179508 305966
rect 178892 286020 178948 286030
rect 178892 281988 178948 285964
rect 178892 236852 178948 281932
rect 178892 236786 178948 236796
rect 177884 233202 177940 233212
rect 177772 226258 177828 226268
rect 177660 221218 177716 221228
rect 179452 216468 179508 305900
rect 179452 216402 179508 216412
rect 177100 216290 177156 216300
rect 177548 213332 177604 213342
rect 177548 211798 177604 213276
rect 177548 211732 177604 211742
rect 179564 209860 179620 317100
rect 179676 271236 179732 571922
rect 180012 569818 180068 569828
rect 179900 279972 179956 279982
rect 179900 279658 179956 279916
rect 179900 279592 179956 279602
rect 179676 271170 179732 271180
rect 180012 263396 180068 569762
rect 184716 550788 184772 550798
rect 184604 543620 184660 543630
rect 180460 507780 180516 507790
rect 180012 263330 180068 263340
rect 180124 316036 180180 316046
rect 180012 262276 180068 262286
rect 179676 256676 179732 256686
rect 179676 218148 179732 256620
rect 179676 218082 179732 218092
rect 180012 212772 180068 262220
rect 180012 212706 180068 212716
rect 179564 209794 179620 209804
rect 176204 209682 176260 209692
rect 174524 209570 174580 209580
rect 174412 209458 174468 209468
rect 172956 209346 173012 209356
rect 180124 209076 180180 315980
rect 180236 307076 180292 307086
rect 180236 211092 180292 307020
rect 180460 288838 180516 507724
rect 180460 284004 180516 288782
rect 180572 500612 180628 500622
rect 180572 286020 180628 500556
rect 184604 399028 184660 543564
rect 184604 398962 184660 398972
rect 184716 397378 184772 550732
rect 186396 522116 186452 522126
rect 186284 421764 186340 421774
rect 184716 397312 184772 397322
rect 185612 414596 185668 414606
rect 184448 364350 184768 364384
rect 184448 364294 184518 364350
rect 184574 364294 184642 364350
rect 184698 364294 184768 364350
rect 184448 364226 184768 364294
rect 184448 364170 184518 364226
rect 184574 364170 184642 364226
rect 184698 364170 184768 364226
rect 184448 364102 184768 364170
rect 184448 364046 184518 364102
rect 184574 364046 184642 364102
rect 184698 364046 184768 364102
rect 184448 363978 184768 364046
rect 184448 363922 184518 363978
rect 184574 363922 184642 363978
rect 184698 363922 184768 363978
rect 184448 363888 184768 363922
rect 184448 346350 184768 346384
rect 184448 346294 184518 346350
rect 184574 346294 184642 346350
rect 184698 346294 184768 346350
rect 184448 346226 184768 346294
rect 184448 346170 184518 346226
rect 184574 346170 184642 346226
rect 184698 346170 184768 346226
rect 184448 346102 184768 346170
rect 184448 346046 184518 346102
rect 184574 346046 184642 346102
rect 184698 346046 184768 346102
rect 184448 345978 184768 346046
rect 184448 345922 184518 345978
rect 184574 345922 184642 345978
rect 184698 345922 184768 345978
rect 184448 345888 184768 345922
rect 184448 328350 184768 328384
rect 184448 328294 184518 328350
rect 184574 328294 184642 328350
rect 184698 328294 184768 328350
rect 184448 328226 184768 328294
rect 184448 328170 184518 328226
rect 184574 328170 184642 328226
rect 184698 328170 184768 328226
rect 184448 328102 184768 328170
rect 184448 328046 184518 328102
rect 184574 328046 184642 328102
rect 184698 328046 184768 328102
rect 184448 327978 184768 328046
rect 184448 327922 184518 327978
rect 184574 327922 184642 327978
rect 184698 327922 184768 327978
rect 184448 327888 184768 327922
rect 184448 310350 184768 310384
rect 184448 310294 184518 310350
rect 184574 310294 184642 310350
rect 184698 310294 184768 310350
rect 184448 310226 184768 310294
rect 184448 310170 184518 310226
rect 184574 310170 184642 310226
rect 184698 310170 184768 310226
rect 184448 310102 184768 310170
rect 184448 310046 184518 310102
rect 184574 310046 184642 310102
rect 184698 310046 184768 310102
rect 184448 309978 184768 310046
rect 184448 309922 184518 309978
rect 184574 309922 184642 309978
rect 184698 309922 184768 309978
rect 184448 309888 184768 309922
rect 184448 292350 184768 292384
rect 184448 292294 184518 292350
rect 184574 292294 184642 292350
rect 184698 292294 184768 292350
rect 184448 292226 184768 292294
rect 184448 292170 184518 292226
rect 184574 292170 184642 292226
rect 184698 292170 184768 292226
rect 184448 292102 184768 292170
rect 184448 292046 184518 292102
rect 184574 292046 184642 292102
rect 184698 292046 184768 292102
rect 184448 291978 184768 292046
rect 184448 291922 184518 291978
rect 184574 291922 184642 291978
rect 184698 291922 184768 291978
rect 184448 291888 184768 291922
rect 184828 290638 184884 290648
rect 180572 285954 180628 285964
rect 183932 287218 183988 287228
rect 180460 283938 180516 283948
rect 183932 279658 183988 287162
rect 180572 265438 180628 265448
rect 180572 265076 180628 265382
rect 180572 265010 180628 265020
rect 180684 261156 180740 261166
rect 180684 261052 180740 261062
rect 180684 260038 180740 260048
rect 180684 259944 180740 259980
rect 180684 258958 180740 258968
rect 180684 258850 180740 258860
rect 180572 257236 180628 257246
rect 180572 257158 180628 257180
rect 180572 257092 180628 257102
rect 180348 255556 180404 255566
rect 180348 214788 180404 255500
rect 180572 252756 180628 252766
rect 180572 252298 180628 252700
rect 180572 252232 180628 252242
rect 180684 252196 180740 252206
rect 180684 252118 180740 252140
rect 180684 252052 180740 252062
rect 183932 235172 183988 279602
rect 184448 274350 184768 274384
rect 184448 274294 184518 274350
rect 184574 274294 184642 274350
rect 184698 274294 184768 274350
rect 184448 274226 184768 274294
rect 184448 274170 184518 274226
rect 184574 274170 184642 274226
rect 184698 274170 184768 274226
rect 184448 274102 184768 274170
rect 184448 274046 184518 274102
rect 184574 274046 184642 274102
rect 184698 274046 184768 274102
rect 184448 273978 184768 274046
rect 184448 273922 184518 273978
rect 184574 273922 184642 273978
rect 184698 273922 184768 273978
rect 184448 273888 184768 273922
rect 184448 256350 184768 256384
rect 184448 256294 184518 256350
rect 184574 256294 184642 256350
rect 184698 256294 184768 256350
rect 184448 256226 184768 256294
rect 184448 256170 184518 256226
rect 184574 256170 184642 256226
rect 184698 256170 184768 256226
rect 184448 256102 184768 256170
rect 184448 256046 184518 256102
rect 184574 256046 184642 256102
rect 184698 256046 184768 256102
rect 184448 255978 184768 256046
rect 184448 255922 184518 255978
rect 184574 255922 184642 255978
rect 184698 255922 184768 255978
rect 184448 255888 184768 255922
rect 184828 240100 184884 290582
rect 185612 290638 185668 414540
rect 186284 394212 186340 421708
rect 186284 394146 186340 394156
rect 186396 390964 186452 522060
rect 187292 493444 187348 493454
rect 186396 390898 186452 390908
rect 187180 479108 187236 479118
rect 187180 393204 187236 479052
rect 185612 290572 185668 290582
rect 187180 285778 187236 393148
rect 187292 287218 187348 493388
rect 188076 486276 188132 486286
rect 187964 471940 188020 471950
rect 187852 464772 187908 464782
rect 187740 457604 187796 457614
rect 187292 287152 187348 287162
rect 187404 450436 187460 450446
rect 187180 285712 187236 285722
rect 187292 283798 187348 283808
rect 187292 283078 187348 283742
rect 187292 283012 187348 283022
rect 186396 282178 186452 282188
rect 186396 280738 186452 282122
rect 187404 282178 187460 450380
rect 187404 282112 187460 282122
rect 187516 443268 187572 443278
rect 184828 240034 184884 240044
rect 186284 279658 186340 279668
rect 186284 278938 186340 279602
rect 186284 239428 186340 278882
rect 186284 239362 186340 239372
rect 186396 239316 186452 280682
rect 187516 278038 187572 443212
rect 187628 436100 187684 436110
rect 187628 279658 187684 436044
rect 187740 281458 187796 457548
rect 187852 283798 187908 464716
rect 187852 283732 187908 283742
rect 187964 283258 188020 471884
rect 188076 286498 188132 486220
rect 188972 409668 189028 590156
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 189420 576436 189476 576446
rect 189196 575428 189252 575438
rect 188972 409602 189028 409612
rect 189084 428932 189140 428942
rect 188076 286432 188132 286442
rect 188076 285778 188132 285788
rect 188076 284698 188132 285722
rect 188076 284632 188132 284642
rect 187964 283192 188020 283202
rect 187740 281392 187796 281402
rect 187628 279592 187684 279602
rect 187404 261118 187460 261128
rect 186396 239250 186452 239260
rect 187292 258958 187348 258968
rect 183932 235106 183988 235116
rect 180348 214722 180404 214732
rect 187292 214676 187348 258902
rect 187404 236628 187460 261062
rect 187516 238308 187572 277982
rect 188076 277318 188132 277328
rect 187516 238242 187572 238252
rect 187628 260038 187684 260048
rect 187404 236562 187460 236572
rect 187628 231058 187684 259982
rect 188076 235732 188132 277262
rect 189084 277318 189140 428876
rect 189196 404218 189252 575372
rect 189196 404152 189252 404162
rect 189308 574868 189364 574878
rect 189308 402612 189364 574812
rect 189308 402546 189364 402556
rect 189420 399252 189476 576380
rect 189420 399186 189476 399196
rect 189532 567924 189588 567934
rect 189420 390538 189476 390548
rect 189084 277252 189140 277262
rect 189308 289018 189364 289028
rect 188076 235666 188132 235676
rect 189308 234948 189364 288962
rect 189420 235844 189476 390482
rect 189532 382900 189588 567868
rect 189532 382834 189588 382844
rect 189738 562350 190358 579922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 202972 591220 203028 591230
rect 202860 587300 202916 587310
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 190428 575204 190484 575214
rect 190428 567028 190484 575148
rect 192892 573300 192948 573310
rect 192668 571284 192724 571294
rect 192556 569940 192612 569950
rect 190428 566962 190484 566972
rect 191324 567252 191380 567262
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 189738 544350 190358 561922
rect 189738 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 190358 544350
rect 189738 544226 190358 544294
rect 189738 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 190358 544226
rect 189738 544102 190358 544170
rect 189738 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 190358 544102
rect 189738 543978 190358 544046
rect 189738 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 190358 543978
rect 189738 526350 190358 543922
rect 189738 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 190358 526350
rect 189738 526226 190358 526294
rect 189738 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 190358 526226
rect 189738 526102 190358 526170
rect 189738 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 190358 526102
rect 189738 525978 190358 526046
rect 189738 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 190358 525978
rect 189738 508350 190358 525922
rect 189738 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 190358 508350
rect 189738 508226 190358 508294
rect 189738 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 190358 508226
rect 189738 508102 190358 508170
rect 189738 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 190358 508102
rect 189738 507978 190358 508046
rect 189738 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 190358 507978
rect 189738 490350 190358 507922
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 189738 454350 190358 471922
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 189738 418350 190358 435922
rect 189738 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 190358 418350
rect 189738 418226 190358 418294
rect 189738 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 190358 418226
rect 189738 418102 190358 418170
rect 189738 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 190358 418102
rect 189738 417978 190358 418046
rect 189738 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 190358 417978
rect 189738 400350 190358 417922
rect 191324 403956 191380 567196
rect 191324 403890 191380 403900
rect 191436 567140 191492 567150
rect 189738 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 190358 400350
rect 189738 400226 190358 400294
rect 189738 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 190358 400226
rect 189738 400102 190358 400170
rect 189738 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 190358 400102
rect 189738 399978 190358 400046
rect 189738 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 190358 399978
rect 189738 382350 190358 399922
rect 191436 390740 191492 567084
rect 192556 407204 192612 569884
rect 192668 409780 192724 571228
rect 192668 409714 192724 409724
rect 192780 568260 192836 568270
rect 192556 407138 192612 407148
rect 192780 404740 192836 568204
rect 192780 404674 192836 404684
rect 192892 400820 192948 573244
rect 193116 572180 193172 572190
rect 192892 400754 192948 400764
rect 193004 571508 193060 571518
rect 193004 397908 193060 571452
rect 193004 397842 193060 397852
rect 192444 393316 192500 393326
rect 191548 392532 191604 392542
rect 191548 391618 191604 392476
rect 191548 391552 191604 391562
rect 191436 390674 191492 390684
rect 189738 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 190358 382350
rect 189738 382226 190358 382294
rect 189738 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 190358 382226
rect 189738 382102 190358 382170
rect 189738 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 190358 382102
rect 189738 381978 190358 382046
rect 189738 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 190358 381978
rect 189420 235778 189476 235788
rect 189532 380548 189588 380558
rect 189308 234882 189364 234892
rect 187628 230992 187684 231002
rect 187292 214610 187348 214620
rect 180236 211026 180292 211036
rect 189532 209972 189588 380492
rect 189532 209906 189588 209916
rect 189738 364350 190358 381922
rect 189738 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 190358 364350
rect 189738 364226 190358 364294
rect 189738 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 190358 364226
rect 189738 364102 190358 364170
rect 189738 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 190358 364102
rect 189738 363978 190358 364046
rect 189738 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 190358 363978
rect 189738 346350 190358 363922
rect 189738 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 190358 346350
rect 189738 346226 190358 346294
rect 189738 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 190358 346226
rect 189738 346102 190358 346170
rect 189738 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 190358 346102
rect 189738 345978 190358 346046
rect 189738 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 190358 345978
rect 189738 328350 190358 345922
rect 189738 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 190358 328350
rect 189738 328226 190358 328294
rect 189738 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 190358 328226
rect 189738 328102 190358 328170
rect 189738 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 190358 328102
rect 189738 327978 190358 328046
rect 189738 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 190358 327978
rect 189738 310350 190358 327922
rect 189738 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 190358 310350
rect 189738 310226 190358 310294
rect 189738 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 190358 310226
rect 189738 310102 190358 310170
rect 189738 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 190358 310102
rect 189738 309978 190358 310046
rect 189738 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 190358 309978
rect 189738 292350 190358 309922
rect 189738 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 190358 292350
rect 189738 292226 190358 292294
rect 189738 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 190358 292226
rect 189738 292102 190358 292170
rect 189738 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 190358 292102
rect 189738 291978 190358 292046
rect 189738 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 190358 291978
rect 189738 274350 190358 291922
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189738 256350 190358 273922
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189738 220350 190358 237922
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 180124 209010 180180 209020
rect 162738 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163358 208350
rect 162738 208226 163358 208294
rect 162738 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163358 208226
rect 162738 208102 163358 208170
rect 162738 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163358 208102
rect 162738 207978 163358 208046
rect 162738 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163358 207978
rect 162738 205590 163358 207922
rect 189738 205590 190358 219922
rect 190764 379540 190820 379550
rect 190764 211078 190820 379484
rect 191324 379540 191380 379550
rect 191324 212518 191380 379484
rect 192108 379540 192164 379550
rect 191548 236852 191604 236862
rect 191548 236292 191604 236796
rect 191548 236226 191604 236236
rect 192108 215938 192164 379484
rect 192444 219604 192500 393260
rect 193116 392532 193172 572124
rect 193116 392466 193172 392476
rect 193458 568350 194078 585922
rect 196476 587188 196532 587198
rect 196252 573188 196308 573198
rect 196028 568708 196084 568718
rect 193458 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 194078 568350
rect 193458 568226 194078 568294
rect 193458 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 194078 568226
rect 193458 568102 194078 568170
rect 193458 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 194078 568102
rect 193458 567978 194078 568046
rect 193458 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 194078 567978
rect 193458 550350 194078 567922
rect 195916 568484 195972 568494
rect 194448 562350 194768 562384
rect 194448 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 194768 562350
rect 194448 562226 194768 562294
rect 194448 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 194768 562226
rect 194448 562102 194768 562170
rect 194448 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 194768 562102
rect 194448 561978 194768 562046
rect 194448 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 194768 561978
rect 194448 561888 194768 561922
rect 193458 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 194078 550350
rect 193458 550226 194078 550294
rect 193458 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 194078 550226
rect 193458 550102 194078 550170
rect 193458 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 194078 550102
rect 193458 549978 194078 550046
rect 193458 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 194078 549978
rect 193458 532350 194078 549922
rect 194448 544350 194768 544384
rect 194448 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 194768 544350
rect 194448 544226 194768 544294
rect 194448 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 194768 544226
rect 194448 544102 194768 544170
rect 194448 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 194768 544102
rect 194448 543978 194768 544046
rect 194448 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 194768 543978
rect 194448 543888 194768 543922
rect 193458 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 194078 532350
rect 193458 532226 194078 532294
rect 193458 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 194078 532226
rect 193458 532102 194078 532170
rect 193458 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 194078 532102
rect 193458 531978 194078 532046
rect 193458 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 194078 531978
rect 193458 514350 194078 531922
rect 194448 526350 194768 526384
rect 194448 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 194768 526350
rect 194448 526226 194768 526294
rect 194448 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 194768 526226
rect 194448 526102 194768 526170
rect 194448 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 194768 526102
rect 194448 525978 194768 526046
rect 194448 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 194768 525978
rect 194448 525888 194768 525922
rect 193458 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 194078 514350
rect 193458 514226 194078 514294
rect 193458 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 194078 514226
rect 193458 514102 194078 514170
rect 193458 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 194078 514102
rect 193458 513978 194078 514046
rect 193458 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 194078 513978
rect 193458 496350 194078 513922
rect 194448 508350 194768 508384
rect 194448 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 194768 508350
rect 194448 508226 194768 508294
rect 194448 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 194768 508226
rect 194448 508102 194768 508170
rect 194448 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 194768 508102
rect 194448 507978 194768 508046
rect 194448 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 194768 507978
rect 194448 507888 194768 507922
rect 193458 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 194078 496350
rect 193458 496226 194078 496294
rect 193458 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 194078 496226
rect 193458 496102 194078 496170
rect 193458 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 194078 496102
rect 193458 495978 194078 496046
rect 193458 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 194078 495978
rect 193458 478350 194078 495922
rect 194448 490350 194768 490384
rect 194448 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 194768 490350
rect 194448 490226 194768 490294
rect 194448 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 194768 490226
rect 194448 490102 194768 490170
rect 194448 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 194768 490102
rect 194448 489978 194768 490046
rect 194448 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 194768 489978
rect 194448 489888 194768 489922
rect 193458 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 194078 478350
rect 193458 478226 194078 478294
rect 193458 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 194078 478226
rect 193458 478102 194078 478170
rect 193458 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 194078 478102
rect 193458 477978 194078 478046
rect 193458 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 194078 477978
rect 193458 460350 194078 477922
rect 194448 472350 194768 472384
rect 194448 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 194768 472350
rect 194448 472226 194768 472294
rect 194448 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 194768 472226
rect 194448 472102 194768 472170
rect 194448 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 194768 472102
rect 194448 471978 194768 472046
rect 194448 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 194768 471978
rect 194448 471888 194768 471922
rect 193458 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 194078 460350
rect 193458 460226 194078 460294
rect 193458 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 194078 460226
rect 193458 460102 194078 460170
rect 193458 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 194078 460102
rect 193458 459978 194078 460046
rect 193458 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 194078 459978
rect 193458 442350 194078 459922
rect 194448 454350 194768 454384
rect 194448 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 194768 454350
rect 194448 454226 194768 454294
rect 194448 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 194768 454226
rect 194448 454102 194768 454170
rect 194448 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 194768 454102
rect 194448 453978 194768 454046
rect 194448 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 194768 453978
rect 194448 453888 194768 453922
rect 193458 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 194078 442350
rect 193458 442226 194078 442294
rect 193458 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 194078 442226
rect 193458 442102 194078 442170
rect 193458 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 194078 442102
rect 193458 441978 194078 442046
rect 193458 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 194078 441978
rect 193458 424350 194078 441922
rect 194448 436350 194768 436384
rect 194448 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 194768 436350
rect 194448 436226 194768 436294
rect 194448 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 194768 436226
rect 194448 436102 194768 436170
rect 194448 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 194768 436102
rect 194448 435978 194768 436046
rect 194448 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 194768 435978
rect 194448 435888 194768 435922
rect 193458 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 194078 424350
rect 193458 424226 194078 424294
rect 193458 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 194078 424226
rect 193458 424102 194078 424170
rect 193458 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 194078 424102
rect 193458 423978 194078 424046
rect 193458 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 194078 423978
rect 193458 406350 194078 423922
rect 194448 418350 194768 418384
rect 194448 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 194768 418350
rect 194448 418226 194768 418294
rect 194448 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 194768 418226
rect 194448 418102 194768 418170
rect 194448 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 194768 418102
rect 194448 417978 194768 418046
rect 194448 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 194768 417978
rect 194448 417888 194768 417922
rect 195916 407876 195972 568428
rect 195916 407810 195972 407820
rect 196028 406756 196084 568652
rect 196028 406690 196084 406700
rect 196140 568372 196196 568382
rect 193458 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 194078 406350
rect 193458 406226 194078 406294
rect 193458 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 194078 406226
rect 193458 406102 194078 406170
rect 193458 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 194078 406102
rect 193458 405978 194078 406046
rect 193458 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 194078 405978
rect 192892 391618 192948 391628
rect 192556 389956 192612 389966
rect 192556 236292 192612 389900
rect 192556 236226 192612 236236
rect 192668 379540 192724 379550
rect 192444 219538 192500 219548
rect 192668 219178 192724 379484
rect 192892 225988 192948 391562
rect 193458 388350 194078 405922
rect 196140 404628 196196 568316
rect 196140 404562 196196 404572
rect 196252 404068 196308 573132
rect 196252 404002 196308 404012
rect 196364 569828 196420 569838
rect 196364 401044 196420 569772
rect 196476 406532 196532 587132
rect 202748 576324 202804 576334
rect 201180 574756 201236 574766
rect 198044 574644 198100 574654
rect 197820 573524 197876 573534
rect 197708 573412 197764 573422
rect 197596 566218 197652 566228
rect 197596 407540 197652 566162
rect 197596 407474 197652 407484
rect 196476 406466 196532 406476
rect 197708 404404 197764 573356
rect 197708 404338 197764 404348
rect 196364 400978 196420 400988
rect 197596 401604 197652 401614
rect 194908 396004 194964 396014
rect 194908 394884 194964 395948
rect 194908 394818 194964 394828
rect 196252 394884 196308 394894
rect 193458 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 194078 388350
rect 193458 388226 194078 388294
rect 193458 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 194078 388226
rect 193458 388102 194078 388170
rect 193458 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 194078 388102
rect 193458 387978 194078 388046
rect 193458 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 194078 387978
rect 193340 379540 193396 379550
rect 192892 225922 192948 225932
rect 193004 379316 193060 379326
rect 192668 219112 192724 219122
rect 192108 215872 192164 215882
rect 193004 214900 193060 379260
rect 193340 216580 193396 379484
rect 193340 216514 193396 216524
rect 193458 370350 194078 387922
rect 196028 388388 196084 388398
rect 193458 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 194078 370350
rect 193458 370226 194078 370294
rect 193458 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 194078 370226
rect 193458 370102 194078 370170
rect 193458 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 194078 370102
rect 193458 369978 194078 370046
rect 193458 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 194078 369978
rect 193458 352350 194078 369922
rect 193458 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 194078 352350
rect 193458 352226 194078 352294
rect 193458 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 194078 352226
rect 193458 352102 194078 352170
rect 193458 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 194078 352102
rect 193458 351978 194078 352046
rect 193458 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 194078 351978
rect 193458 334350 194078 351922
rect 193458 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 194078 334350
rect 193458 334226 194078 334294
rect 193458 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 194078 334226
rect 193458 334102 194078 334170
rect 193458 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 194078 334102
rect 193458 333978 194078 334046
rect 193458 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 194078 333978
rect 193458 316350 194078 333922
rect 193458 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 194078 316350
rect 193458 316226 194078 316294
rect 193458 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 194078 316226
rect 193458 316102 194078 316170
rect 193458 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 194078 316102
rect 193458 315978 194078 316046
rect 193458 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 194078 315978
rect 193458 298350 194078 315922
rect 193458 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 194078 298350
rect 193458 298226 194078 298294
rect 193458 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 194078 298226
rect 193458 298102 194078 298170
rect 193458 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 194078 298102
rect 193458 297978 194078 298046
rect 193458 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 194078 297978
rect 193458 280350 194078 297922
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193458 262350 194078 279922
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 193458 244350 194078 261922
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 193004 214834 193060 214844
rect 191324 212452 191380 212462
rect 190764 211012 190820 211022
rect 193458 208350 194078 225922
rect 194684 379540 194740 379550
rect 194684 222964 194740 379484
rect 195244 379540 195300 379550
rect 195244 289018 195300 379484
rect 195244 288952 195300 288962
rect 196028 288838 196084 388332
rect 196028 288772 196084 288782
rect 196140 379316 196196 379326
rect 195916 286498 195972 286508
rect 195692 285778 195748 285788
rect 195692 232708 195748 285722
rect 195916 282358 195972 286442
rect 195692 232642 195748 232652
rect 195804 257158 195860 257168
rect 194684 222898 194740 222908
rect 195804 218372 195860 257102
rect 195916 246898 195972 282302
rect 195916 246832 195972 246842
rect 196140 229460 196196 379260
rect 196252 239338 196308 394828
rect 196476 391748 196532 391758
rect 196252 239272 196308 239282
rect 196364 379540 196420 379550
rect 196140 229394 196196 229404
rect 195804 218306 195860 218316
rect 196364 214452 196420 379484
rect 196364 214386 196420 214396
rect 193458 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 194078 208350
rect 193458 208226 194078 208294
rect 193458 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 194078 208226
rect 193458 208102 194078 208170
rect 193458 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 194078 208102
rect 193458 207978 194078 208046
rect 193458 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 194078 207978
rect 193458 205590 194078 207922
rect 196476 206578 196532 391692
rect 197484 388052 197540 388062
rect 197484 386820 197540 387996
rect 197484 386754 197540 386764
rect 197372 383236 197428 383246
rect 197372 240548 197428 383180
rect 197372 240482 197428 240492
rect 197596 231700 197652 401548
rect 197820 399364 197876 573468
rect 197820 399298 197876 399308
rect 197932 571620 197988 571630
rect 197932 396004 197988 571564
rect 197932 395938 197988 395948
rect 198044 396452 198100 574588
rect 199612 573636 199668 573646
rect 199388 571732 199444 571742
rect 198044 395892 198100 396396
rect 198044 395826 198100 395836
rect 198156 568036 198212 568046
rect 197708 392338 197764 392348
rect 197708 382228 197764 392282
rect 197932 386820 197988 386830
rect 197708 382162 197764 382172
rect 197820 386578 197876 386588
rect 197708 380660 197764 380670
rect 197708 236740 197764 380604
rect 197708 236674 197764 236684
rect 197820 233492 197876 386522
rect 197820 233426 197876 233436
rect 197596 231634 197652 231644
rect 197932 224756 197988 386764
rect 198156 382228 198212 567980
rect 199276 567364 199332 567374
rect 199276 408996 199332 567308
rect 199276 408930 199332 408940
rect 199388 407764 199444 571676
rect 199388 407698 199444 407708
rect 199500 569940 199556 569950
rect 199500 404180 199556 569884
rect 199612 404852 199668 573580
rect 200956 572068 201012 572078
rect 199836 571396 199892 571406
rect 199612 404786 199668 404796
rect 199724 571258 199780 571268
rect 199500 404114 199556 404124
rect 199276 399140 199332 399150
rect 199276 398244 199332 399084
rect 198156 382162 198212 382172
rect 199052 383796 199108 383806
rect 198156 380098 198212 380108
rect 198044 233492 198100 233502
rect 198044 232820 198100 233436
rect 198044 232754 198100 232764
rect 197932 224690 197988 224700
rect 198156 221508 198212 380042
rect 198940 288838 198996 288848
rect 198940 236180 198996 288782
rect 198940 236114 198996 236124
rect 199052 233380 199108 383740
rect 199164 379738 199220 379748
rect 199164 283798 199220 379682
rect 199164 240436 199220 283742
rect 199276 253738 199332 398188
rect 199612 390964 199668 390974
rect 199500 390404 199556 390414
rect 199388 390292 199444 390302
rect 199388 282358 199444 390236
rect 199388 282292 199444 282302
rect 199276 253672 199332 253682
rect 199164 240370 199220 240380
rect 199276 252298 199332 252308
rect 199052 233314 199108 233324
rect 198156 221442 198212 221452
rect 199276 212660 199332 252242
rect 199388 246898 199444 246908
rect 199388 236516 199444 246842
rect 199388 236450 199444 236460
rect 199500 221396 199556 390348
rect 199500 221330 199556 221340
rect 199612 389818 199668 390908
rect 199612 217558 199668 389762
rect 199724 382228 199780 571202
rect 199836 382340 199892 571340
rect 200732 568148 200788 568158
rect 199836 382274 199892 382284
rect 199948 404218 200004 404228
rect 199724 382162 199780 382172
rect 199948 382228 200004 404162
rect 199948 382162 200004 382172
rect 199808 370350 200128 370384
rect 199808 370294 199878 370350
rect 199934 370294 200002 370350
rect 200058 370294 200128 370350
rect 199808 370226 200128 370294
rect 199808 370170 199878 370226
rect 199934 370170 200002 370226
rect 200058 370170 200128 370226
rect 199808 370102 200128 370170
rect 199808 370046 199878 370102
rect 199934 370046 200002 370102
rect 200058 370046 200128 370102
rect 199808 369978 200128 370046
rect 199808 369922 199878 369978
rect 199934 369922 200002 369978
rect 200058 369922 200128 369978
rect 199808 369888 200128 369922
rect 199808 352350 200128 352384
rect 199808 352294 199878 352350
rect 199934 352294 200002 352350
rect 200058 352294 200128 352350
rect 199808 352226 200128 352294
rect 199808 352170 199878 352226
rect 199934 352170 200002 352226
rect 200058 352170 200128 352226
rect 199808 352102 200128 352170
rect 199808 352046 199878 352102
rect 199934 352046 200002 352102
rect 200058 352046 200128 352102
rect 199808 351978 200128 352046
rect 199808 351922 199878 351978
rect 199934 351922 200002 351978
rect 200058 351922 200128 351978
rect 199808 351888 200128 351922
rect 199808 334350 200128 334384
rect 199808 334294 199878 334350
rect 199934 334294 200002 334350
rect 200058 334294 200128 334350
rect 199808 334226 200128 334294
rect 199808 334170 199878 334226
rect 199934 334170 200002 334226
rect 200058 334170 200128 334226
rect 199808 334102 200128 334170
rect 199808 334046 199878 334102
rect 199934 334046 200002 334102
rect 200058 334046 200128 334102
rect 199808 333978 200128 334046
rect 199808 333922 199878 333978
rect 199934 333922 200002 333978
rect 200058 333922 200128 333978
rect 199808 333888 200128 333922
rect 199808 316350 200128 316384
rect 199808 316294 199878 316350
rect 199934 316294 200002 316350
rect 200058 316294 200128 316350
rect 199808 316226 200128 316294
rect 199808 316170 199878 316226
rect 199934 316170 200002 316226
rect 200058 316170 200128 316226
rect 199808 316102 200128 316170
rect 199808 316046 199878 316102
rect 199934 316046 200002 316102
rect 200058 316046 200128 316102
rect 199808 315978 200128 316046
rect 199808 315922 199878 315978
rect 199934 315922 200002 315978
rect 200058 315922 200128 315978
rect 199808 315888 200128 315922
rect 199808 298350 200128 298384
rect 199808 298294 199878 298350
rect 199934 298294 200002 298350
rect 200058 298294 200128 298350
rect 199808 298226 200128 298294
rect 199808 298170 199878 298226
rect 199934 298170 200002 298226
rect 200058 298170 200128 298226
rect 199808 298102 200128 298170
rect 199808 298046 199878 298102
rect 199934 298046 200002 298102
rect 200058 298046 200128 298102
rect 199808 297978 200128 298046
rect 199808 297922 199878 297978
rect 199934 297922 200002 297978
rect 200058 297922 200128 297978
rect 199808 297888 200128 297922
rect 199808 280350 200128 280384
rect 199808 280294 199878 280350
rect 199934 280294 200002 280350
rect 200058 280294 200128 280350
rect 199808 280226 200128 280294
rect 199808 280170 199878 280226
rect 199934 280170 200002 280226
rect 200058 280170 200128 280226
rect 199808 280102 200128 280170
rect 199808 280046 199878 280102
rect 199934 280046 200002 280102
rect 200058 280046 200128 280102
rect 199808 279978 200128 280046
rect 199808 279922 199878 279978
rect 199934 279922 200002 279978
rect 200058 279922 200128 279978
rect 199808 279888 200128 279922
rect 200732 265438 200788 568092
rect 200956 398132 201012 572012
rect 201068 571956 201124 571966
rect 201068 409220 201124 571900
rect 201180 409332 201236 574700
rect 201180 409266 201236 409276
rect 201292 571844 201348 571854
rect 201068 409154 201124 409164
rect 200956 398066 201012 398076
rect 201292 397684 201348 571788
rect 202412 570358 202468 570368
rect 201516 570052 201572 570062
rect 201292 397618 201348 397628
rect 201404 400708 201460 400718
rect 201404 399924 201460 400652
rect 201068 390852 201124 390862
rect 201068 389998 201124 390796
rect 200732 265372 200788 265382
rect 200844 383158 200900 383168
rect 199808 262350 200128 262384
rect 199808 262294 199878 262350
rect 199934 262294 200002 262350
rect 200058 262294 200128 262350
rect 199808 262226 200128 262294
rect 199808 262170 199878 262226
rect 199934 262170 200002 262226
rect 200058 262170 200128 262226
rect 199808 262102 200128 262170
rect 199808 262046 199878 262102
rect 199934 262046 200002 262102
rect 200058 262046 200128 262102
rect 199808 261978 200128 262046
rect 199808 261922 199878 261978
rect 199934 261922 200002 261978
rect 200058 261922 200128 261978
rect 199808 261888 200128 261922
rect 200732 253738 200788 253748
rect 199808 244350 200128 244384
rect 199808 244294 199878 244350
rect 199934 244294 200002 244350
rect 200058 244294 200128 244350
rect 199808 244226 200128 244294
rect 199808 244170 199878 244226
rect 199934 244170 200002 244226
rect 200058 244170 200128 244226
rect 199808 244102 200128 244170
rect 199808 244046 199878 244102
rect 199934 244046 200002 244102
rect 200058 244046 200128 244102
rect 199808 243978 200128 244046
rect 199808 243922 199878 243978
rect 199934 243922 200002 243978
rect 200058 243922 200128 243978
rect 199808 243888 200128 243922
rect 200732 221060 200788 253682
rect 200844 222598 200900 383102
rect 201068 351118 201124 389942
rect 201292 390516 201348 390526
rect 201068 351052 201124 351062
rect 201180 388836 201236 388846
rect 201068 307378 201124 307388
rect 201068 305938 201124 307322
rect 201068 231140 201124 305882
rect 201180 300898 201236 388780
rect 201180 300832 201236 300842
rect 201068 231074 201124 231084
rect 201180 265618 201236 265628
rect 201180 226100 201236 265562
rect 201180 226034 201236 226044
rect 201292 224218 201348 390460
rect 201292 224152 201348 224162
rect 200844 222532 200900 222542
rect 200732 220994 200788 221004
rect 199612 217492 199668 217502
rect 201404 214138 201460 399868
rect 201516 382452 201572 569996
rect 201516 382386 201572 382396
rect 202300 410698 202356 410708
rect 202300 410004 202356 410642
rect 201628 351118 201684 351128
rect 201628 283798 201684 351062
rect 201516 283742 201684 283798
rect 201740 300898 201796 300908
rect 201516 227638 201572 283742
rect 201740 265618 201796 300842
rect 201740 265552 201796 265562
rect 201516 227572 201572 227582
rect 202300 222852 202356 409948
rect 202412 404964 202468 570302
rect 202412 307378 202468 404908
rect 202524 570164 202580 570174
rect 202524 404292 202580 570108
rect 202524 404226 202580 404236
rect 202636 568596 202692 568606
rect 202636 400708 202692 568540
rect 202748 406738 202804 576268
rect 202860 409556 202916 587244
rect 202972 409780 203028 591164
rect 203196 590884 203252 590894
rect 202972 409714 203028 409724
rect 203084 590660 203140 590670
rect 202860 409490 202916 409500
rect 203084 409444 203140 590604
rect 203084 409378 203140 409388
rect 203196 407204 203252 590828
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 203196 407138 203252 407148
rect 203532 570276 203588 570286
rect 203308 406738 203364 406748
rect 202748 406682 203308 406738
rect 202636 400642 202692 400652
rect 202748 405860 202804 405870
rect 202748 405076 202804 405804
rect 202748 396508 202804 405020
rect 202860 398132 202916 398142
rect 202860 397796 202916 398076
rect 202860 397730 202916 397740
rect 202748 396452 203028 396508
rect 202524 387298 202580 387308
rect 202524 376318 202580 387242
rect 202748 384958 202804 384968
rect 202524 376252 202580 376262
rect 202636 377938 202692 377948
rect 202636 372178 202692 377882
rect 202636 372112 202692 372122
rect 202412 307312 202468 307322
rect 202524 283258 202580 283268
rect 202412 281458 202468 281468
rect 202412 240100 202468 281402
rect 202524 240548 202580 283202
rect 202524 240482 202580 240492
rect 202636 252118 202692 252128
rect 202412 240034 202468 240044
rect 202524 235172 202580 235182
rect 202524 234388 202580 235116
rect 202524 234322 202580 234332
rect 202300 222786 202356 222796
rect 202636 215012 202692 252062
rect 202748 235172 202804 384902
rect 202748 235106 202804 235116
rect 202860 382676 202916 382686
rect 202860 226548 202916 382620
rect 202972 236404 203028 396452
rect 203308 390538 203364 406682
rect 203532 397572 203588 570220
rect 220458 568502 221078 579922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 568502 224798 585922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 568502 251798 579922
rect 253708 590212 253764 590222
rect 253708 570358 253764 590156
rect 253708 570292 253764 570302
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 568502 255518 585922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 568502 282518 579922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 568502 286238 585922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 568502 313238 579922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 568502 316958 585922
rect 341068 590212 341124 590222
rect 341068 571978 341124 590156
rect 341068 571912 341124 571922
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 568502 343958 579922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 568502 347678 585922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 568502 374678 579922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 568502 378398 585922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 568502 405398 579922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 568502 409118 585922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 568502 436118 579922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 568502 439838 585922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 568502 466838 579922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 568502 470558 585922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 478828 575204 478884 575214
rect 225168 562350 225488 562384
rect 225168 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 225488 562350
rect 225168 562226 225488 562294
rect 225168 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 225488 562226
rect 225168 562102 225488 562170
rect 225168 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 225488 562102
rect 225168 561978 225488 562046
rect 225168 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 225488 561978
rect 225168 561888 225488 561922
rect 255888 562350 256208 562384
rect 255888 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 256208 562350
rect 255888 562226 256208 562294
rect 255888 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 256208 562226
rect 255888 562102 256208 562170
rect 255888 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 256208 562102
rect 255888 561978 256208 562046
rect 255888 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 256208 561978
rect 255888 561888 256208 561922
rect 286608 562350 286928 562384
rect 286608 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 286928 562350
rect 286608 562226 286928 562294
rect 286608 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 286928 562226
rect 286608 562102 286928 562170
rect 286608 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 286928 562102
rect 286608 561978 286928 562046
rect 286608 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 286928 561978
rect 286608 561888 286928 561922
rect 317328 562350 317648 562384
rect 317328 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 317648 562350
rect 317328 562226 317648 562294
rect 317328 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 317648 562226
rect 317328 562102 317648 562170
rect 317328 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 317648 562102
rect 317328 561978 317648 562046
rect 317328 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 317648 561978
rect 317328 561888 317648 561922
rect 348048 562350 348368 562384
rect 348048 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 348368 562350
rect 348048 562226 348368 562294
rect 348048 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 348368 562226
rect 348048 562102 348368 562170
rect 348048 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 348368 562102
rect 348048 561978 348368 562046
rect 348048 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 348368 561978
rect 348048 561888 348368 561922
rect 378768 562350 379088 562384
rect 378768 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 379088 562350
rect 378768 562226 379088 562294
rect 378768 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 379088 562226
rect 378768 562102 379088 562170
rect 378768 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 379088 562102
rect 378768 561978 379088 562046
rect 378768 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 379088 561978
rect 378768 561888 379088 561922
rect 409488 562350 409808 562384
rect 409488 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 409808 562350
rect 409488 562226 409808 562294
rect 409488 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 409808 562226
rect 409488 562102 409808 562170
rect 409488 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 409808 562102
rect 409488 561978 409808 562046
rect 409488 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 409808 561978
rect 409488 561888 409808 561922
rect 440208 562350 440528 562384
rect 440208 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 440528 562350
rect 440208 562226 440528 562294
rect 440208 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 440528 562226
rect 440208 562102 440528 562170
rect 440208 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 440528 562102
rect 440208 561978 440528 562046
rect 440208 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 440528 561978
rect 440208 561888 440528 561922
rect 470928 562350 471248 562384
rect 470928 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 471248 562350
rect 470928 562226 471248 562294
rect 470928 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 471248 562226
rect 470928 562102 471248 562170
rect 470928 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 471248 562102
rect 470928 561978 471248 562046
rect 470928 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 471248 561978
rect 470928 561888 471248 561922
rect 209808 550350 210128 550384
rect 209808 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 210128 550350
rect 209808 550226 210128 550294
rect 209808 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 210128 550226
rect 209808 550102 210128 550170
rect 209808 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 210128 550102
rect 209808 549978 210128 550046
rect 209808 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 210128 549978
rect 209808 549888 210128 549922
rect 240528 550350 240848 550384
rect 240528 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 240848 550350
rect 240528 550226 240848 550294
rect 240528 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 240848 550226
rect 240528 550102 240848 550170
rect 240528 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 240848 550102
rect 240528 549978 240848 550046
rect 240528 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 240848 549978
rect 240528 549888 240848 549922
rect 271248 550350 271568 550384
rect 271248 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 271568 550350
rect 271248 550226 271568 550294
rect 271248 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 271568 550226
rect 271248 550102 271568 550170
rect 271248 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 271568 550102
rect 271248 549978 271568 550046
rect 271248 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 271568 549978
rect 271248 549888 271568 549922
rect 301968 550350 302288 550384
rect 301968 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 302288 550350
rect 301968 550226 302288 550294
rect 301968 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 302288 550226
rect 301968 550102 302288 550170
rect 301968 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 302288 550102
rect 301968 549978 302288 550046
rect 301968 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 302288 549978
rect 301968 549888 302288 549922
rect 332688 550350 333008 550384
rect 332688 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 333008 550350
rect 332688 550226 333008 550294
rect 332688 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 333008 550226
rect 332688 550102 333008 550170
rect 332688 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 333008 550102
rect 332688 549978 333008 550046
rect 332688 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 333008 549978
rect 332688 549888 333008 549922
rect 363408 550350 363728 550384
rect 363408 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 363728 550350
rect 363408 550226 363728 550294
rect 363408 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 363728 550226
rect 363408 550102 363728 550170
rect 363408 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 363728 550102
rect 363408 549978 363728 550046
rect 363408 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 363728 549978
rect 363408 549888 363728 549922
rect 394128 550350 394448 550384
rect 394128 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 394448 550350
rect 394128 550226 394448 550294
rect 394128 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 394448 550226
rect 394128 550102 394448 550170
rect 394128 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 394448 550102
rect 394128 549978 394448 550046
rect 394128 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 394448 549978
rect 394128 549888 394448 549922
rect 424848 550350 425168 550384
rect 424848 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 425168 550350
rect 424848 550226 425168 550294
rect 424848 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 425168 550226
rect 424848 550102 425168 550170
rect 424848 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 425168 550102
rect 424848 549978 425168 550046
rect 424848 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 425168 549978
rect 424848 549888 425168 549922
rect 455568 550350 455888 550384
rect 455568 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 455888 550350
rect 455568 550226 455888 550294
rect 455568 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 455888 550226
rect 455568 550102 455888 550170
rect 455568 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 455888 550102
rect 455568 549978 455888 550046
rect 455568 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 455888 549978
rect 455568 549888 455888 549922
rect 225168 544350 225488 544384
rect 225168 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 225488 544350
rect 225168 544226 225488 544294
rect 225168 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 225488 544226
rect 225168 544102 225488 544170
rect 225168 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 225488 544102
rect 225168 543978 225488 544046
rect 225168 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 225488 543978
rect 225168 543888 225488 543922
rect 255888 544350 256208 544384
rect 255888 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 256208 544350
rect 255888 544226 256208 544294
rect 255888 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 256208 544226
rect 255888 544102 256208 544170
rect 255888 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 256208 544102
rect 255888 543978 256208 544046
rect 255888 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 256208 543978
rect 255888 543888 256208 543922
rect 286608 544350 286928 544384
rect 286608 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 286928 544350
rect 286608 544226 286928 544294
rect 286608 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 286928 544226
rect 286608 544102 286928 544170
rect 286608 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 286928 544102
rect 286608 543978 286928 544046
rect 286608 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 286928 543978
rect 286608 543888 286928 543922
rect 317328 544350 317648 544384
rect 317328 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 317648 544350
rect 317328 544226 317648 544294
rect 317328 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 317648 544226
rect 317328 544102 317648 544170
rect 317328 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 317648 544102
rect 317328 543978 317648 544046
rect 317328 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 317648 543978
rect 317328 543888 317648 543922
rect 348048 544350 348368 544384
rect 348048 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 348368 544350
rect 348048 544226 348368 544294
rect 348048 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 348368 544226
rect 348048 544102 348368 544170
rect 348048 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 348368 544102
rect 348048 543978 348368 544046
rect 348048 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 348368 543978
rect 348048 543888 348368 543922
rect 378768 544350 379088 544384
rect 378768 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 379088 544350
rect 378768 544226 379088 544294
rect 378768 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 379088 544226
rect 378768 544102 379088 544170
rect 378768 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 379088 544102
rect 378768 543978 379088 544046
rect 378768 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 379088 543978
rect 378768 543888 379088 543922
rect 409488 544350 409808 544384
rect 409488 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 409808 544350
rect 409488 544226 409808 544294
rect 409488 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 409808 544226
rect 409488 544102 409808 544170
rect 409488 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 409808 544102
rect 409488 543978 409808 544046
rect 409488 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 409808 543978
rect 409488 543888 409808 543922
rect 440208 544350 440528 544384
rect 440208 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 440528 544350
rect 440208 544226 440528 544294
rect 440208 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 440528 544226
rect 440208 544102 440528 544170
rect 440208 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 440528 544102
rect 440208 543978 440528 544046
rect 440208 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 440528 543978
rect 440208 543888 440528 543922
rect 470928 544350 471248 544384
rect 470928 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 471248 544350
rect 470928 544226 471248 544294
rect 470928 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 471248 544226
rect 470928 544102 471248 544170
rect 470928 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 471248 544102
rect 470928 543978 471248 544046
rect 470928 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 471248 543978
rect 470928 543888 471248 543922
rect 209808 532350 210128 532384
rect 209808 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 210128 532350
rect 209808 532226 210128 532294
rect 209808 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 210128 532226
rect 209808 532102 210128 532170
rect 209808 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 210128 532102
rect 209808 531978 210128 532046
rect 209808 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 210128 531978
rect 209808 531888 210128 531922
rect 240528 532350 240848 532384
rect 240528 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 240848 532350
rect 240528 532226 240848 532294
rect 240528 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 240848 532226
rect 240528 532102 240848 532170
rect 240528 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 240848 532102
rect 240528 531978 240848 532046
rect 240528 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 240848 531978
rect 240528 531888 240848 531922
rect 271248 532350 271568 532384
rect 271248 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 271568 532350
rect 271248 532226 271568 532294
rect 271248 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 271568 532226
rect 271248 532102 271568 532170
rect 271248 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 271568 532102
rect 271248 531978 271568 532046
rect 271248 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 271568 531978
rect 271248 531888 271568 531922
rect 301968 532350 302288 532384
rect 301968 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 302288 532350
rect 301968 532226 302288 532294
rect 301968 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 302288 532226
rect 301968 532102 302288 532170
rect 301968 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 302288 532102
rect 301968 531978 302288 532046
rect 301968 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 302288 531978
rect 301968 531888 302288 531922
rect 332688 532350 333008 532384
rect 332688 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 333008 532350
rect 332688 532226 333008 532294
rect 332688 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 333008 532226
rect 332688 532102 333008 532170
rect 332688 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 333008 532102
rect 332688 531978 333008 532046
rect 332688 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 333008 531978
rect 332688 531888 333008 531922
rect 363408 532350 363728 532384
rect 363408 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 363728 532350
rect 363408 532226 363728 532294
rect 363408 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 363728 532226
rect 363408 532102 363728 532170
rect 363408 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 363728 532102
rect 363408 531978 363728 532046
rect 363408 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 363728 531978
rect 363408 531888 363728 531922
rect 394128 532350 394448 532384
rect 394128 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 394448 532350
rect 394128 532226 394448 532294
rect 394128 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 394448 532226
rect 394128 532102 394448 532170
rect 394128 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 394448 532102
rect 394128 531978 394448 532046
rect 394128 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 394448 531978
rect 394128 531888 394448 531922
rect 424848 532350 425168 532384
rect 424848 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 425168 532350
rect 424848 532226 425168 532294
rect 424848 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 425168 532226
rect 424848 532102 425168 532170
rect 424848 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 425168 532102
rect 424848 531978 425168 532046
rect 424848 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 425168 531978
rect 424848 531888 425168 531922
rect 455568 532350 455888 532384
rect 455568 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 455888 532350
rect 455568 532226 455888 532294
rect 455568 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 455888 532226
rect 455568 532102 455888 532170
rect 455568 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 455888 532102
rect 455568 531978 455888 532046
rect 455568 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 455888 531978
rect 455568 531888 455888 531922
rect 225168 526350 225488 526384
rect 225168 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 225488 526350
rect 225168 526226 225488 526294
rect 225168 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 225488 526226
rect 225168 526102 225488 526170
rect 225168 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 225488 526102
rect 225168 525978 225488 526046
rect 225168 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 225488 525978
rect 225168 525888 225488 525922
rect 255888 526350 256208 526384
rect 255888 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 256208 526350
rect 255888 526226 256208 526294
rect 255888 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 256208 526226
rect 255888 526102 256208 526170
rect 255888 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 256208 526102
rect 255888 525978 256208 526046
rect 255888 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 256208 525978
rect 255888 525888 256208 525922
rect 286608 526350 286928 526384
rect 286608 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 286928 526350
rect 286608 526226 286928 526294
rect 286608 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 286928 526226
rect 286608 526102 286928 526170
rect 286608 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 286928 526102
rect 286608 525978 286928 526046
rect 286608 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 286928 525978
rect 286608 525888 286928 525922
rect 317328 526350 317648 526384
rect 317328 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 317648 526350
rect 317328 526226 317648 526294
rect 317328 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 317648 526226
rect 317328 526102 317648 526170
rect 317328 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 317648 526102
rect 317328 525978 317648 526046
rect 317328 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 317648 525978
rect 317328 525888 317648 525922
rect 348048 526350 348368 526384
rect 348048 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 348368 526350
rect 348048 526226 348368 526294
rect 348048 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 348368 526226
rect 348048 526102 348368 526170
rect 348048 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 348368 526102
rect 348048 525978 348368 526046
rect 348048 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 348368 525978
rect 348048 525888 348368 525922
rect 378768 526350 379088 526384
rect 378768 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 379088 526350
rect 378768 526226 379088 526294
rect 378768 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 379088 526226
rect 378768 526102 379088 526170
rect 378768 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 379088 526102
rect 378768 525978 379088 526046
rect 378768 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 379088 525978
rect 378768 525888 379088 525922
rect 409488 526350 409808 526384
rect 409488 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 409808 526350
rect 409488 526226 409808 526294
rect 409488 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 409808 526226
rect 409488 526102 409808 526170
rect 409488 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 409808 526102
rect 409488 525978 409808 526046
rect 409488 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 409808 525978
rect 409488 525888 409808 525922
rect 440208 526350 440528 526384
rect 440208 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 440528 526350
rect 440208 526226 440528 526294
rect 440208 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 440528 526226
rect 440208 526102 440528 526170
rect 440208 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 440528 526102
rect 440208 525978 440528 526046
rect 440208 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 440528 525978
rect 440208 525888 440528 525922
rect 470928 526350 471248 526384
rect 470928 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 471248 526350
rect 470928 526226 471248 526294
rect 470928 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 471248 526226
rect 470928 526102 471248 526170
rect 470928 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 471248 526102
rect 470928 525978 471248 526046
rect 470928 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 471248 525978
rect 470928 525888 471248 525922
rect 209808 514350 210128 514384
rect 209808 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 210128 514350
rect 209808 514226 210128 514294
rect 209808 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 210128 514226
rect 209808 514102 210128 514170
rect 209808 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 210128 514102
rect 209808 513978 210128 514046
rect 209808 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 210128 513978
rect 209808 513888 210128 513922
rect 240528 514350 240848 514384
rect 240528 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 240848 514350
rect 240528 514226 240848 514294
rect 240528 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 240848 514226
rect 240528 514102 240848 514170
rect 240528 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 240848 514102
rect 240528 513978 240848 514046
rect 240528 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 240848 513978
rect 240528 513888 240848 513922
rect 271248 514350 271568 514384
rect 271248 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 271568 514350
rect 271248 514226 271568 514294
rect 271248 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 271568 514226
rect 271248 514102 271568 514170
rect 271248 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 271568 514102
rect 271248 513978 271568 514046
rect 271248 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 271568 513978
rect 271248 513888 271568 513922
rect 301968 514350 302288 514384
rect 301968 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 302288 514350
rect 301968 514226 302288 514294
rect 301968 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 302288 514226
rect 301968 514102 302288 514170
rect 301968 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 302288 514102
rect 301968 513978 302288 514046
rect 301968 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 302288 513978
rect 301968 513888 302288 513922
rect 332688 514350 333008 514384
rect 332688 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 333008 514350
rect 332688 514226 333008 514294
rect 332688 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 333008 514226
rect 332688 514102 333008 514170
rect 332688 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 333008 514102
rect 332688 513978 333008 514046
rect 332688 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 333008 513978
rect 332688 513888 333008 513922
rect 363408 514350 363728 514384
rect 363408 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 363728 514350
rect 363408 514226 363728 514294
rect 363408 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 363728 514226
rect 363408 514102 363728 514170
rect 363408 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 363728 514102
rect 363408 513978 363728 514046
rect 363408 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 363728 513978
rect 363408 513888 363728 513922
rect 394128 514350 394448 514384
rect 394128 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 394448 514350
rect 394128 514226 394448 514294
rect 394128 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 394448 514226
rect 394128 514102 394448 514170
rect 394128 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 394448 514102
rect 394128 513978 394448 514046
rect 394128 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 394448 513978
rect 394128 513888 394448 513922
rect 424848 514350 425168 514384
rect 424848 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 425168 514350
rect 424848 514226 425168 514294
rect 424848 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 425168 514226
rect 424848 514102 425168 514170
rect 424848 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 425168 514102
rect 424848 513978 425168 514046
rect 424848 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 425168 513978
rect 424848 513888 425168 513922
rect 455568 514350 455888 514384
rect 455568 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 455888 514350
rect 455568 514226 455888 514294
rect 455568 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 455888 514226
rect 455568 514102 455888 514170
rect 455568 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 455888 514102
rect 455568 513978 455888 514046
rect 455568 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 455888 513978
rect 455568 513888 455888 513922
rect 225168 508350 225488 508384
rect 225168 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 225488 508350
rect 225168 508226 225488 508294
rect 225168 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 225488 508226
rect 225168 508102 225488 508170
rect 225168 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 225488 508102
rect 225168 507978 225488 508046
rect 225168 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 225488 507978
rect 225168 507888 225488 507922
rect 255888 508350 256208 508384
rect 255888 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 256208 508350
rect 255888 508226 256208 508294
rect 255888 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 256208 508226
rect 255888 508102 256208 508170
rect 255888 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 256208 508102
rect 255888 507978 256208 508046
rect 255888 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 256208 507978
rect 255888 507888 256208 507922
rect 286608 508350 286928 508384
rect 286608 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 286928 508350
rect 286608 508226 286928 508294
rect 286608 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 286928 508226
rect 286608 508102 286928 508170
rect 286608 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 286928 508102
rect 286608 507978 286928 508046
rect 286608 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 286928 507978
rect 286608 507888 286928 507922
rect 317328 508350 317648 508384
rect 317328 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 317648 508350
rect 317328 508226 317648 508294
rect 317328 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 317648 508226
rect 317328 508102 317648 508170
rect 317328 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 317648 508102
rect 317328 507978 317648 508046
rect 317328 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 317648 507978
rect 317328 507888 317648 507922
rect 348048 508350 348368 508384
rect 348048 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 348368 508350
rect 348048 508226 348368 508294
rect 348048 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 348368 508226
rect 348048 508102 348368 508170
rect 348048 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 348368 508102
rect 348048 507978 348368 508046
rect 348048 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 348368 507978
rect 348048 507888 348368 507922
rect 378768 508350 379088 508384
rect 378768 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 379088 508350
rect 378768 508226 379088 508294
rect 378768 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 379088 508226
rect 378768 508102 379088 508170
rect 378768 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 379088 508102
rect 378768 507978 379088 508046
rect 378768 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 379088 507978
rect 378768 507888 379088 507922
rect 409488 508350 409808 508384
rect 409488 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 409808 508350
rect 409488 508226 409808 508294
rect 409488 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 409808 508226
rect 409488 508102 409808 508170
rect 409488 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 409808 508102
rect 409488 507978 409808 508046
rect 409488 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 409808 507978
rect 409488 507888 409808 507922
rect 440208 508350 440528 508384
rect 440208 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 440528 508350
rect 440208 508226 440528 508294
rect 440208 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 440528 508226
rect 440208 508102 440528 508170
rect 440208 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 440528 508102
rect 440208 507978 440528 508046
rect 440208 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 440528 507978
rect 440208 507888 440528 507922
rect 470928 508350 471248 508384
rect 470928 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 471248 508350
rect 470928 508226 471248 508294
rect 470928 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 471248 508226
rect 470928 508102 471248 508170
rect 470928 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 471248 508102
rect 470928 507978 471248 508046
rect 470928 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 471248 507978
rect 470928 507888 471248 507922
rect 209808 496350 210128 496384
rect 209808 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 210128 496350
rect 209808 496226 210128 496294
rect 209808 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 210128 496226
rect 209808 496102 210128 496170
rect 209808 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 210128 496102
rect 209808 495978 210128 496046
rect 209808 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 210128 495978
rect 209808 495888 210128 495922
rect 240528 496350 240848 496384
rect 240528 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 240848 496350
rect 240528 496226 240848 496294
rect 240528 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 240848 496226
rect 240528 496102 240848 496170
rect 240528 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 240848 496102
rect 240528 495978 240848 496046
rect 240528 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 240848 495978
rect 240528 495888 240848 495922
rect 271248 496350 271568 496384
rect 271248 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 271568 496350
rect 271248 496226 271568 496294
rect 271248 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 271568 496226
rect 271248 496102 271568 496170
rect 271248 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 271568 496102
rect 271248 495978 271568 496046
rect 271248 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 271568 495978
rect 271248 495888 271568 495922
rect 301968 496350 302288 496384
rect 301968 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 302288 496350
rect 301968 496226 302288 496294
rect 301968 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 302288 496226
rect 301968 496102 302288 496170
rect 301968 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 302288 496102
rect 301968 495978 302288 496046
rect 301968 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 302288 495978
rect 301968 495888 302288 495922
rect 332688 496350 333008 496384
rect 332688 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 333008 496350
rect 332688 496226 333008 496294
rect 332688 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 333008 496226
rect 332688 496102 333008 496170
rect 332688 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 333008 496102
rect 332688 495978 333008 496046
rect 332688 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 333008 495978
rect 332688 495888 333008 495922
rect 363408 496350 363728 496384
rect 363408 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 363728 496350
rect 363408 496226 363728 496294
rect 363408 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 363728 496226
rect 363408 496102 363728 496170
rect 363408 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 363728 496102
rect 363408 495978 363728 496046
rect 363408 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 363728 495978
rect 363408 495888 363728 495922
rect 394128 496350 394448 496384
rect 394128 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 394448 496350
rect 394128 496226 394448 496294
rect 394128 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 394448 496226
rect 394128 496102 394448 496170
rect 394128 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 394448 496102
rect 394128 495978 394448 496046
rect 394128 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 394448 495978
rect 394128 495888 394448 495922
rect 424848 496350 425168 496384
rect 424848 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 425168 496350
rect 424848 496226 425168 496294
rect 424848 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 425168 496226
rect 424848 496102 425168 496170
rect 424848 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 425168 496102
rect 424848 495978 425168 496046
rect 424848 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 425168 495978
rect 424848 495888 425168 495922
rect 455568 496350 455888 496384
rect 455568 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 455888 496350
rect 455568 496226 455888 496294
rect 455568 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 455888 496226
rect 455568 496102 455888 496170
rect 455568 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 455888 496102
rect 455568 495978 455888 496046
rect 455568 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 455888 495978
rect 455568 495888 455888 495922
rect 225168 490350 225488 490384
rect 225168 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 225488 490350
rect 225168 490226 225488 490294
rect 225168 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 225488 490226
rect 225168 490102 225488 490170
rect 225168 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 225488 490102
rect 225168 489978 225488 490046
rect 225168 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 225488 489978
rect 225168 489888 225488 489922
rect 255888 490350 256208 490384
rect 255888 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 256208 490350
rect 255888 490226 256208 490294
rect 255888 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 256208 490226
rect 255888 490102 256208 490170
rect 255888 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 256208 490102
rect 255888 489978 256208 490046
rect 255888 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 256208 489978
rect 255888 489888 256208 489922
rect 286608 490350 286928 490384
rect 286608 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 286928 490350
rect 286608 490226 286928 490294
rect 286608 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 286928 490226
rect 286608 490102 286928 490170
rect 286608 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 286928 490102
rect 286608 489978 286928 490046
rect 286608 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 286928 489978
rect 286608 489888 286928 489922
rect 317328 490350 317648 490384
rect 317328 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 317648 490350
rect 317328 490226 317648 490294
rect 317328 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 317648 490226
rect 317328 490102 317648 490170
rect 317328 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 317648 490102
rect 317328 489978 317648 490046
rect 317328 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 317648 489978
rect 317328 489888 317648 489922
rect 348048 490350 348368 490384
rect 348048 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 348368 490350
rect 348048 490226 348368 490294
rect 348048 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 348368 490226
rect 348048 490102 348368 490170
rect 348048 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 348368 490102
rect 348048 489978 348368 490046
rect 348048 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 348368 489978
rect 348048 489888 348368 489922
rect 378768 490350 379088 490384
rect 378768 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 379088 490350
rect 378768 490226 379088 490294
rect 378768 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 379088 490226
rect 378768 490102 379088 490170
rect 378768 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 379088 490102
rect 378768 489978 379088 490046
rect 378768 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 379088 489978
rect 378768 489888 379088 489922
rect 409488 490350 409808 490384
rect 409488 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 409808 490350
rect 409488 490226 409808 490294
rect 409488 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 409808 490226
rect 409488 490102 409808 490170
rect 409488 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 409808 490102
rect 409488 489978 409808 490046
rect 409488 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 409808 489978
rect 409488 489888 409808 489922
rect 440208 490350 440528 490384
rect 440208 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 440528 490350
rect 440208 490226 440528 490294
rect 440208 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 440528 490226
rect 440208 490102 440528 490170
rect 440208 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 440528 490102
rect 440208 489978 440528 490046
rect 440208 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 440528 489978
rect 440208 489888 440528 489922
rect 470928 490350 471248 490384
rect 470928 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 471248 490350
rect 470928 490226 471248 490294
rect 470928 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 471248 490226
rect 470928 490102 471248 490170
rect 470928 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 471248 490102
rect 470928 489978 471248 490046
rect 470928 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 471248 489978
rect 470928 489888 471248 489922
rect 209808 478350 210128 478384
rect 209808 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 210128 478350
rect 209808 478226 210128 478294
rect 209808 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 210128 478226
rect 209808 478102 210128 478170
rect 209808 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 210128 478102
rect 209808 477978 210128 478046
rect 209808 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 210128 477978
rect 209808 477888 210128 477922
rect 240528 478350 240848 478384
rect 240528 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 240848 478350
rect 240528 478226 240848 478294
rect 240528 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 240848 478226
rect 240528 478102 240848 478170
rect 240528 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 240848 478102
rect 240528 477978 240848 478046
rect 240528 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 240848 477978
rect 240528 477888 240848 477922
rect 271248 478350 271568 478384
rect 271248 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 271568 478350
rect 271248 478226 271568 478294
rect 271248 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 271568 478226
rect 271248 478102 271568 478170
rect 271248 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 271568 478102
rect 271248 477978 271568 478046
rect 271248 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 271568 477978
rect 271248 477888 271568 477922
rect 301968 478350 302288 478384
rect 301968 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 302288 478350
rect 301968 478226 302288 478294
rect 301968 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 302288 478226
rect 301968 478102 302288 478170
rect 301968 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 302288 478102
rect 301968 477978 302288 478046
rect 301968 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 302288 477978
rect 301968 477888 302288 477922
rect 332688 478350 333008 478384
rect 332688 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 333008 478350
rect 332688 478226 333008 478294
rect 332688 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 333008 478226
rect 332688 478102 333008 478170
rect 332688 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 333008 478102
rect 332688 477978 333008 478046
rect 332688 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 333008 477978
rect 332688 477888 333008 477922
rect 363408 478350 363728 478384
rect 363408 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 363728 478350
rect 363408 478226 363728 478294
rect 363408 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 363728 478226
rect 363408 478102 363728 478170
rect 363408 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 363728 478102
rect 363408 477978 363728 478046
rect 363408 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 363728 477978
rect 363408 477888 363728 477922
rect 394128 478350 394448 478384
rect 394128 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 394448 478350
rect 394128 478226 394448 478294
rect 394128 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 394448 478226
rect 394128 478102 394448 478170
rect 394128 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 394448 478102
rect 394128 477978 394448 478046
rect 394128 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 394448 477978
rect 394128 477888 394448 477922
rect 424848 478350 425168 478384
rect 424848 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 425168 478350
rect 424848 478226 425168 478294
rect 424848 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 425168 478226
rect 424848 478102 425168 478170
rect 424848 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 425168 478102
rect 424848 477978 425168 478046
rect 424848 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 425168 477978
rect 424848 477888 425168 477922
rect 455568 478350 455888 478384
rect 455568 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 455888 478350
rect 455568 478226 455888 478294
rect 455568 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 455888 478226
rect 455568 478102 455888 478170
rect 455568 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 455888 478102
rect 455568 477978 455888 478046
rect 455568 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 455888 477978
rect 455568 477888 455888 477922
rect 225168 472350 225488 472384
rect 225168 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 225488 472350
rect 225168 472226 225488 472294
rect 225168 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 225488 472226
rect 225168 472102 225488 472170
rect 225168 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 225488 472102
rect 225168 471978 225488 472046
rect 225168 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 225488 471978
rect 225168 471888 225488 471922
rect 255888 472350 256208 472384
rect 255888 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 256208 472350
rect 255888 472226 256208 472294
rect 255888 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 256208 472226
rect 255888 472102 256208 472170
rect 255888 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 256208 472102
rect 255888 471978 256208 472046
rect 255888 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 256208 471978
rect 255888 471888 256208 471922
rect 286608 472350 286928 472384
rect 286608 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 286928 472350
rect 286608 472226 286928 472294
rect 286608 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 286928 472226
rect 286608 472102 286928 472170
rect 286608 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 286928 472102
rect 286608 471978 286928 472046
rect 286608 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 286928 471978
rect 286608 471888 286928 471922
rect 317328 472350 317648 472384
rect 317328 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 317648 472350
rect 317328 472226 317648 472294
rect 317328 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 317648 472226
rect 317328 472102 317648 472170
rect 317328 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 317648 472102
rect 317328 471978 317648 472046
rect 317328 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 317648 471978
rect 317328 471888 317648 471922
rect 348048 472350 348368 472384
rect 348048 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 348368 472350
rect 348048 472226 348368 472294
rect 348048 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 348368 472226
rect 348048 472102 348368 472170
rect 348048 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 348368 472102
rect 348048 471978 348368 472046
rect 348048 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 348368 471978
rect 348048 471888 348368 471922
rect 378768 472350 379088 472384
rect 378768 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 379088 472350
rect 378768 472226 379088 472294
rect 378768 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 379088 472226
rect 378768 472102 379088 472170
rect 378768 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 379088 472102
rect 378768 471978 379088 472046
rect 378768 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 379088 471978
rect 378768 471888 379088 471922
rect 409488 472350 409808 472384
rect 409488 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 409808 472350
rect 409488 472226 409808 472294
rect 409488 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 409808 472226
rect 409488 472102 409808 472170
rect 409488 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 409808 472102
rect 409488 471978 409808 472046
rect 409488 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 409808 471978
rect 409488 471888 409808 471922
rect 440208 472350 440528 472384
rect 440208 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 440528 472350
rect 440208 472226 440528 472294
rect 440208 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 440528 472226
rect 440208 472102 440528 472170
rect 440208 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 440528 472102
rect 440208 471978 440528 472046
rect 440208 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 440528 471978
rect 440208 471888 440528 471922
rect 470928 472350 471248 472384
rect 470928 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 471248 472350
rect 470928 472226 471248 472294
rect 470928 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 471248 472226
rect 470928 472102 471248 472170
rect 470928 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 471248 472102
rect 470928 471978 471248 472046
rect 470928 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 471248 471978
rect 470928 471888 471248 471922
rect 209808 460350 210128 460384
rect 209808 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 210128 460350
rect 209808 460226 210128 460294
rect 209808 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 210128 460226
rect 209808 460102 210128 460170
rect 209808 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 210128 460102
rect 209808 459978 210128 460046
rect 209808 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 210128 459978
rect 209808 459888 210128 459922
rect 240528 460350 240848 460384
rect 240528 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 240848 460350
rect 240528 460226 240848 460294
rect 240528 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 240848 460226
rect 240528 460102 240848 460170
rect 240528 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 240848 460102
rect 240528 459978 240848 460046
rect 240528 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 240848 459978
rect 240528 459888 240848 459922
rect 271248 460350 271568 460384
rect 271248 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 271568 460350
rect 271248 460226 271568 460294
rect 271248 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 271568 460226
rect 271248 460102 271568 460170
rect 271248 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 271568 460102
rect 271248 459978 271568 460046
rect 271248 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 271568 459978
rect 271248 459888 271568 459922
rect 301968 460350 302288 460384
rect 301968 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 302288 460350
rect 301968 460226 302288 460294
rect 301968 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 302288 460226
rect 301968 460102 302288 460170
rect 301968 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 302288 460102
rect 301968 459978 302288 460046
rect 301968 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 302288 459978
rect 301968 459888 302288 459922
rect 332688 460350 333008 460384
rect 332688 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 333008 460350
rect 332688 460226 333008 460294
rect 332688 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 333008 460226
rect 332688 460102 333008 460170
rect 332688 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 333008 460102
rect 332688 459978 333008 460046
rect 332688 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 333008 459978
rect 332688 459888 333008 459922
rect 363408 460350 363728 460384
rect 363408 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 363728 460350
rect 363408 460226 363728 460294
rect 363408 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 363728 460226
rect 363408 460102 363728 460170
rect 363408 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 363728 460102
rect 363408 459978 363728 460046
rect 363408 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 363728 459978
rect 363408 459888 363728 459922
rect 394128 460350 394448 460384
rect 394128 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 394448 460350
rect 394128 460226 394448 460294
rect 394128 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 394448 460226
rect 394128 460102 394448 460170
rect 394128 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 394448 460102
rect 394128 459978 394448 460046
rect 394128 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 394448 459978
rect 394128 459888 394448 459922
rect 424848 460350 425168 460384
rect 424848 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 425168 460350
rect 424848 460226 425168 460294
rect 424848 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 425168 460226
rect 424848 460102 425168 460170
rect 424848 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 425168 460102
rect 424848 459978 425168 460046
rect 424848 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 425168 459978
rect 424848 459888 425168 459922
rect 455568 460350 455888 460384
rect 455568 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 455888 460350
rect 455568 460226 455888 460294
rect 455568 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 455888 460226
rect 455568 460102 455888 460170
rect 455568 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 455888 460102
rect 455568 459978 455888 460046
rect 455568 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 455888 459978
rect 455568 459888 455888 459922
rect 225168 454350 225488 454384
rect 225168 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 225488 454350
rect 225168 454226 225488 454294
rect 225168 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 225488 454226
rect 225168 454102 225488 454170
rect 225168 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 225488 454102
rect 225168 453978 225488 454046
rect 225168 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 225488 453978
rect 225168 453888 225488 453922
rect 255888 454350 256208 454384
rect 255888 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 256208 454350
rect 255888 454226 256208 454294
rect 255888 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 256208 454226
rect 255888 454102 256208 454170
rect 255888 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 256208 454102
rect 255888 453978 256208 454046
rect 255888 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 256208 453978
rect 255888 453888 256208 453922
rect 286608 454350 286928 454384
rect 286608 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 286928 454350
rect 286608 454226 286928 454294
rect 286608 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 286928 454226
rect 286608 454102 286928 454170
rect 286608 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 286928 454102
rect 286608 453978 286928 454046
rect 286608 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 286928 453978
rect 286608 453888 286928 453922
rect 317328 454350 317648 454384
rect 317328 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 317648 454350
rect 317328 454226 317648 454294
rect 317328 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 317648 454226
rect 317328 454102 317648 454170
rect 317328 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 317648 454102
rect 317328 453978 317648 454046
rect 317328 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 317648 453978
rect 317328 453888 317648 453922
rect 348048 454350 348368 454384
rect 348048 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 348368 454350
rect 348048 454226 348368 454294
rect 348048 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 348368 454226
rect 348048 454102 348368 454170
rect 348048 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 348368 454102
rect 348048 453978 348368 454046
rect 348048 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 348368 453978
rect 348048 453888 348368 453922
rect 378768 454350 379088 454384
rect 378768 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 379088 454350
rect 378768 454226 379088 454294
rect 378768 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 379088 454226
rect 378768 454102 379088 454170
rect 378768 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 379088 454102
rect 378768 453978 379088 454046
rect 378768 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 379088 453978
rect 378768 453888 379088 453922
rect 409488 454350 409808 454384
rect 409488 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 409808 454350
rect 409488 454226 409808 454294
rect 409488 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 409808 454226
rect 409488 454102 409808 454170
rect 409488 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 409808 454102
rect 409488 453978 409808 454046
rect 409488 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 409808 453978
rect 409488 453888 409808 453922
rect 440208 454350 440528 454384
rect 440208 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 440528 454350
rect 440208 454226 440528 454294
rect 440208 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 440528 454226
rect 440208 454102 440528 454170
rect 440208 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 440528 454102
rect 440208 453978 440528 454046
rect 440208 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 440528 453978
rect 440208 453888 440528 453922
rect 470928 454350 471248 454384
rect 470928 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 471248 454350
rect 470928 454226 471248 454294
rect 470928 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 471248 454226
rect 470928 454102 471248 454170
rect 470928 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 471248 454102
rect 470928 453978 471248 454046
rect 470928 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 471248 453978
rect 470928 453888 471248 453922
rect 209808 442350 210128 442384
rect 209808 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 210128 442350
rect 209808 442226 210128 442294
rect 209808 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 210128 442226
rect 209808 442102 210128 442170
rect 209808 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 210128 442102
rect 209808 441978 210128 442046
rect 209808 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 210128 441978
rect 209808 441888 210128 441922
rect 240528 442350 240848 442384
rect 240528 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 240848 442350
rect 240528 442226 240848 442294
rect 240528 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 240848 442226
rect 240528 442102 240848 442170
rect 240528 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 240848 442102
rect 240528 441978 240848 442046
rect 240528 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 240848 441978
rect 240528 441888 240848 441922
rect 271248 442350 271568 442384
rect 271248 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 271568 442350
rect 271248 442226 271568 442294
rect 271248 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 271568 442226
rect 271248 442102 271568 442170
rect 271248 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 271568 442102
rect 271248 441978 271568 442046
rect 271248 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 271568 441978
rect 271248 441888 271568 441922
rect 301968 442350 302288 442384
rect 301968 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 302288 442350
rect 301968 442226 302288 442294
rect 301968 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 302288 442226
rect 301968 442102 302288 442170
rect 301968 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 302288 442102
rect 301968 441978 302288 442046
rect 301968 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 302288 441978
rect 301968 441888 302288 441922
rect 332688 442350 333008 442384
rect 332688 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 333008 442350
rect 332688 442226 333008 442294
rect 332688 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 333008 442226
rect 332688 442102 333008 442170
rect 332688 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 333008 442102
rect 332688 441978 333008 442046
rect 332688 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 333008 441978
rect 332688 441888 333008 441922
rect 363408 442350 363728 442384
rect 363408 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 363728 442350
rect 363408 442226 363728 442294
rect 363408 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 363728 442226
rect 363408 442102 363728 442170
rect 363408 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 363728 442102
rect 363408 441978 363728 442046
rect 363408 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 363728 441978
rect 363408 441888 363728 441922
rect 394128 442350 394448 442384
rect 394128 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 394448 442350
rect 394128 442226 394448 442294
rect 394128 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 394448 442226
rect 394128 442102 394448 442170
rect 394128 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 394448 442102
rect 394128 441978 394448 442046
rect 394128 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 394448 441978
rect 394128 441888 394448 441922
rect 424848 442350 425168 442384
rect 424848 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 425168 442350
rect 424848 442226 425168 442294
rect 424848 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 425168 442226
rect 424848 442102 425168 442170
rect 424848 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 425168 442102
rect 424848 441978 425168 442046
rect 424848 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 425168 441978
rect 424848 441888 425168 441922
rect 455568 442350 455888 442384
rect 455568 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 455888 442350
rect 455568 442226 455888 442294
rect 455568 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 455888 442226
rect 455568 442102 455888 442170
rect 455568 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 455888 442102
rect 455568 441978 455888 442046
rect 455568 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 455888 441978
rect 455568 441888 455888 441922
rect 225168 436350 225488 436384
rect 225168 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 225488 436350
rect 225168 436226 225488 436294
rect 225168 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 225488 436226
rect 225168 436102 225488 436170
rect 225168 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 225488 436102
rect 225168 435978 225488 436046
rect 225168 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 225488 435978
rect 225168 435888 225488 435922
rect 255888 436350 256208 436384
rect 255888 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 256208 436350
rect 255888 436226 256208 436294
rect 255888 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 256208 436226
rect 255888 436102 256208 436170
rect 255888 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 256208 436102
rect 255888 435978 256208 436046
rect 255888 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 256208 435978
rect 255888 435888 256208 435922
rect 286608 436350 286928 436384
rect 286608 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 286928 436350
rect 286608 436226 286928 436294
rect 286608 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 286928 436226
rect 286608 436102 286928 436170
rect 286608 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 286928 436102
rect 286608 435978 286928 436046
rect 286608 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 286928 435978
rect 286608 435888 286928 435922
rect 317328 436350 317648 436384
rect 317328 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 317648 436350
rect 317328 436226 317648 436294
rect 317328 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 317648 436226
rect 317328 436102 317648 436170
rect 317328 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 317648 436102
rect 317328 435978 317648 436046
rect 317328 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 317648 435978
rect 317328 435888 317648 435922
rect 348048 436350 348368 436384
rect 348048 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 348368 436350
rect 348048 436226 348368 436294
rect 348048 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 348368 436226
rect 348048 436102 348368 436170
rect 348048 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 348368 436102
rect 348048 435978 348368 436046
rect 348048 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 348368 435978
rect 348048 435888 348368 435922
rect 378768 436350 379088 436384
rect 378768 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 379088 436350
rect 378768 436226 379088 436294
rect 378768 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 379088 436226
rect 378768 436102 379088 436170
rect 378768 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 379088 436102
rect 378768 435978 379088 436046
rect 378768 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 379088 435978
rect 378768 435888 379088 435922
rect 409488 436350 409808 436384
rect 409488 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 409808 436350
rect 409488 436226 409808 436294
rect 409488 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 409808 436226
rect 409488 436102 409808 436170
rect 409488 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 409808 436102
rect 409488 435978 409808 436046
rect 409488 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 409808 435978
rect 409488 435888 409808 435922
rect 440208 436350 440528 436384
rect 440208 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 440528 436350
rect 440208 436226 440528 436294
rect 440208 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 440528 436226
rect 440208 436102 440528 436170
rect 440208 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 440528 436102
rect 440208 435978 440528 436046
rect 440208 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 440528 435978
rect 440208 435888 440528 435922
rect 470928 436350 471248 436384
rect 470928 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 471248 436350
rect 470928 436226 471248 436294
rect 470928 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 471248 436226
rect 470928 436102 471248 436170
rect 470928 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 471248 436102
rect 470928 435978 471248 436046
rect 470928 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 471248 435978
rect 470928 435888 471248 435922
rect 209808 424350 210128 424384
rect 209808 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 210128 424350
rect 209808 424226 210128 424294
rect 209808 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 210128 424226
rect 209808 424102 210128 424170
rect 209808 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 210128 424102
rect 209808 423978 210128 424046
rect 209808 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 210128 423978
rect 209808 423888 210128 423922
rect 240528 424350 240848 424384
rect 240528 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 240848 424350
rect 240528 424226 240848 424294
rect 240528 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 240848 424226
rect 240528 424102 240848 424170
rect 240528 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 240848 424102
rect 240528 423978 240848 424046
rect 240528 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 240848 423978
rect 240528 423888 240848 423922
rect 271248 424350 271568 424384
rect 271248 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 271568 424350
rect 271248 424226 271568 424294
rect 271248 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 271568 424226
rect 271248 424102 271568 424170
rect 271248 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 271568 424102
rect 271248 423978 271568 424046
rect 271248 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 271568 423978
rect 271248 423888 271568 423922
rect 301968 424350 302288 424384
rect 301968 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 302288 424350
rect 301968 424226 302288 424294
rect 301968 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 302288 424226
rect 301968 424102 302288 424170
rect 301968 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 302288 424102
rect 301968 423978 302288 424046
rect 301968 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 302288 423978
rect 301968 423888 302288 423922
rect 332688 424350 333008 424384
rect 332688 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 333008 424350
rect 332688 424226 333008 424294
rect 332688 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 333008 424226
rect 332688 424102 333008 424170
rect 332688 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 333008 424102
rect 332688 423978 333008 424046
rect 332688 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 333008 423978
rect 332688 423888 333008 423922
rect 363408 424350 363728 424384
rect 363408 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 363728 424350
rect 363408 424226 363728 424294
rect 363408 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 363728 424226
rect 363408 424102 363728 424170
rect 363408 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 363728 424102
rect 363408 423978 363728 424046
rect 363408 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 363728 423978
rect 363408 423888 363728 423922
rect 394128 424350 394448 424384
rect 394128 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 394448 424350
rect 394128 424226 394448 424294
rect 394128 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 394448 424226
rect 394128 424102 394448 424170
rect 394128 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 394448 424102
rect 394128 423978 394448 424046
rect 394128 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 394448 423978
rect 394128 423888 394448 423922
rect 424848 424350 425168 424384
rect 424848 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 425168 424350
rect 424848 424226 425168 424294
rect 424848 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 425168 424226
rect 424848 424102 425168 424170
rect 424848 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 425168 424102
rect 424848 423978 425168 424046
rect 424848 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 425168 423978
rect 424848 423888 425168 423922
rect 455568 424350 455888 424384
rect 455568 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 455888 424350
rect 455568 424226 455888 424294
rect 455568 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 455888 424226
rect 455568 424102 455888 424170
rect 455568 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 455888 424102
rect 455568 423978 455888 424046
rect 455568 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 455888 423978
rect 455568 423888 455888 423922
rect 225168 418350 225488 418384
rect 225168 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 225488 418350
rect 225168 418226 225488 418294
rect 225168 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 225488 418226
rect 225168 418102 225488 418170
rect 225168 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 225488 418102
rect 225168 417978 225488 418046
rect 225168 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 225488 417978
rect 225168 417888 225488 417922
rect 255888 418350 256208 418384
rect 255888 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 256208 418350
rect 255888 418226 256208 418294
rect 255888 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 256208 418226
rect 255888 418102 256208 418170
rect 255888 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 256208 418102
rect 255888 417978 256208 418046
rect 255888 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 256208 417978
rect 255888 417888 256208 417922
rect 286608 418350 286928 418384
rect 286608 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 286928 418350
rect 286608 418226 286928 418294
rect 286608 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 286928 418226
rect 286608 418102 286928 418170
rect 286608 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 286928 418102
rect 286608 417978 286928 418046
rect 286608 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 286928 417978
rect 286608 417888 286928 417922
rect 317328 418350 317648 418384
rect 317328 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 317648 418350
rect 317328 418226 317648 418294
rect 317328 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 317648 418226
rect 317328 418102 317648 418170
rect 317328 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 317648 418102
rect 317328 417978 317648 418046
rect 317328 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 317648 417978
rect 317328 417888 317648 417922
rect 348048 418350 348368 418384
rect 348048 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 348368 418350
rect 348048 418226 348368 418294
rect 348048 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 348368 418226
rect 348048 418102 348368 418170
rect 348048 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 348368 418102
rect 348048 417978 348368 418046
rect 348048 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 348368 417978
rect 348048 417888 348368 417922
rect 378768 418350 379088 418384
rect 378768 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 379088 418350
rect 378768 418226 379088 418294
rect 378768 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 379088 418226
rect 378768 418102 379088 418170
rect 378768 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 379088 418102
rect 378768 417978 379088 418046
rect 378768 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 379088 417978
rect 378768 417888 379088 417922
rect 409488 418350 409808 418384
rect 409488 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 409808 418350
rect 409488 418226 409808 418294
rect 409488 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 409808 418226
rect 409488 418102 409808 418170
rect 409488 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 409808 418102
rect 409488 417978 409808 418046
rect 409488 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 409808 417978
rect 409488 417888 409808 417922
rect 440208 418350 440528 418384
rect 440208 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 440528 418350
rect 440208 418226 440528 418294
rect 440208 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 440528 418226
rect 440208 418102 440528 418170
rect 440208 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 440528 418102
rect 440208 417978 440528 418046
rect 440208 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 440528 417978
rect 440208 417888 440528 417922
rect 470928 418350 471248 418384
rect 470928 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 471248 418350
rect 470928 418226 471248 418294
rect 470928 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 471248 418226
rect 470928 418102 471248 418170
rect 470928 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 471248 418102
rect 470928 417978 471248 418046
rect 470928 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 471248 417978
rect 470928 417888 471248 417922
rect 336924 410518 336980 410528
rect 297276 410338 297332 410348
rect 261996 409618 262052 409628
rect 240268 409332 240324 409342
rect 206668 404038 206724 404048
rect 203532 397506 203588 397516
rect 204764 398132 204820 398142
rect 203308 390472 203364 390482
rect 204540 386820 204596 386830
rect 204428 385252 204484 385262
rect 202972 236338 203028 236348
rect 203084 383518 203140 383528
rect 202860 226482 202916 226492
rect 202636 214946 202692 214956
rect 201404 214072 201460 214082
rect 199276 212594 199332 212604
rect 196476 206512 196532 206522
rect 203084 205858 203140 383462
rect 204092 382228 204148 382238
rect 204092 302518 204148 382172
rect 203308 236068 203364 236078
rect 203308 235732 203364 236012
rect 204092 235956 204148 302462
rect 204316 378756 204372 378766
rect 204316 239428 204372 378700
rect 204428 239988 204484 385196
rect 204428 239922 204484 239932
rect 204316 239362 204372 239372
rect 204540 236068 204596 386764
rect 204540 236002 204596 236012
rect 204652 379378 204708 379388
rect 204092 235890 204148 235900
rect 203308 235666 203364 235676
rect 204652 226436 204708 379322
rect 204764 238420 204820 398076
rect 206668 383012 206724 403982
rect 208348 402418 208404 402428
rect 208348 384244 208404 402362
rect 208348 384178 208404 384188
rect 220458 400350 221078 409194
rect 220458 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 221078 400350
rect 220458 400226 221078 400294
rect 220458 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 221078 400226
rect 220458 400102 221078 400170
rect 220458 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 221078 400102
rect 220458 399978 221078 400046
rect 220458 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 221078 399978
rect 206668 382946 206724 382956
rect 214508 383338 214564 383348
rect 214508 381444 214564 383282
rect 214508 381378 214564 381388
rect 216524 383158 216580 383168
rect 216524 381444 216580 383102
rect 216524 381378 216580 381388
rect 220458 382350 221078 399922
rect 220458 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 221078 382350
rect 220458 382226 221078 382294
rect 220458 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 221078 382226
rect 220458 382102 221078 382170
rect 220458 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 221078 382102
rect 220458 381978 221078 382046
rect 220458 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 221078 381978
rect 209132 380548 209188 380558
rect 209132 380100 209188 380492
rect 209132 380034 209188 380044
rect 215852 380278 215908 380288
rect 215852 379988 215908 380222
rect 204764 238354 204820 238364
rect 204876 379918 204932 379928
rect 215852 379922 215908 379932
rect 204652 226370 204708 226380
rect 204876 220052 204932 379862
rect 218540 379918 218596 379928
rect 218540 379652 218596 379862
rect 218540 379586 218596 379596
rect 217196 379378 217252 379388
rect 213164 379316 213220 379326
rect 213164 379198 213220 379260
rect 213164 379132 213220 379142
rect 213836 379316 213892 379326
rect 213836 378838 213892 379260
rect 215180 379316 215236 379326
rect 215180 379018 215236 379260
rect 217196 379316 217252 379322
rect 217196 379250 217252 379260
rect 220458 379126 221078 381922
rect 224178 406350 224798 409194
rect 240268 407458 240324 409276
rect 240268 407392 240324 407402
rect 243516 409078 243572 409088
rect 232316 407316 232372 407326
rect 232316 406738 232372 407260
rect 232316 406672 232372 406682
rect 224178 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 224798 406350
rect 224178 406226 224798 406294
rect 224178 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 224798 406226
rect 224178 406102 224798 406170
rect 224178 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 224798 406102
rect 224178 405978 224798 406046
rect 224178 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 224798 405978
rect 224178 388350 224798 405922
rect 224178 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 224798 388350
rect 224178 388226 224798 388294
rect 224178 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 224798 388226
rect 224178 388102 224798 388170
rect 224178 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 224798 388102
rect 224178 387978 224798 388046
rect 224178 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 224798 387978
rect 224178 379126 224798 387922
rect 237692 383012 237748 383022
rect 237692 382116 237748 382956
rect 237692 382050 237748 382060
rect 243516 382004 243572 409022
rect 246876 407278 246932 407288
rect 246876 406532 246932 407222
rect 246876 406466 246932 406476
rect 243516 381938 243572 381948
rect 251178 400350 251798 409194
rect 251178 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 251798 400350
rect 251178 400226 251798 400294
rect 251178 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 251798 400226
rect 251178 400102 251798 400170
rect 251178 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 251798 400102
rect 251178 399978 251798 400046
rect 251178 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 251798 399978
rect 251178 382350 251798 399922
rect 251178 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 251798 382350
rect 251178 382226 251798 382294
rect 251178 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 251798 382226
rect 251178 382102 251798 382170
rect 251178 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 251798 382102
rect 251178 381978 251798 382046
rect 251178 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 251798 381978
rect 251178 379126 251798 381922
rect 254898 406350 255518 409194
rect 254898 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 255518 406350
rect 254898 406226 255518 406294
rect 254898 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 255518 406226
rect 254898 406102 255518 406170
rect 254898 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 255518 406102
rect 254898 405978 255518 406046
rect 254898 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 255518 405978
rect 254898 388350 255518 405922
rect 254898 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 255518 388350
rect 254898 388226 255518 388294
rect 254898 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 255518 388226
rect 254898 388102 255518 388170
rect 254898 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 255518 388102
rect 254898 387978 255518 388046
rect 254898 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 255518 387978
rect 254898 379126 255518 387922
rect 261996 381668 262052 409562
rect 278908 409438 278964 409448
rect 278908 407876 278964 409382
rect 288092 409258 288148 409268
rect 278908 407810 278964 407820
rect 278796 402418 278852 402428
rect 263676 400618 263732 400628
rect 263676 382004 263732 400562
rect 263676 381938 263732 381948
rect 278796 382004 278852 402362
rect 278796 381938 278852 381948
rect 281898 400350 282518 409194
rect 281898 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 282518 400350
rect 281898 400226 282518 400294
rect 281898 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 282518 400226
rect 281898 400102 282518 400170
rect 281898 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 282518 400102
rect 281898 399978 282518 400046
rect 281898 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 282518 399978
rect 281898 382350 282518 399922
rect 281898 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 282518 382350
rect 281898 382226 282518 382294
rect 281898 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 282518 382226
rect 281898 382102 282518 382170
rect 281898 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 282518 382102
rect 281898 381978 282518 382046
rect 261996 381602 262052 381612
rect 281898 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 282518 381978
rect 281898 379126 282518 381922
rect 285618 406350 286238 409194
rect 288092 408100 288148 409202
rect 288092 408034 288148 408044
rect 295596 408718 295652 408728
rect 285618 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 286238 406350
rect 285618 406226 286238 406294
rect 285618 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 286238 406226
rect 285618 406102 286238 406170
rect 285618 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 286238 406102
rect 285618 405978 286238 406046
rect 285618 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 286238 405978
rect 285618 388350 286238 405922
rect 285618 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 286238 388350
rect 285618 388226 286238 388294
rect 285618 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 286238 388226
rect 285618 388102 286238 388170
rect 285618 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 286238 388102
rect 285618 387978 286238 388046
rect 285618 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 286238 387978
rect 285618 379126 286238 387922
rect 293916 402778 293972 402788
rect 293916 381444 293972 402722
rect 295596 381668 295652 408662
rect 297276 382004 297332 410282
rect 297276 381938 297332 381948
rect 298956 408358 299012 408368
rect 298956 382004 299012 408302
rect 305676 407638 305732 407648
rect 302316 407098 302372 407108
rect 302204 406918 302260 406928
rect 298956 381938 299012 381948
rect 300636 404038 300692 404048
rect 300636 382004 300692 403982
rect 300636 381938 300692 381948
rect 302204 382004 302260 406862
rect 302316 382116 302372 407042
rect 303996 405658 304052 405668
rect 302316 382050 302372 382060
rect 303884 400798 303940 400808
rect 303884 382116 303940 400742
rect 303884 382050 303940 382060
rect 302204 381938 302260 381948
rect 303996 382004 304052 405602
rect 303996 381938 304052 381948
rect 295596 381602 295652 381612
rect 305676 381668 305732 407582
rect 305676 381602 305732 381612
rect 312618 400350 313238 409194
rect 312618 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 313238 400350
rect 312618 400226 313238 400294
rect 312618 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 313238 400226
rect 312618 400102 313238 400170
rect 312618 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 313238 400102
rect 312618 399978 313238 400046
rect 312618 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 313238 399978
rect 312618 382350 313238 399922
rect 316338 406350 316958 409194
rect 316338 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 316958 406350
rect 316338 406226 316958 406294
rect 316338 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 316958 406226
rect 316338 406102 316958 406170
rect 316338 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 316958 406102
rect 316338 405978 316958 406046
rect 316338 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 316958 405978
rect 312618 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 313238 382350
rect 312618 382226 313238 382294
rect 312618 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 313238 382226
rect 312618 382102 313238 382170
rect 312618 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 313238 382102
rect 312618 381978 313238 382046
rect 312618 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 313238 381978
rect 313404 395578 313460 395588
rect 313404 382004 313460 395522
rect 313404 381938 313460 381948
rect 316338 388350 316958 405922
rect 316338 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 316958 388350
rect 316338 388226 316958 388294
rect 328524 407652 328580 407662
rect 316338 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 316958 388226
rect 316338 388102 316958 388170
rect 316338 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 316958 388102
rect 316338 387978 316958 388046
rect 316338 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 316958 387978
rect 293916 381378 293972 381388
rect 312618 379126 313238 381922
rect 316338 379126 316958 387922
rect 317436 388276 317492 388286
rect 317436 387298 317492 388220
rect 317436 387232 317492 387242
rect 327404 385252 327460 385262
rect 215180 378952 215236 378962
rect 213836 378772 213892 378782
rect 230528 370350 230848 370384
rect 230528 370294 230598 370350
rect 230654 370294 230722 370350
rect 230778 370294 230848 370350
rect 230528 370226 230848 370294
rect 230528 370170 230598 370226
rect 230654 370170 230722 370226
rect 230778 370170 230848 370226
rect 230528 370102 230848 370170
rect 230528 370046 230598 370102
rect 230654 370046 230722 370102
rect 230778 370046 230848 370102
rect 230528 369978 230848 370046
rect 230528 369922 230598 369978
rect 230654 369922 230722 369978
rect 230778 369922 230848 369978
rect 230528 369888 230848 369922
rect 261248 370350 261568 370384
rect 261248 370294 261318 370350
rect 261374 370294 261442 370350
rect 261498 370294 261568 370350
rect 261248 370226 261568 370294
rect 261248 370170 261318 370226
rect 261374 370170 261442 370226
rect 261498 370170 261568 370226
rect 261248 370102 261568 370170
rect 261248 370046 261318 370102
rect 261374 370046 261442 370102
rect 261498 370046 261568 370102
rect 261248 369978 261568 370046
rect 261248 369922 261318 369978
rect 261374 369922 261442 369978
rect 261498 369922 261568 369978
rect 261248 369888 261568 369922
rect 291968 370350 292288 370384
rect 291968 370294 292038 370350
rect 292094 370294 292162 370350
rect 292218 370294 292288 370350
rect 291968 370226 292288 370294
rect 291968 370170 292038 370226
rect 292094 370170 292162 370226
rect 292218 370170 292288 370226
rect 291968 370102 292288 370170
rect 291968 370046 292038 370102
rect 292094 370046 292162 370102
rect 292218 370046 292288 370102
rect 291968 369978 292288 370046
rect 291968 369922 292038 369978
rect 292094 369922 292162 369978
rect 292218 369922 292288 369978
rect 291968 369888 292288 369922
rect 322688 370350 323008 370384
rect 322688 370294 322758 370350
rect 322814 370294 322882 370350
rect 322938 370294 323008 370350
rect 322688 370226 323008 370294
rect 322688 370170 322758 370226
rect 322814 370170 322882 370226
rect 322938 370170 323008 370226
rect 322688 370102 323008 370170
rect 322688 370046 322758 370102
rect 322814 370046 322882 370102
rect 322938 370046 323008 370102
rect 322688 369978 323008 370046
rect 322688 369922 322758 369978
rect 322814 369922 322882 369978
rect 322938 369922 323008 369978
rect 322688 369888 323008 369922
rect 215168 364350 215488 364384
rect 215168 364294 215238 364350
rect 215294 364294 215362 364350
rect 215418 364294 215488 364350
rect 215168 364226 215488 364294
rect 215168 364170 215238 364226
rect 215294 364170 215362 364226
rect 215418 364170 215488 364226
rect 215168 364102 215488 364170
rect 215168 364046 215238 364102
rect 215294 364046 215362 364102
rect 215418 364046 215488 364102
rect 215168 363978 215488 364046
rect 215168 363922 215238 363978
rect 215294 363922 215362 363978
rect 215418 363922 215488 363978
rect 215168 363888 215488 363922
rect 245888 364350 246208 364384
rect 245888 364294 245958 364350
rect 246014 364294 246082 364350
rect 246138 364294 246208 364350
rect 245888 364226 246208 364294
rect 245888 364170 245958 364226
rect 246014 364170 246082 364226
rect 246138 364170 246208 364226
rect 245888 364102 246208 364170
rect 245888 364046 245958 364102
rect 246014 364046 246082 364102
rect 246138 364046 246208 364102
rect 245888 363978 246208 364046
rect 245888 363922 245958 363978
rect 246014 363922 246082 363978
rect 246138 363922 246208 363978
rect 245888 363888 246208 363922
rect 276608 364350 276928 364384
rect 276608 364294 276678 364350
rect 276734 364294 276802 364350
rect 276858 364294 276928 364350
rect 276608 364226 276928 364294
rect 276608 364170 276678 364226
rect 276734 364170 276802 364226
rect 276858 364170 276928 364226
rect 276608 364102 276928 364170
rect 276608 364046 276678 364102
rect 276734 364046 276802 364102
rect 276858 364046 276928 364102
rect 276608 363978 276928 364046
rect 276608 363922 276678 363978
rect 276734 363922 276802 363978
rect 276858 363922 276928 363978
rect 276608 363888 276928 363922
rect 307328 364350 307648 364384
rect 307328 364294 307398 364350
rect 307454 364294 307522 364350
rect 307578 364294 307648 364350
rect 307328 364226 307648 364294
rect 307328 364170 307398 364226
rect 307454 364170 307522 364226
rect 307578 364170 307648 364226
rect 307328 364102 307648 364170
rect 307328 364046 307398 364102
rect 307454 364046 307522 364102
rect 307578 364046 307648 364102
rect 307328 363978 307648 364046
rect 307328 363922 307398 363978
rect 307454 363922 307522 363978
rect 307578 363922 307648 363978
rect 307328 363888 307648 363922
rect 327404 360838 327460 385196
rect 327404 360772 327460 360782
rect 328412 379738 328468 379748
rect 230528 352350 230848 352384
rect 230528 352294 230598 352350
rect 230654 352294 230722 352350
rect 230778 352294 230848 352350
rect 230528 352226 230848 352294
rect 230528 352170 230598 352226
rect 230654 352170 230722 352226
rect 230778 352170 230848 352226
rect 230528 352102 230848 352170
rect 230528 352046 230598 352102
rect 230654 352046 230722 352102
rect 230778 352046 230848 352102
rect 230528 351978 230848 352046
rect 230528 351922 230598 351978
rect 230654 351922 230722 351978
rect 230778 351922 230848 351978
rect 230528 351888 230848 351922
rect 261248 352350 261568 352384
rect 261248 352294 261318 352350
rect 261374 352294 261442 352350
rect 261498 352294 261568 352350
rect 261248 352226 261568 352294
rect 261248 352170 261318 352226
rect 261374 352170 261442 352226
rect 261498 352170 261568 352226
rect 261248 352102 261568 352170
rect 261248 352046 261318 352102
rect 261374 352046 261442 352102
rect 261498 352046 261568 352102
rect 261248 351978 261568 352046
rect 261248 351922 261318 351978
rect 261374 351922 261442 351978
rect 261498 351922 261568 351978
rect 261248 351888 261568 351922
rect 291968 352350 292288 352384
rect 291968 352294 292038 352350
rect 292094 352294 292162 352350
rect 292218 352294 292288 352350
rect 291968 352226 292288 352294
rect 291968 352170 292038 352226
rect 292094 352170 292162 352226
rect 292218 352170 292288 352226
rect 291968 352102 292288 352170
rect 291968 352046 292038 352102
rect 292094 352046 292162 352102
rect 292218 352046 292288 352102
rect 291968 351978 292288 352046
rect 291968 351922 292038 351978
rect 292094 351922 292162 351978
rect 292218 351922 292288 351978
rect 291968 351888 292288 351922
rect 322688 352350 323008 352384
rect 322688 352294 322758 352350
rect 322814 352294 322882 352350
rect 322938 352294 323008 352350
rect 322688 352226 323008 352294
rect 322688 352170 322758 352226
rect 322814 352170 322882 352226
rect 322938 352170 323008 352226
rect 322688 352102 323008 352170
rect 322688 352046 322758 352102
rect 322814 352046 322882 352102
rect 322938 352046 323008 352102
rect 322688 351978 323008 352046
rect 322688 351922 322758 351978
rect 322814 351922 322882 351978
rect 322938 351922 323008 351978
rect 322688 351888 323008 351922
rect 215168 346350 215488 346384
rect 215168 346294 215238 346350
rect 215294 346294 215362 346350
rect 215418 346294 215488 346350
rect 215168 346226 215488 346294
rect 215168 346170 215238 346226
rect 215294 346170 215362 346226
rect 215418 346170 215488 346226
rect 215168 346102 215488 346170
rect 215168 346046 215238 346102
rect 215294 346046 215362 346102
rect 215418 346046 215488 346102
rect 215168 345978 215488 346046
rect 215168 345922 215238 345978
rect 215294 345922 215362 345978
rect 215418 345922 215488 345978
rect 215168 345888 215488 345922
rect 245888 346350 246208 346384
rect 245888 346294 245958 346350
rect 246014 346294 246082 346350
rect 246138 346294 246208 346350
rect 245888 346226 246208 346294
rect 245888 346170 245958 346226
rect 246014 346170 246082 346226
rect 246138 346170 246208 346226
rect 245888 346102 246208 346170
rect 245888 346046 245958 346102
rect 246014 346046 246082 346102
rect 246138 346046 246208 346102
rect 245888 345978 246208 346046
rect 245888 345922 245958 345978
rect 246014 345922 246082 345978
rect 246138 345922 246208 345978
rect 245888 345888 246208 345922
rect 276608 346350 276928 346384
rect 276608 346294 276678 346350
rect 276734 346294 276802 346350
rect 276858 346294 276928 346350
rect 276608 346226 276928 346294
rect 276608 346170 276678 346226
rect 276734 346170 276802 346226
rect 276858 346170 276928 346226
rect 276608 346102 276928 346170
rect 276608 346046 276678 346102
rect 276734 346046 276802 346102
rect 276858 346046 276928 346102
rect 276608 345978 276928 346046
rect 276608 345922 276678 345978
rect 276734 345922 276802 345978
rect 276858 345922 276928 345978
rect 276608 345888 276928 345922
rect 307328 346350 307648 346384
rect 307328 346294 307398 346350
rect 307454 346294 307522 346350
rect 307578 346294 307648 346350
rect 307328 346226 307648 346294
rect 307328 346170 307398 346226
rect 307454 346170 307522 346226
rect 307578 346170 307648 346226
rect 307328 346102 307648 346170
rect 307328 346046 307398 346102
rect 307454 346046 307522 346102
rect 307578 346046 307648 346102
rect 307328 345978 307648 346046
rect 307328 345922 307398 345978
rect 307454 345922 307522 345978
rect 307578 345922 307648 345978
rect 307328 345888 307648 345922
rect 230528 334350 230848 334384
rect 230528 334294 230598 334350
rect 230654 334294 230722 334350
rect 230778 334294 230848 334350
rect 230528 334226 230848 334294
rect 230528 334170 230598 334226
rect 230654 334170 230722 334226
rect 230778 334170 230848 334226
rect 230528 334102 230848 334170
rect 230528 334046 230598 334102
rect 230654 334046 230722 334102
rect 230778 334046 230848 334102
rect 230528 333978 230848 334046
rect 230528 333922 230598 333978
rect 230654 333922 230722 333978
rect 230778 333922 230848 333978
rect 230528 333888 230848 333922
rect 261248 334350 261568 334384
rect 261248 334294 261318 334350
rect 261374 334294 261442 334350
rect 261498 334294 261568 334350
rect 261248 334226 261568 334294
rect 261248 334170 261318 334226
rect 261374 334170 261442 334226
rect 261498 334170 261568 334226
rect 261248 334102 261568 334170
rect 261248 334046 261318 334102
rect 261374 334046 261442 334102
rect 261498 334046 261568 334102
rect 261248 333978 261568 334046
rect 261248 333922 261318 333978
rect 261374 333922 261442 333978
rect 261498 333922 261568 333978
rect 261248 333888 261568 333922
rect 291968 334350 292288 334384
rect 291968 334294 292038 334350
rect 292094 334294 292162 334350
rect 292218 334294 292288 334350
rect 291968 334226 292288 334294
rect 291968 334170 292038 334226
rect 292094 334170 292162 334226
rect 292218 334170 292288 334226
rect 291968 334102 292288 334170
rect 291968 334046 292038 334102
rect 292094 334046 292162 334102
rect 292218 334046 292288 334102
rect 291968 333978 292288 334046
rect 291968 333922 292038 333978
rect 292094 333922 292162 333978
rect 292218 333922 292288 333978
rect 291968 333888 292288 333922
rect 322688 334350 323008 334384
rect 322688 334294 322758 334350
rect 322814 334294 322882 334350
rect 322938 334294 323008 334350
rect 322688 334226 323008 334294
rect 322688 334170 322758 334226
rect 322814 334170 322882 334226
rect 322938 334170 323008 334226
rect 322688 334102 323008 334170
rect 322688 334046 322758 334102
rect 322814 334046 322882 334102
rect 322938 334046 323008 334102
rect 322688 333978 323008 334046
rect 322688 333922 322758 333978
rect 322814 333922 322882 333978
rect 322938 333922 323008 333978
rect 322688 333888 323008 333922
rect 215168 328350 215488 328384
rect 215168 328294 215238 328350
rect 215294 328294 215362 328350
rect 215418 328294 215488 328350
rect 215168 328226 215488 328294
rect 215168 328170 215238 328226
rect 215294 328170 215362 328226
rect 215418 328170 215488 328226
rect 215168 328102 215488 328170
rect 215168 328046 215238 328102
rect 215294 328046 215362 328102
rect 215418 328046 215488 328102
rect 215168 327978 215488 328046
rect 215168 327922 215238 327978
rect 215294 327922 215362 327978
rect 215418 327922 215488 327978
rect 215168 327888 215488 327922
rect 245888 328350 246208 328384
rect 245888 328294 245958 328350
rect 246014 328294 246082 328350
rect 246138 328294 246208 328350
rect 245888 328226 246208 328294
rect 245888 328170 245958 328226
rect 246014 328170 246082 328226
rect 246138 328170 246208 328226
rect 245888 328102 246208 328170
rect 245888 328046 245958 328102
rect 246014 328046 246082 328102
rect 246138 328046 246208 328102
rect 245888 327978 246208 328046
rect 245888 327922 245958 327978
rect 246014 327922 246082 327978
rect 246138 327922 246208 327978
rect 245888 327888 246208 327922
rect 276608 328350 276928 328384
rect 276608 328294 276678 328350
rect 276734 328294 276802 328350
rect 276858 328294 276928 328350
rect 276608 328226 276928 328294
rect 276608 328170 276678 328226
rect 276734 328170 276802 328226
rect 276858 328170 276928 328226
rect 276608 328102 276928 328170
rect 276608 328046 276678 328102
rect 276734 328046 276802 328102
rect 276858 328046 276928 328102
rect 276608 327978 276928 328046
rect 276608 327922 276678 327978
rect 276734 327922 276802 327978
rect 276858 327922 276928 327978
rect 276608 327888 276928 327922
rect 307328 328350 307648 328384
rect 307328 328294 307398 328350
rect 307454 328294 307522 328350
rect 307578 328294 307648 328350
rect 307328 328226 307648 328294
rect 307328 328170 307398 328226
rect 307454 328170 307522 328226
rect 307578 328170 307648 328226
rect 307328 328102 307648 328170
rect 307328 328046 307398 328102
rect 307454 328046 307522 328102
rect 307578 328046 307648 328102
rect 307328 327978 307648 328046
rect 307328 327922 307398 327978
rect 307454 327922 307522 327978
rect 307578 327922 307648 327978
rect 307328 327888 307648 327922
rect 230528 316350 230848 316384
rect 230528 316294 230598 316350
rect 230654 316294 230722 316350
rect 230778 316294 230848 316350
rect 230528 316226 230848 316294
rect 230528 316170 230598 316226
rect 230654 316170 230722 316226
rect 230778 316170 230848 316226
rect 230528 316102 230848 316170
rect 230528 316046 230598 316102
rect 230654 316046 230722 316102
rect 230778 316046 230848 316102
rect 230528 315978 230848 316046
rect 230528 315922 230598 315978
rect 230654 315922 230722 315978
rect 230778 315922 230848 315978
rect 230528 315888 230848 315922
rect 261248 316350 261568 316384
rect 261248 316294 261318 316350
rect 261374 316294 261442 316350
rect 261498 316294 261568 316350
rect 261248 316226 261568 316294
rect 261248 316170 261318 316226
rect 261374 316170 261442 316226
rect 261498 316170 261568 316226
rect 261248 316102 261568 316170
rect 261248 316046 261318 316102
rect 261374 316046 261442 316102
rect 261498 316046 261568 316102
rect 261248 315978 261568 316046
rect 261248 315922 261318 315978
rect 261374 315922 261442 315978
rect 261498 315922 261568 315978
rect 261248 315888 261568 315922
rect 291968 316350 292288 316384
rect 291968 316294 292038 316350
rect 292094 316294 292162 316350
rect 292218 316294 292288 316350
rect 291968 316226 292288 316294
rect 291968 316170 292038 316226
rect 292094 316170 292162 316226
rect 292218 316170 292288 316226
rect 291968 316102 292288 316170
rect 291968 316046 292038 316102
rect 292094 316046 292162 316102
rect 292218 316046 292288 316102
rect 291968 315978 292288 316046
rect 291968 315922 292038 315978
rect 292094 315922 292162 315978
rect 292218 315922 292288 315978
rect 291968 315888 292288 315922
rect 322688 316350 323008 316384
rect 322688 316294 322758 316350
rect 322814 316294 322882 316350
rect 322938 316294 323008 316350
rect 322688 316226 323008 316294
rect 322688 316170 322758 316226
rect 322814 316170 322882 316226
rect 322938 316170 323008 316226
rect 322688 316102 323008 316170
rect 322688 316046 322758 316102
rect 322814 316046 322882 316102
rect 322938 316046 323008 316102
rect 322688 315978 323008 316046
rect 322688 315922 322758 315978
rect 322814 315922 322882 315978
rect 322938 315922 323008 315978
rect 322688 315888 323008 315922
rect 328076 311698 328132 311708
rect 215168 310350 215488 310384
rect 215168 310294 215238 310350
rect 215294 310294 215362 310350
rect 215418 310294 215488 310350
rect 215168 310226 215488 310294
rect 215168 310170 215238 310226
rect 215294 310170 215362 310226
rect 215418 310170 215488 310226
rect 215168 310102 215488 310170
rect 215168 310046 215238 310102
rect 215294 310046 215362 310102
rect 215418 310046 215488 310102
rect 215168 309978 215488 310046
rect 215168 309922 215238 309978
rect 215294 309922 215362 309978
rect 215418 309922 215488 309978
rect 215168 309888 215488 309922
rect 245888 310350 246208 310384
rect 245888 310294 245958 310350
rect 246014 310294 246082 310350
rect 246138 310294 246208 310350
rect 245888 310226 246208 310294
rect 245888 310170 245958 310226
rect 246014 310170 246082 310226
rect 246138 310170 246208 310226
rect 245888 310102 246208 310170
rect 245888 310046 245958 310102
rect 246014 310046 246082 310102
rect 246138 310046 246208 310102
rect 245888 309978 246208 310046
rect 245888 309922 245958 309978
rect 246014 309922 246082 309978
rect 246138 309922 246208 309978
rect 245888 309888 246208 309922
rect 276608 310350 276928 310384
rect 276608 310294 276678 310350
rect 276734 310294 276802 310350
rect 276858 310294 276928 310350
rect 276608 310226 276928 310294
rect 276608 310170 276678 310226
rect 276734 310170 276802 310226
rect 276858 310170 276928 310226
rect 276608 310102 276928 310170
rect 276608 310046 276678 310102
rect 276734 310046 276802 310102
rect 276858 310046 276928 310102
rect 276608 309978 276928 310046
rect 276608 309922 276678 309978
rect 276734 309922 276802 309978
rect 276858 309922 276928 309978
rect 276608 309888 276928 309922
rect 307328 310350 307648 310384
rect 307328 310294 307398 310350
rect 307454 310294 307522 310350
rect 307578 310294 307648 310350
rect 307328 310226 307648 310294
rect 307328 310170 307398 310226
rect 307454 310170 307522 310226
rect 307578 310170 307648 310226
rect 307328 310102 307648 310170
rect 307328 310046 307398 310102
rect 307454 310046 307522 310102
rect 307578 310046 307648 310102
rect 307328 309978 307648 310046
rect 307328 309922 307398 309978
rect 307454 309922 307522 309978
rect 307578 309922 307648 309978
rect 307328 309888 307648 309922
rect 230528 298350 230848 298384
rect 230528 298294 230598 298350
rect 230654 298294 230722 298350
rect 230778 298294 230848 298350
rect 230528 298226 230848 298294
rect 230528 298170 230598 298226
rect 230654 298170 230722 298226
rect 230778 298170 230848 298226
rect 230528 298102 230848 298170
rect 230528 298046 230598 298102
rect 230654 298046 230722 298102
rect 230778 298046 230848 298102
rect 230528 297978 230848 298046
rect 230528 297922 230598 297978
rect 230654 297922 230722 297978
rect 230778 297922 230848 297978
rect 230528 297888 230848 297922
rect 261248 298350 261568 298384
rect 261248 298294 261318 298350
rect 261374 298294 261442 298350
rect 261498 298294 261568 298350
rect 261248 298226 261568 298294
rect 261248 298170 261318 298226
rect 261374 298170 261442 298226
rect 261498 298170 261568 298226
rect 261248 298102 261568 298170
rect 261248 298046 261318 298102
rect 261374 298046 261442 298102
rect 261498 298046 261568 298102
rect 261248 297978 261568 298046
rect 261248 297922 261318 297978
rect 261374 297922 261442 297978
rect 261498 297922 261568 297978
rect 261248 297888 261568 297922
rect 291968 298350 292288 298384
rect 291968 298294 292038 298350
rect 292094 298294 292162 298350
rect 292218 298294 292288 298350
rect 291968 298226 292288 298294
rect 291968 298170 292038 298226
rect 292094 298170 292162 298226
rect 292218 298170 292288 298226
rect 291968 298102 292288 298170
rect 291968 298046 292038 298102
rect 292094 298046 292162 298102
rect 292218 298046 292288 298102
rect 291968 297978 292288 298046
rect 291968 297922 292038 297978
rect 292094 297922 292162 297978
rect 292218 297922 292288 297978
rect 291968 297888 292288 297922
rect 322688 298350 323008 298384
rect 322688 298294 322758 298350
rect 322814 298294 322882 298350
rect 322938 298294 323008 298350
rect 322688 298226 323008 298294
rect 322688 298170 322758 298226
rect 322814 298170 322882 298226
rect 322938 298170 323008 298226
rect 322688 298102 323008 298170
rect 322688 298046 322758 298102
rect 322814 298046 322882 298102
rect 322938 298046 323008 298102
rect 322688 297978 323008 298046
rect 322688 297922 322758 297978
rect 322814 297922 322882 297978
rect 322938 297922 323008 297978
rect 322688 297888 323008 297922
rect 215168 292350 215488 292384
rect 215168 292294 215238 292350
rect 215294 292294 215362 292350
rect 215418 292294 215488 292350
rect 215168 292226 215488 292294
rect 215168 292170 215238 292226
rect 215294 292170 215362 292226
rect 215418 292170 215488 292226
rect 215168 292102 215488 292170
rect 215168 292046 215238 292102
rect 215294 292046 215362 292102
rect 215418 292046 215488 292102
rect 215168 291978 215488 292046
rect 215168 291922 215238 291978
rect 215294 291922 215362 291978
rect 215418 291922 215488 291978
rect 215168 291888 215488 291922
rect 245888 292350 246208 292384
rect 245888 292294 245958 292350
rect 246014 292294 246082 292350
rect 246138 292294 246208 292350
rect 245888 292226 246208 292294
rect 245888 292170 245958 292226
rect 246014 292170 246082 292226
rect 246138 292170 246208 292226
rect 245888 292102 246208 292170
rect 245888 292046 245958 292102
rect 246014 292046 246082 292102
rect 246138 292046 246208 292102
rect 245888 291978 246208 292046
rect 245888 291922 245958 291978
rect 246014 291922 246082 291978
rect 246138 291922 246208 291978
rect 245888 291888 246208 291922
rect 276608 292350 276928 292384
rect 276608 292294 276678 292350
rect 276734 292294 276802 292350
rect 276858 292294 276928 292350
rect 276608 292226 276928 292294
rect 276608 292170 276678 292226
rect 276734 292170 276802 292226
rect 276858 292170 276928 292226
rect 276608 292102 276928 292170
rect 276608 292046 276678 292102
rect 276734 292046 276802 292102
rect 276858 292046 276928 292102
rect 276608 291978 276928 292046
rect 276608 291922 276678 291978
rect 276734 291922 276802 291978
rect 276858 291922 276928 291978
rect 276608 291888 276928 291922
rect 307328 292350 307648 292384
rect 307328 292294 307398 292350
rect 307454 292294 307522 292350
rect 307578 292294 307648 292350
rect 307328 292226 307648 292294
rect 307328 292170 307398 292226
rect 307454 292170 307522 292226
rect 307578 292170 307648 292226
rect 307328 292102 307648 292170
rect 307328 292046 307398 292102
rect 307454 292046 307522 292102
rect 307578 292046 307648 292102
rect 307328 291978 307648 292046
rect 307328 291922 307398 291978
rect 307454 291922 307522 291978
rect 307578 291922 307648 291978
rect 307328 291888 307648 291922
rect 230528 280350 230848 280384
rect 230528 280294 230598 280350
rect 230654 280294 230722 280350
rect 230778 280294 230848 280350
rect 230528 280226 230848 280294
rect 230528 280170 230598 280226
rect 230654 280170 230722 280226
rect 230778 280170 230848 280226
rect 230528 280102 230848 280170
rect 230528 280046 230598 280102
rect 230654 280046 230722 280102
rect 230778 280046 230848 280102
rect 230528 279978 230848 280046
rect 230528 279922 230598 279978
rect 230654 279922 230722 279978
rect 230778 279922 230848 279978
rect 230528 279888 230848 279922
rect 261248 280350 261568 280384
rect 261248 280294 261318 280350
rect 261374 280294 261442 280350
rect 261498 280294 261568 280350
rect 261248 280226 261568 280294
rect 261248 280170 261318 280226
rect 261374 280170 261442 280226
rect 261498 280170 261568 280226
rect 261248 280102 261568 280170
rect 261248 280046 261318 280102
rect 261374 280046 261442 280102
rect 261498 280046 261568 280102
rect 261248 279978 261568 280046
rect 261248 279922 261318 279978
rect 261374 279922 261442 279978
rect 261498 279922 261568 279978
rect 261248 279888 261568 279922
rect 291968 280350 292288 280384
rect 291968 280294 292038 280350
rect 292094 280294 292162 280350
rect 292218 280294 292288 280350
rect 291968 280226 292288 280294
rect 291968 280170 292038 280226
rect 292094 280170 292162 280226
rect 292218 280170 292288 280226
rect 291968 280102 292288 280170
rect 291968 280046 292038 280102
rect 292094 280046 292162 280102
rect 292218 280046 292288 280102
rect 291968 279978 292288 280046
rect 291968 279922 292038 279978
rect 292094 279922 292162 279978
rect 292218 279922 292288 279978
rect 291968 279888 292288 279922
rect 322688 280350 323008 280384
rect 322688 280294 322758 280350
rect 322814 280294 322882 280350
rect 322938 280294 323008 280350
rect 322688 280226 323008 280294
rect 322688 280170 322758 280226
rect 322814 280170 322882 280226
rect 322938 280170 323008 280226
rect 322688 280102 323008 280170
rect 322688 280046 322758 280102
rect 322814 280046 322882 280102
rect 322938 280046 323008 280102
rect 322688 279978 323008 280046
rect 322688 279922 322758 279978
rect 322814 279922 322882 279978
rect 322938 279922 323008 279978
rect 322688 279888 323008 279922
rect 215168 274350 215488 274384
rect 215168 274294 215238 274350
rect 215294 274294 215362 274350
rect 215418 274294 215488 274350
rect 215168 274226 215488 274294
rect 215168 274170 215238 274226
rect 215294 274170 215362 274226
rect 215418 274170 215488 274226
rect 215168 274102 215488 274170
rect 215168 274046 215238 274102
rect 215294 274046 215362 274102
rect 215418 274046 215488 274102
rect 215168 273978 215488 274046
rect 215168 273922 215238 273978
rect 215294 273922 215362 273978
rect 215418 273922 215488 273978
rect 215168 273888 215488 273922
rect 245888 274350 246208 274384
rect 245888 274294 245958 274350
rect 246014 274294 246082 274350
rect 246138 274294 246208 274350
rect 245888 274226 246208 274294
rect 245888 274170 245958 274226
rect 246014 274170 246082 274226
rect 246138 274170 246208 274226
rect 245888 274102 246208 274170
rect 245888 274046 245958 274102
rect 246014 274046 246082 274102
rect 246138 274046 246208 274102
rect 245888 273978 246208 274046
rect 245888 273922 245958 273978
rect 246014 273922 246082 273978
rect 246138 273922 246208 273978
rect 245888 273888 246208 273922
rect 276608 274350 276928 274384
rect 276608 274294 276678 274350
rect 276734 274294 276802 274350
rect 276858 274294 276928 274350
rect 276608 274226 276928 274294
rect 276608 274170 276678 274226
rect 276734 274170 276802 274226
rect 276858 274170 276928 274226
rect 276608 274102 276928 274170
rect 276608 274046 276678 274102
rect 276734 274046 276802 274102
rect 276858 274046 276928 274102
rect 276608 273978 276928 274046
rect 276608 273922 276678 273978
rect 276734 273922 276802 273978
rect 276858 273922 276928 273978
rect 276608 273888 276928 273922
rect 307328 274350 307648 274384
rect 307328 274294 307398 274350
rect 307454 274294 307522 274350
rect 307578 274294 307648 274350
rect 307328 274226 307648 274294
rect 307328 274170 307398 274226
rect 307454 274170 307522 274226
rect 307578 274170 307648 274226
rect 307328 274102 307648 274170
rect 307328 274046 307398 274102
rect 307454 274046 307522 274102
rect 307578 274046 307648 274102
rect 307328 273978 307648 274046
rect 307328 273922 307398 273978
rect 307454 273922 307522 273978
rect 307578 273922 307648 273978
rect 307328 273888 307648 273922
rect 230528 262350 230848 262384
rect 230528 262294 230598 262350
rect 230654 262294 230722 262350
rect 230778 262294 230848 262350
rect 230528 262226 230848 262294
rect 230528 262170 230598 262226
rect 230654 262170 230722 262226
rect 230778 262170 230848 262226
rect 230528 262102 230848 262170
rect 230528 262046 230598 262102
rect 230654 262046 230722 262102
rect 230778 262046 230848 262102
rect 230528 261978 230848 262046
rect 230528 261922 230598 261978
rect 230654 261922 230722 261978
rect 230778 261922 230848 261978
rect 230528 261888 230848 261922
rect 261248 262350 261568 262384
rect 261248 262294 261318 262350
rect 261374 262294 261442 262350
rect 261498 262294 261568 262350
rect 261248 262226 261568 262294
rect 261248 262170 261318 262226
rect 261374 262170 261442 262226
rect 261498 262170 261568 262226
rect 261248 262102 261568 262170
rect 261248 262046 261318 262102
rect 261374 262046 261442 262102
rect 261498 262046 261568 262102
rect 261248 261978 261568 262046
rect 261248 261922 261318 261978
rect 261374 261922 261442 261978
rect 261498 261922 261568 261978
rect 261248 261888 261568 261922
rect 291968 262350 292288 262384
rect 291968 262294 292038 262350
rect 292094 262294 292162 262350
rect 292218 262294 292288 262350
rect 291968 262226 292288 262294
rect 291968 262170 292038 262226
rect 292094 262170 292162 262226
rect 292218 262170 292288 262226
rect 291968 262102 292288 262170
rect 291968 262046 292038 262102
rect 292094 262046 292162 262102
rect 292218 262046 292288 262102
rect 291968 261978 292288 262046
rect 291968 261922 292038 261978
rect 292094 261922 292162 261978
rect 292218 261922 292288 261978
rect 291968 261888 292288 261922
rect 322688 262350 323008 262384
rect 322688 262294 322758 262350
rect 322814 262294 322882 262350
rect 322938 262294 323008 262350
rect 322688 262226 323008 262294
rect 322688 262170 322758 262226
rect 322814 262170 322882 262226
rect 322938 262170 323008 262226
rect 322688 262102 323008 262170
rect 322688 262046 322758 262102
rect 322814 262046 322882 262102
rect 322938 262046 323008 262102
rect 322688 261978 323008 262046
rect 322688 261922 322758 261978
rect 322814 261922 322882 261978
rect 322938 261922 323008 261978
rect 322688 261888 323008 261922
rect 327964 260398 328020 260408
rect 215168 256350 215488 256384
rect 215168 256294 215238 256350
rect 215294 256294 215362 256350
rect 215418 256294 215488 256350
rect 215168 256226 215488 256294
rect 215168 256170 215238 256226
rect 215294 256170 215362 256226
rect 215418 256170 215488 256226
rect 215168 256102 215488 256170
rect 215168 256046 215238 256102
rect 215294 256046 215362 256102
rect 215418 256046 215488 256102
rect 215168 255978 215488 256046
rect 215168 255922 215238 255978
rect 215294 255922 215362 255978
rect 215418 255922 215488 255978
rect 215168 255888 215488 255922
rect 245888 256350 246208 256384
rect 245888 256294 245958 256350
rect 246014 256294 246082 256350
rect 246138 256294 246208 256350
rect 245888 256226 246208 256294
rect 245888 256170 245958 256226
rect 246014 256170 246082 256226
rect 246138 256170 246208 256226
rect 245888 256102 246208 256170
rect 245888 256046 245958 256102
rect 246014 256046 246082 256102
rect 246138 256046 246208 256102
rect 245888 255978 246208 256046
rect 245888 255922 245958 255978
rect 246014 255922 246082 255978
rect 246138 255922 246208 255978
rect 245888 255888 246208 255922
rect 276608 256350 276928 256384
rect 276608 256294 276678 256350
rect 276734 256294 276802 256350
rect 276858 256294 276928 256350
rect 276608 256226 276928 256294
rect 276608 256170 276678 256226
rect 276734 256170 276802 256226
rect 276858 256170 276928 256226
rect 276608 256102 276928 256170
rect 276608 256046 276678 256102
rect 276734 256046 276802 256102
rect 276858 256046 276928 256102
rect 276608 255978 276928 256046
rect 276608 255922 276678 255978
rect 276734 255922 276802 255978
rect 276858 255922 276928 255978
rect 276608 255888 276928 255922
rect 307328 256350 307648 256384
rect 307328 256294 307398 256350
rect 307454 256294 307522 256350
rect 307578 256294 307648 256350
rect 307328 256226 307648 256294
rect 307328 256170 307398 256226
rect 307454 256170 307522 256226
rect 307578 256170 307648 256226
rect 307328 256102 307648 256170
rect 307328 256046 307398 256102
rect 307454 256046 307522 256102
rect 307578 256046 307648 256102
rect 307328 255978 307648 256046
rect 307328 255922 307398 255978
rect 307454 255922 307522 255978
rect 307578 255922 307648 255978
rect 307328 255888 307648 255922
rect 327404 248158 327460 248168
rect 230528 244350 230848 244384
rect 230528 244294 230598 244350
rect 230654 244294 230722 244350
rect 230778 244294 230848 244350
rect 230528 244226 230848 244294
rect 230528 244170 230598 244226
rect 230654 244170 230722 244226
rect 230778 244170 230848 244226
rect 230528 244102 230848 244170
rect 230528 244046 230598 244102
rect 230654 244046 230722 244102
rect 230778 244046 230848 244102
rect 230528 243978 230848 244046
rect 230528 243922 230598 243978
rect 230654 243922 230722 243978
rect 230778 243922 230848 243978
rect 230528 243888 230848 243922
rect 261248 244350 261568 244384
rect 261248 244294 261318 244350
rect 261374 244294 261442 244350
rect 261498 244294 261568 244350
rect 261248 244226 261568 244294
rect 261248 244170 261318 244226
rect 261374 244170 261442 244226
rect 261498 244170 261568 244226
rect 261248 244102 261568 244170
rect 261248 244046 261318 244102
rect 261374 244046 261442 244102
rect 261498 244046 261568 244102
rect 261248 243978 261568 244046
rect 261248 243922 261318 243978
rect 261374 243922 261442 243978
rect 261498 243922 261568 243978
rect 261248 243888 261568 243922
rect 291968 244350 292288 244384
rect 291968 244294 292038 244350
rect 292094 244294 292162 244350
rect 292218 244294 292288 244350
rect 291968 244226 292288 244294
rect 291968 244170 292038 244226
rect 292094 244170 292162 244226
rect 292218 244170 292288 244226
rect 291968 244102 292288 244170
rect 291968 244046 292038 244102
rect 292094 244046 292162 244102
rect 292218 244046 292288 244102
rect 291968 243978 292288 244046
rect 291968 243922 292038 243978
rect 292094 243922 292162 243978
rect 292218 243922 292288 243978
rect 291968 243888 292288 243922
rect 322688 244350 323008 244384
rect 322688 244294 322758 244350
rect 322814 244294 322882 244350
rect 322938 244294 323008 244350
rect 322688 244226 323008 244294
rect 322688 244170 322758 244226
rect 322814 244170 322882 244226
rect 322938 244170 323008 244226
rect 322688 244102 323008 244170
rect 322688 244046 322758 244102
rect 322814 244046 322882 244102
rect 322938 244046 323008 244102
rect 322688 243978 323008 244046
rect 322688 243922 322758 243978
rect 322814 243922 322882 243978
rect 322938 243922 323008 243978
rect 322688 243888 323008 243922
rect 326732 240958 326788 240968
rect 326620 240778 326676 240788
rect 326508 240660 326564 240670
rect 294812 240436 294868 240446
rect 268044 239764 268100 239774
rect 204876 219986 204932 219996
rect 220458 238350 221078 239082
rect 220458 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 221078 238350
rect 220458 238226 221078 238294
rect 220458 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 221078 238226
rect 220458 238102 221078 238170
rect 220458 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 221078 238102
rect 220458 237978 221078 238046
rect 220458 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 221078 237978
rect 220458 220350 221078 237922
rect 220458 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 221078 220350
rect 220458 220226 221078 220294
rect 220458 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 221078 220226
rect 220458 220102 221078 220170
rect 220458 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 221078 220102
rect 203084 205792 203140 205802
rect 220458 219978 221078 220046
rect 220458 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 221078 219978
rect 220458 205590 221078 219922
rect 224178 226350 224798 239082
rect 251178 238350 251798 239082
rect 251178 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 251798 238350
rect 251178 238226 251798 238294
rect 251178 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 251798 238226
rect 251178 238102 251798 238170
rect 251178 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 251798 238102
rect 251178 237978 251798 238046
rect 251178 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 251798 237978
rect 235116 237188 235172 237198
rect 235116 237094 235172 237122
rect 234220 237076 234276 237086
rect 234220 236998 234276 237020
rect 224178 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 224798 226350
rect 224178 226226 224798 226294
rect 224178 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 224798 226226
rect 224178 226102 224798 226170
rect 224178 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 224798 226102
rect 224178 225978 224798 226046
rect 224178 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 224798 225978
rect 224178 208350 224798 225922
rect 224178 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 224798 208350
rect 224178 208226 224798 208294
rect 224178 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 224798 208226
rect 224178 208102 224798 208170
rect 224178 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 224798 208102
rect 224178 207978 224798 208046
rect 224178 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 224798 207978
rect 224178 205590 224798 207922
rect 226716 236964 226772 236974
rect 226716 204058 226772 236908
rect 231756 236964 231812 236974
rect 231756 206578 231812 236908
rect 233436 236964 233492 236974
rect 234220 236932 234276 236942
rect 233436 207478 233492 236908
rect 251178 220350 251798 237922
rect 251178 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 251798 220350
rect 251178 220226 251798 220294
rect 251178 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 251798 220226
rect 251178 220102 251798 220170
rect 251178 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 251798 220102
rect 251178 219978 251798 220046
rect 251178 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 251798 219978
rect 241388 210084 241444 210094
rect 241388 208964 241444 210028
rect 241388 208898 241444 208908
rect 233436 207412 233492 207422
rect 231756 206512 231812 206522
rect 251178 205590 251798 219922
rect 254492 234276 254548 234286
rect 254492 204238 254548 234220
rect 254898 226350 255518 239082
rect 267148 237178 267204 237188
rect 254898 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 255518 226350
rect 254898 226226 255518 226294
rect 254898 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 255518 226226
rect 254898 226102 255518 226170
rect 254898 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 255518 226102
rect 254898 225978 255518 226046
rect 254898 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 255518 225978
rect 254898 208350 255518 225922
rect 254898 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 255518 208350
rect 254898 208226 255518 208294
rect 254898 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 255518 208226
rect 254898 208102 255518 208170
rect 254898 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 255518 208102
rect 254898 207978 255518 208046
rect 254898 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 255518 207978
rect 254898 205590 255518 207922
rect 265244 237076 265300 237086
rect 265244 206578 265300 237020
rect 265244 206512 265300 206522
rect 265356 236964 265412 236974
rect 265356 204418 265412 236908
rect 266812 236964 266868 236974
rect 266812 206218 266868 236908
rect 267036 236964 267092 236974
rect 266812 206152 266868 206162
rect 266924 235060 266980 235070
rect 265356 204352 265412 204362
rect 254492 204172 254548 204182
rect 226716 203992 226772 204002
rect 44448 202350 44768 202384
rect 44448 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 44768 202350
rect 44448 202226 44768 202294
rect 44448 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 44768 202226
rect 44448 202102 44768 202170
rect 44448 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 44768 202102
rect 44448 201978 44768 202046
rect 44448 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 44768 201978
rect 44448 201888 44768 201922
rect 75168 202350 75488 202384
rect 75168 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 75488 202350
rect 75168 202226 75488 202294
rect 75168 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 75488 202226
rect 75168 202102 75488 202170
rect 75168 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 75488 202102
rect 75168 201978 75488 202046
rect 75168 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 75488 201978
rect 75168 201888 75488 201922
rect 105888 202350 106208 202384
rect 105888 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 106208 202350
rect 105888 202226 106208 202294
rect 105888 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 106208 202226
rect 105888 202102 106208 202170
rect 105888 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 106208 202102
rect 105888 201978 106208 202046
rect 105888 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 106208 201978
rect 105888 201888 106208 201922
rect 136608 202350 136928 202384
rect 136608 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 136928 202350
rect 136608 202226 136928 202294
rect 136608 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 136928 202226
rect 136608 202102 136928 202170
rect 136608 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 136928 202102
rect 136608 201978 136928 202046
rect 136608 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 136928 201978
rect 136608 201888 136928 201922
rect 167328 202350 167648 202384
rect 167328 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 167648 202350
rect 167328 202226 167648 202294
rect 167328 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 167648 202226
rect 167328 202102 167648 202170
rect 167328 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 167648 202102
rect 167328 201978 167648 202046
rect 167328 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 167648 201978
rect 167328 201888 167648 201922
rect 198048 202350 198368 202384
rect 198048 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 198368 202350
rect 198048 202226 198368 202294
rect 198048 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 198368 202226
rect 198048 202102 198368 202170
rect 198048 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 198368 202102
rect 198048 201978 198368 202046
rect 198048 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 198368 201978
rect 198048 201888 198368 201922
rect 228768 202350 229088 202384
rect 228768 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 229088 202350
rect 228768 202226 229088 202294
rect 228768 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 229088 202226
rect 228768 202102 229088 202170
rect 228768 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 229088 202102
rect 228768 201978 229088 202046
rect 228768 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 229088 201978
rect 228768 201888 229088 201922
rect 259488 202350 259808 202384
rect 259488 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 259808 202350
rect 259488 202226 259808 202294
rect 259488 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 259808 202226
rect 259488 202102 259808 202170
rect 259488 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 259808 202102
rect 259488 201978 259808 202046
rect 259488 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 259808 201978
rect 259488 201888 259808 201922
rect 59808 190350 60128 190384
rect 59808 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 60128 190350
rect 59808 190226 60128 190294
rect 59808 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 60128 190226
rect 59808 190102 60128 190170
rect 59808 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 60128 190102
rect 59808 189978 60128 190046
rect 59808 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 60128 189978
rect 59808 189888 60128 189922
rect 90528 190350 90848 190384
rect 90528 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 90848 190350
rect 90528 190226 90848 190294
rect 90528 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 90848 190226
rect 90528 190102 90848 190170
rect 90528 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 90848 190102
rect 90528 189978 90848 190046
rect 90528 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 90848 189978
rect 90528 189888 90848 189922
rect 121248 190350 121568 190384
rect 121248 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 121568 190350
rect 121248 190226 121568 190294
rect 121248 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 121568 190226
rect 121248 190102 121568 190170
rect 121248 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 121568 190102
rect 121248 189978 121568 190046
rect 121248 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 121568 189978
rect 121248 189888 121568 189922
rect 151968 190350 152288 190384
rect 151968 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 152288 190350
rect 151968 190226 152288 190294
rect 151968 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 152288 190226
rect 151968 190102 152288 190170
rect 151968 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 152288 190102
rect 151968 189978 152288 190046
rect 151968 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 152288 189978
rect 151968 189888 152288 189922
rect 182688 190350 183008 190384
rect 182688 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 183008 190350
rect 182688 190226 183008 190294
rect 182688 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 183008 190226
rect 182688 190102 183008 190170
rect 182688 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 183008 190102
rect 182688 189978 183008 190046
rect 182688 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 183008 189978
rect 182688 189888 183008 189922
rect 213408 190350 213728 190384
rect 213408 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 213728 190350
rect 213408 190226 213728 190294
rect 213408 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 213728 190226
rect 213408 190102 213728 190170
rect 213408 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 213728 190102
rect 213408 189978 213728 190046
rect 213408 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 213728 189978
rect 213408 189888 213728 189922
rect 244128 190350 244448 190384
rect 244128 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 244448 190350
rect 244128 190226 244448 190294
rect 244128 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 244448 190226
rect 244128 190102 244448 190170
rect 244128 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 244448 190102
rect 244128 189978 244448 190046
rect 244128 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 244448 189978
rect 244128 189888 244448 189922
rect 44448 184350 44768 184384
rect 44448 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 44768 184350
rect 44448 184226 44768 184294
rect 44448 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 44768 184226
rect 44448 184102 44768 184170
rect 44448 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 44768 184102
rect 44448 183978 44768 184046
rect 44448 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 44768 183978
rect 44448 183888 44768 183922
rect 75168 184350 75488 184384
rect 75168 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 75488 184350
rect 75168 184226 75488 184294
rect 75168 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 75488 184226
rect 75168 184102 75488 184170
rect 75168 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 75488 184102
rect 75168 183978 75488 184046
rect 75168 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 75488 183978
rect 75168 183888 75488 183922
rect 105888 184350 106208 184384
rect 105888 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 106208 184350
rect 105888 184226 106208 184294
rect 105888 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 106208 184226
rect 105888 184102 106208 184170
rect 105888 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 106208 184102
rect 105888 183978 106208 184046
rect 105888 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 106208 183978
rect 105888 183888 106208 183922
rect 136608 184350 136928 184384
rect 136608 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 136928 184350
rect 136608 184226 136928 184294
rect 136608 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 136928 184226
rect 136608 184102 136928 184170
rect 136608 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 136928 184102
rect 136608 183978 136928 184046
rect 136608 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 136928 183978
rect 136608 183888 136928 183922
rect 167328 184350 167648 184384
rect 167328 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 167648 184350
rect 167328 184226 167648 184294
rect 167328 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 167648 184226
rect 167328 184102 167648 184170
rect 167328 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 167648 184102
rect 167328 183978 167648 184046
rect 167328 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 167648 183978
rect 167328 183888 167648 183922
rect 198048 184350 198368 184384
rect 198048 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 198368 184350
rect 198048 184226 198368 184294
rect 198048 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 198368 184226
rect 198048 184102 198368 184170
rect 198048 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 198368 184102
rect 198048 183978 198368 184046
rect 198048 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 198368 183978
rect 198048 183888 198368 183922
rect 228768 184350 229088 184384
rect 228768 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 229088 184350
rect 228768 184226 229088 184294
rect 228768 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 229088 184226
rect 228768 184102 229088 184170
rect 228768 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 229088 184102
rect 228768 183978 229088 184046
rect 228768 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 229088 183978
rect 228768 183888 229088 183922
rect 259488 184350 259808 184384
rect 259488 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 259808 184350
rect 259488 184226 259808 184294
rect 259488 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 259808 184226
rect 259488 184102 259808 184170
rect 259488 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 259808 184102
rect 259488 183978 259808 184046
rect 259488 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 259808 183978
rect 259488 183888 259808 183922
rect 59808 172350 60128 172384
rect 59808 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 60128 172350
rect 59808 172226 60128 172294
rect 59808 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 60128 172226
rect 59808 172102 60128 172170
rect 59808 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 60128 172102
rect 59808 171978 60128 172046
rect 59808 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 60128 171978
rect 59808 171888 60128 171922
rect 90528 172350 90848 172384
rect 90528 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 90848 172350
rect 90528 172226 90848 172294
rect 90528 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 90848 172226
rect 90528 172102 90848 172170
rect 90528 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 90848 172102
rect 90528 171978 90848 172046
rect 90528 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 90848 171978
rect 90528 171888 90848 171922
rect 121248 172350 121568 172384
rect 121248 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 121568 172350
rect 121248 172226 121568 172294
rect 121248 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 121568 172226
rect 121248 172102 121568 172170
rect 121248 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 121568 172102
rect 121248 171978 121568 172046
rect 121248 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 121568 171978
rect 121248 171888 121568 171922
rect 151968 172350 152288 172384
rect 151968 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 152288 172350
rect 151968 172226 152288 172294
rect 151968 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 152288 172226
rect 151968 172102 152288 172170
rect 151968 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 152288 172102
rect 151968 171978 152288 172046
rect 151968 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 152288 171978
rect 151968 171888 152288 171922
rect 182688 172350 183008 172384
rect 182688 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 183008 172350
rect 182688 172226 183008 172294
rect 182688 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 183008 172226
rect 182688 172102 183008 172170
rect 182688 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 183008 172102
rect 182688 171978 183008 172046
rect 182688 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 183008 171978
rect 182688 171888 183008 171922
rect 213408 172350 213728 172384
rect 213408 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 213728 172350
rect 213408 172226 213728 172294
rect 213408 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 213728 172226
rect 213408 172102 213728 172170
rect 213408 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 213728 172102
rect 213408 171978 213728 172046
rect 213408 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 213728 171978
rect 213408 171888 213728 171922
rect 244128 172350 244448 172384
rect 244128 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 244448 172350
rect 244128 172226 244448 172294
rect 244128 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 244448 172226
rect 244128 172102 244448 172170
rect 244128 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 244448 172102
rect 244128 171978 244448 172046
rect 244128 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 244448 171978
rect 244128 171888 244448 171922
rect 44448 166350 44768 166384
rect 44448 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 44768 166350
rect 44448 166226 44768 166294
rect 44448 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 44768 166226
rect 44448 166102 44768 166170
rect 44448 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 44768 166102
rect 44448 165978 44768 166046
rect 44448 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 44768 165978
rect 44448 165888 44768 165922
rect 75168 166350 75488 166384
rect 75168 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 75488 166350
rect 75168 166226 75488 166294
rect 75168 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 75488 166226
rect 75168 166102 75488 166170
rect 75168 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 75488 166102
rect 75168 165978 75488 166046
rect 75168 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 75488 165978
rect 75168 165888 75488 165922
rect 105888 166350 106208 166384
rect 105888 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 106208 166350
rect 105888 166226 106208 166294
rect 105888 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 106208 166226
rect 105888 166102 106208 166170
rect 105888 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 106208 166102
rect 105888 165978 106208 166046
rect 105888 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 106208 165978
rect 105888 165888 106208 165922
rect 136608 166350 136928 166384
rect 136608 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 136928 166350
rect 136608 166226 136928 166294
rect 136608 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 136928 166226
rect 136608 166102 136928 166170
rect 136608 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 136928 166102
rect 136608 165978 136928 166046
rect 136608 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 136928 165978
rect 136608 165888 136928 165922
rect 167328 166350 167648 166384
rect 167328 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 167648 166350
rect 167328 166226 167648 166294
rect 167328 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 167648 166226
rect 167328 166102 167648 166170
rect 167328 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 167648 166102
rect 167328 165978 167648 166046
rect 167328 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 167648 165978
rect 167328 165888 167648 165922
rect 198048 166350 198368 166384
rect 198048 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 198368 166350
rect 198048 166226 198368 166294
rect 198048 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 198368 166226
rect 198048 166102 198368 166170
rect 198048 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 198368 166102
rect 198048 165978 198368 166046
rect 198048 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 198368 165978
rect 198048 165888 198368 165922
rect 228768 166350 229088 166384
rect 228768 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 229088 166350
rect 228768 166226 229088 166294
rect 228768 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 229088 166226
rect 228768 166102 229088 166170
rect 228768 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 229088 166102
rect 228768 165978 229088 166046
rect 228768 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 229088 165978
rect 228768 165888 229088 165922
rect 259488 166350 259808 166384
rect 259488 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 259808 166350
rect 259488 166226 259808 166294
rect 259488 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 259808 166226
rect 259488 166102 259808 166170
rect 259488 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 259808 166102
rect 259488 165978 259808 166046
rect 259488 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 259808 165978
rect 259488 165888 259808 165922
rect 59808 154350 60128 154384
rect 59808 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 60128 154350
rect 59808 154226 60128 154294
rect 59808 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 60128 154226
rect 59808 154102 60128 154170
rect 59808 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 60128 154102
rect 59808 153978 60128 154046
rect 59808 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 60128 153978
rect 59808 153888 60128 153922
rect 90528 154350 90848 154384
rect 90528 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 90848 154350
rect 90528 154226 90848 154294
rect 90528 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 90848 154226
rect 90528 154102 90848 154170
rect 90528 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 90848 154102
rect 90528 153978 90848 154046
rect 90528 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 90848 153978
rect 90528 153888 90848 153922
rect 121248 154350 121568 154384
rect 121248 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 121568 154350
rect 121248 154226 121568 154294
rect 121248 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 121568 154226
rect 121248 154102 121568 154170
rect 121248 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 121568 154102
rect 121248 153978 121568 154046
rect 121248 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 121568 153978
rect 121248 153888 121568 153922
rect 151968 154350 152288 154384
rect 151968 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 152288 154350
rect 151968 154226 152288 154294
rect 151968 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 152288 154226
rect 151968 154102 152288 154170
rect 151968 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 152288 154102
rect 151968 153978 152288 154046
rect 151968 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 152288 153978
rect 151968 153888 152288 153922
rect 182688 154350 183008 154384
rect 182688 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 183008 154350
rect 182688 154226 183008 154294
rect 182688 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 183008 154226
rect 182688 154102 183008 154170
rect 182688 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 183008 154102
rect 182688 153978 183008 154046
rect 182688 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 183008 153978
rect 182688 153888 183008 153922
rect 213408 154350 213728 154384
rect 213408 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 213728 154350
rect 213408 154226 213728 154294
rect 213408 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 213728 154226
rect 213408 154102 213728 154170
rect 213408 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 213728 154102
rect 213408 153978 213728 154046
rect 213408 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 213728 153978
rect 213408 153888 213728 153922
rect 244128 154350 244448 154384
rect 244128 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 244448 154350
rect 244128 154226 244448 154294
rect 244128 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 244448 154226
rect 244128 154102 244448 154170
rect 244128 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 244448 154102
rect 244128 153978 244448 154046
rect 244128 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 244448 153978
rect 244128 153888 244448 153922
rect 44448 148350 44768 148384
rect 44448 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 44768 148350
rect 44448 148226 44768 148294
rect 44448 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 44768 148226
rect 44448 148102 44768 148170
rect 44448 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 44768 148102
rect 44448 147978 44768 148046
rect 44448 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 44768 147978
rect 44448 147888 44768 147922
rect 75168 148350 75488 148384
rect 75168 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 75488 148350
rect 75168 148226 75488 148294
rect 75168 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 75488 148226
rect 75168 148102 75488 148170
rect 75168 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 75488 148102
rect 75168 147978 75488 148046
rect 75168 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 75488 147978
rect 75168 147888 75488 147922
rect 105888 148350 106208 148384
rect 105888 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 106208 148350
rect 105888 148226 106208 148294
rect 105888 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 106208 148226
rect 105888 148102 106208 148170
rect 105888 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 106208 148102
rect 105888 147978 106208 148046
rect 105888 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 106208 147978
rect 105888 147888 106208 147922
rect 136608 148350 136928 148384
rect 136608 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 136928 148350
rect 136608 148226 136928 148294
rect 136608 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 136928 148226
rect 136608 148102 136928 148170
rect 136608 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 136928 148102
rect 136608 147978 136928 148046
rect 136608 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 136928 147978
rect 136608 147888 136928 147922
rect 167328 148350 167648 148384
rect 167328 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 167648 148350
rect 167328 148226 167648 148294
rect 167328 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 167648 148226
rect 167328 148102 167648 148170
rect 167328 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 167648 148102
rect 167328 147978 167648 148046
rect 167328 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 167648 147978
rect 167328 147888 167648 147922
rect 198048 148350 198368 148384
rect 198048 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 198368 148350
rect 198048 148226 198368 148294
rect 198048 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 198368 148226
rect 198048 148102 198368 148170
rect 198048 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 198368 148102
rect 198048 147978 198368 148046
rect 198048 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 198368 147978
rect 198048 147888 198368 147922
rect 228768 148350 229088 148384
rect 228768 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 229088 148350
rect 228768 148226 229088 148294
rect 228768 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 229088 148226
rect 228768 148102 229088 148170
rect 228768 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 229088 148102
rect 228768 147978 229088 148046
rect 228768 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 229088 147978
rect 228768 147888 229088 147922
rect 259488 148350 259808 148384
rect 259488 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 259808 148350
rect 259488 148226 259808 148294
rect 259488 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 259808 148226
rect 259488 148102 259808 148170
rect 259488 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 259808 148102
rect 259488 147978 259808 148046
rect 259488 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 259808 147978
rect 259488 147888 259808 147922
rect 59808 136350 60128 136384
rect 59808 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 60128 136350
rect 59808 136226 60128 136294
rect 59808 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 60128 136226
rect 59808 136102 60128 136170
rect 59808 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 60128 136102
rect 59808 135978 60128 136046
rect 59808 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 60128 135978
rect 59808 135888 60128 135922
rect 90528 136350 90848 136384
rect 90528 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 90848 136350
rect 90528 136226 90848 136294
rect 90528 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 90848 136226
rect 90528 136102 90848 136170
rect 90528 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 90848 136102
rect 90528 135978 90848 136046
rect 90528 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 90848 135978
rect 90528 135888 90848 135922
rect 121248 136350 121568 136384
rect 121248 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 121568 136350
rect 121248 136226 121568 136294
rect 121248 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 121568 136226
rect 121248 136102 121568 136170
rect 121248 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 121568 136102
rect 121248 135978 121568 136046
rect 121248 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 121568 135978
rect 121248 135888 121568 135922
rect 151968 136350 152288 136384
rect 151968 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 152288 136350
rect 151968 136226 152288 136294
rect 151968 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 152288 136226
rect 151968 136102 152288 136170
rect 151968 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 152288 136102
rect 151968 135978 152288 136046
rect 151968 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 152288 135978
rect 151968 135888 152288 135922
rect 182688 136350 183008 136384
rect 182688 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 183008 136350
rect 182688 136226 183008 136294
rect 182688 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 183008 136226
rect 182688 136102 183008 136170
rect 182688 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 183008 136102
rect 182688 135978 183008 136046
rect 182688 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 183008 135978
rect 182688 135888 183008 135922
rect 213408 136350 213728 136384
rect 213408 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 213728 136350
rect 213408 136226 213728 136294
rect 213408 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 213728 136226
rect 213408 136102 213728 136170
rect 213408 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 213728 136102
rect 213408 135978 213728 136046
rect 213408 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 213728 135978
rect 213408 135888 213728 135922
rect 244128 136350 244448 136384
rect 244128 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 244448 136350
rect 244128 136226 244448 136294
rect 244128 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 244448 136226
rect 244128 136102 244448 136170
rect 244128 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 244448 136102
rect 244128 135978 244448 136046
rect 244128 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 244448 135978
rect 244128 135888 244448 135922
rect 44448 130350 44768 130384
rect 44448 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 44768 130350
rect 44448 130226 44768 130294
rect 44448 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 44768 130226
rect 44448 130102 44768 130170
rect 44448 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 44768 130102
rect 44448 129978 44768 130046
rect 44448 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 44768 129978
rect 44448 129888 44768 129922
rect 75168 130350 75488 130384
rect 75168 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 75488 130350
rect 75168 130226 75488 130294
rect 75168 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 75488 130226
rect 75168 130102 75488 130170
rect 75168 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 75488 130102
rect 75168 129978 75488 130046
rect 75168 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 75488 129978
rect 75168 129888 75488 129922
rect 105888 130350 106208 130384
rect 105888 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 106208 130350
rect 105888 130226 106208 130294
rect 105888 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 106208 130226
rect 105888 130102 106208 130170
rect 105888 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 106208 130102
rect 105888 129978 106208 130046
rect 105888 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 106208 129978
rect 105888 129888 106208 129922
rect 136608 130350 136928 130384
rect 136608 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 136928 130350
rect 136608 130226 136928 130294
rect 136608 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 136928 130226
rect 136608 130102 136928 130170
rect 136608 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 136928 130102
rect 136608 129978 136928 130046
rect 136608 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 136928 129978
rect 136608 129888 136928 129922
rect 167328 130350 167648 130384
rect 167328 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 167648 130350
rect 167328 130226 167648 130294
rect 167328 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 167648 130226
rect 167328 130102 167648 130170
rect 167328 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 167648 130102
rect 167328 129978 167648 130046
rect 167328 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 167648 129978
rect 167328 129888 167648 129922
rect 198048 130350 198368 130384
rect 198048 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 198368 130350
rect 198048 130226 198368 130294
rect 198048 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 198368 130226
rect 198048 130102 198368 130170
rect 198048 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 198368 130102
rect 198048 129978 198368 130046
rect 198048 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 198368 129978
rect 198048 129888 198368 129922
rect 228768 130350 229088 130384
rect 228768 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 229088 130350
rect 228768 130226 229088 130294
rect 228768 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 229088 130226
rect 228768 130102 229088 130170
rect 228768 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 229088 130102
rect 228768 129978 229088 130046
rect 228768 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 229088 129978
rect 228768 129888 229088 129922
rect 259488 130350 259808 130384
rect 259488 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 259808 130350
rect 259488 130226 259808 130294
rect 259488 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 259808 130226
rect 259488 130102 259808 130170
rect 259488 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 259808 130102
rect 259488 129978 259808 130046
rect 259488 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 259808 129978
rect 259488 129888 259808 129922
rect 59808 118350 60128 118384
rect 59808 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 60128 118350
rect 59808 118226 60128 118294
rect 59808 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 60128 118226
rect 59808 118102 60128 118170
rect 59808 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 60128 118102
rect 59808 117978 60128 118046
rect 59808 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 60128 117978
rect 59808 117888 60128 117922
rect 90528 118350 90848 118384
rect 90528 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 90848 118350
rect 90528 118226 90848 118294
rect 90528 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 90848 118226
rect 90528 118102 90848 118170
rect 90528 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 90848 118102
rect 90528 117978 90848 118046
rect 90528 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 90848 117978
rect 90528 117888 90848 117922
rect 121248 118350 121568 118384
rect 121248 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 121568 118350
rect 121248 118226 121568 118294
rect 121248 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 121568 118226
rect 121248 118102 121568 118170
rect 121248 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 121568 118102
rect 121248 117978 121568 118046
rect 121248 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 121568 117978
rect 121248 117888 121568 117922
rect 151968 118350 152288 118384
rect 151968 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 152288 118350
rect 151968 118226 152288 118294
rect 151968 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 152288 118226
rect 151968 118102 152288 118170
rect 151968 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 152288 118102
rect 151968 117978 152288 118046
rect 151968 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 152288 117978
rect 151968 117888 152288 117922
rect 182688 118350 183008 118384
rect 182688 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 183008 118350
rect 182688 118226 183008 118294
rect 182688 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 183008 118226
rect 182688 118102 183008 118170
rect 182688 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 183008 118102
rect 182688 117978 183008 118046
rect 182688 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 183008 117978
rect 182688 117888 183008 117922
rect 213408 118350 213728 118384
rect 213408 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 213728 118350
rect 213408 118226 213728 118294
rect 213408 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 213728 118226
rect 213408 118102 213728 118170
rect 213408 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 213728 118102
rect 213408 117978 213728 118046
rect 213408 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 213728 117978
rect 213408 117888 213728 117922
rect 244128 118350 244448 118384
rect 244128 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 244448 118350
rect 244128 118226 244448 118294
rect 244128 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 244448 118226
rect 244128 118102 244448 118170
rect 244128 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 244448 118102
rect 244128 117978 244448 118046
rect 244128 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 244448 117978
rect 244128 117888 244448 117922
rect 44448 112350 44768 112384
rect 44448 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 44768 112350
rect 44448 112226 44768 112294
rect 44448 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 44768 112226
rect 44448 112102 44768 112170
rect 44448 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 44768 112102
rect 44448 111978 44768 112046
rect 44448 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 44768 111978
rect 44448 111888 44768 111922
rect 75168 112350 75488 112384
rect 75168 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 75488 112350
rect 75168 112226 75488 112294
rect 75168 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 75488 112226
rect 75168 112102 75488 112170
rect 75168 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 75488 112102
rect 75168 111978 75488 112046
rect 75168 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 75488 111978
rect 75168 111888 75488 111922
rect 105888 112350 106208 112384
rect 105888 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 106208 112350
rect 105888 112226 106208 112294
rect 105888 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 106208 112226
rect 105888 112102 106208 112170
rect 105888 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 106208 112102
rect 105888 111978 106208 112046
rect 105888 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 106208 111978
rect 105888 111888 106208 111922
rect 136608 112350 136928 112384
rect 136608 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 136928 112350
rect 136608 112226 136928 112294
rect 136608 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 136928 112226
rect 136608 112102 136928 112170
rect 136608 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 136928 112102
rect 136608 111978 136928 112046
rect 136608 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 136928 111978
rect 136608 111888 136928 111922
rect 167328 112350 167648 112384
rect 167328 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 167648 112350
rect 167328 112226 167648 112294
rect 167328 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 167648 112226
rect 167328 112102 167648 112170
rect 167328 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 167648 112102
rect 167328 111978 167648 112046
rect 167328 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 167648 111978
rect 167328 111888 167648 111922
rect 198048 112350 198368 112384
rect 198048 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 198368 112350
rect 198048 112226 198368 112294
rect 198048 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 198368 112226
rect 198048 112102 198368 112170
rect 198048 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 198368 112102
rect 198048 111978 198368 112046
rect 198048 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 198368 111978
rect 198048 111888 198368 111922
rect 228768 112350 229088 112384
rect 228768 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 229088 112350
rect 228768 112226 229088 112294
rect 228768 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 229088 112226
rect 228768 112102 229088 112170
rect 228768 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 229088 112102
rect 228768 111978 229088 112046
rect 228768 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 229088 111978
rect 228768 111888 229088 111922
rect 259488 112350 259808 112384
rect 259488 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 259808 112350
rect 259488 112226 259808 112294
rect 259488 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 259808 112226
rect 259488 112102 259808 112170
rect 259488 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 259808 112102
rect 259488 111978 259808 112046
rect 259488 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 259808 111978
rect 259488 111888 259808 111922
rect 59808 100350 60128 100384
rect 59808 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 60128 100350
rect 59808 100226 60128 100294
rect 59808 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 60128 100226
rect 59808 100102 60128 100170
rect 59808 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 60128 100102
rect 59808 99978 60128 100046
rect 59808 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 60128 99978
rect 59808 99888 60128 99922
rect 90528 100350 90848 100384
rect 90528 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 90848 100350
rect 90528 100226 90848 100294
rect 90528 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 90848 100226
rect 90528 100102 90848 100170
rect 90528 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 90848 100102
rect 90528 99978 90848 100046
rect 90528 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 90848 99978
rect 90528 99888 90848 99922
rect 121248 100350 121568 100384
rect 121248 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 121568 100350
rect 121248 100226 121568 100294
rect 121248 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 121568 100226
rect 121248 100102 121568 100170
rect 121248 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 121568 100102
rect 121248 99978 121568 100046
rect 121248 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 121568 99978
rect 121248 99888 121568 99922
rect 151968 100350 152288 100384
rect 151968 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 152288 100350
rect 151968 100226 152288 100294
rect 151968 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 152288 100226
rect 151968 100102 152288 100170
rect 151968 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 152288 100102
rect 151968 99978 152288 100046
rect 151968 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 152288 99978
rect 151968 99888 152288 99922
rect 182688 100350 183008 100384
rect 182688 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 183008 100350
rect 182688 100226 183008 100294
rect 182688 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 183008 100226
rect 182688 100102 183008 100170
rect 182688 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 183008 100102
rect 182688 99978 183008 100046
rect 182688 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 183008 99978
rect 182688 99888 183008 99922
rect 213408 100350 213728 100384
rect 213408 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 213728 100350
rect 213408 100226 213728 100294
rect 213408 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 213728 100226
rect 213408 100102 213728 100170
rect 213408 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 213728 100102
rect 213408 99978 213728 100046
rect 213408 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 213728 99978
rect 213408 99888 213728 99922
rect 244128 100350 244448 100384
rect 244128 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 244448 100350
rect 244128 100226 244448 100294
rect 244128 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 244448 100226
rect 244128 100102 244448 100170
rect 244128 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 244448 100102
rect 244128 99978 244448 100046
rect 244128 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 244448 99978
rect 244128 99888 244448 99922
rect 44448 94350 44768 94384
rect 44448 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 44768 94350
rect 44448 94226 44768 94294
rect 44448 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 44768 94226
rect 44448 94102 44768 94170
rect 44448 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 44768 94102
rect 44448 93978 44768 94046
rect 44448 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 44768 93978
rect 44448 93888 44768 93922
rect 75168 94350 75488 94384
rect 75168 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 75488 94350
rect 75168 94226 75488 94294
rect 75168 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 75488 94226
rect 75168 94102 75488 94170
rect 75168 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 75488 94102
rect 75168 93978 75488 94046
rect 75168 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 75488 93978
rect 75168 93888 75488 93922
rect 105888 94350 106208 94384
rect 105888 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 106208 94350
rect 105888 94226 106208 94294
rect 105888 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 106208 94226
rect 105888 94102 106208 94170
rect 105888 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 106208 94102
rect 105888 93978 106208 94046
rect 105888 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 106208 93978
rect 105888 93888 106208 93922
rect 136608 94350 136928 94384
rect 136608 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 136928 94350
rect 136608 94226 136928 94294
rect 136608 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 136928 94226
rect 136608 94102 136928 94170
rect 136608 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 136928 94102
rect 136608 93978 136928 94046
rect 136608 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 136928 93978
rect 136608 93888 136928 93922
rect 167328 94350 167648 94384
rect 167328 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 167648 94350
rect 167328 94226 167648 94294
rect 167328 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 167648 94226
rect 167328 94102 167648 94170
rect 167328 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 167648 94102
rect 167328 93978 167648 94046
rect 167328 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 167648 93978
rect 167328 93888 167648 93922
rect 198048 94350 198368 94384
rect 198048 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 198368 94350
rect 198048 94226 198368 94294
rect 198048 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 198368 94226
rect 198048 94102 198368 94170
rect 198048 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 198368 94102
rect 198048 93978 198368 94046
rect 198048 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 198368 93978
rect 198048 93888 198368 93922
rect 228768 94350 229088 94384
rect 228768 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 229088 94350
rect 228768 94226 229088 94294
rect 228768 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 229088 94226
rect 228768 94102 229088 94170
rect 228768 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 229088 94102
rect 228768 93978 229088 94046
rect 228768 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 229088 93978
rect 228768 93888 229088 93922
rect 259488 94350 259808 94384
rect 259488 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 259808 94350
rect 259488 94226 259808 94294
rect 259488 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 259808 94226
rect 259488 94102 259808 94170
rect 259488 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 259808 94102
rect 259488 93978 259808 94046
rect 259488 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 259808 93978
rect 259488 93888 259808 93922
rect 59808 82350 60128 82384
rect 59808 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 60128 82350
rect 59808 82226 60128 82294
rect 59808 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 60128 82226
rect 59808 82102 60128 82170
rect 59808 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 60128 82102
rect 59808 81978 60128 82046
rect 59808 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 60128 81978
rect 59808 81888 60128 81922
rect 90528 82350 90848 82384
rect 90528 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 90848 82350
rect 90528 82226 90848 82294
rect 90528 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 90848 82226
rect 90528 82102 90848 82170
rect 90528 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 90848 82102
rect 90528 81978 90848 82046
rect 90528 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 90848 81978
rect 90528 81888 90848 81922
rect 121248 82350 121568 82384
rect 121248 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 121568 82350
rect 121248 82226 121568 82294
rect 121248 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 121568 82226
rect 121248 82102 121568 82170
rect 121248 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 121568 82102
rect 121248 81978 121568 82046
rect 121248 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 121568 81978
rect 121248 81888 121568 81922
rect 151968 82350 152288 82384
rect 151968 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 152288 82350
rect 151968 82226 152288 82294
rect 151968 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 152288 82226
rect 151968 82102 152288 82170
rect 151968 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 152288 82102
rect 151968 81978 152288 82046
rect 151968 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 152288 81978
rect 151968 81888 152288 81922
rect 182688 82350 183008 82384
rect 182688 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 183008 82350
rect 182688 82226 183008 82294
rect 182688 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 183008 82226
rect 182688 82102 183008 82170
rect 182688 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 183008 82102
rect 182688 81978 183008 82046
rect 182688 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 183008 81978
rect 182688 81888 183008 81922
rect 213408 82350 213728 82384
rect 213408 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 213728 82350
rect 213408 82226 213728 82294
rect 213408 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 213728 82226
rect 213408 82102 213728 82170
rect 213408 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 213728 82102
rect 213408 81978 213728 82046
rect 213408 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 213728 81978
rect 213408 81888 213728 81922
rect 244128 82350 244448 82384
rect 244128 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 244448 82350
rect 244128 82226 244448 82294
rect 244128 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 244448 82226
rect 244128 82102 244448 82170
rect 244128 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 244448 82102
rect 244128 81978 244448 82046
rect 244128 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 244448 81978
rect 244128 81888 244448 81922
rect 44448 76350 44768 76384
rect 44448 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 44768 76350
rect 44448 76226 44768 76294
rect 44448 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 44768 76226
rect 44448 76102 44768 76170
rect 44448 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 44768 76102
rect 44448 75978 44768 76046
rect 44448 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 44768 75978
rect 44448 75888 44768 75922
rect 75168 76350 75488 76384
rect 75168 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 75488 76350
rect 75168 76226 75488 76294
rect 75168 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 75488 76226
rect 75168 76102 75488 76170
rect 75168 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 75488 76102
rect 75168 75978 75488 76046
rect 75168 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 75488 75978
rect 75168 75888 75488 75922
rect 105888 76350 106208 76384
rect 105888 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 106208 76350
rect 105888 76226 106208 76294
rect 105888 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 106208 76226
rect 105888 76102 106208 76170
rect 105888 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 106208 76102
rect 105888 75978 106208 76046
rect 105888 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 106208 75978
rect 105888 75888 106208 75922
rect 136608 76350 136928 76384
rect 136608 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 136928 76350
rect 136608 76226 136928 76294
rect 136608 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 136928 76226
rect 136608 76102 136928 76170
rect 136608 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 136928 76102
rect 136608 75978 136928 76046
rect 136608 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 136928 75978
rect 136608 75888 136928 75922
rect 167328 76350 167648 76384
rect 167328 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 167648 76350
rect 167328 76226 167648 76294
rect 167328 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 167648 76226
rect 167328 76102 167648 76170
rect 167328 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 167648 76102
rect 167328 75978 167648 76046
rect 167328 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 167648 75978
rect 167328 75888 167648 75922
rect 198048 76350 198368 76384
rect 198048 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 198368 76350
rect 198048 76226 198368 76294
rect 198048 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 198368 76226
rect 198048 76102 198368 76170
rect 198048 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 198368 76102
rect 198048 75978 198368 76046
rect 198048 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 198368 75978
rect 198048 75888 198368 75922
rect 228768 76350 229088 76384
rect 228768 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 229088 76350
rect 228768 76226 229088 76294
rect 228768 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 229088 76226
rect 228768 76102 229088 76170
rect 228768 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 229088 76102
rect 228768 75978 229088 76046
rect 228768 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 229088 75978
rect 228768 75888 229088 75922
rect 259488 76350 259808 76384
rect 259488 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 259808 76350
rect 259488 76226 259808 76294
rect 259488 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 259808 76226
rect 259488 76102 259808 76170
rect 259488 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 259808 76102
rect 259488 75978 259808 76046
rect 259488 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 259808 75978
rect 259488 75888 259808 75922
rect 59808 64350 60128 64384
rect 59808 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 60128 64350
rect 59808 64226 60128 64294
rect 59808 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 60128 64226
rect 59808 64102 60128 64170
rect 59808 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 60128 64102
rect 59808 63978 60128 64046
rect 59808 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 60128 63978
rect 59808 63888 60128 63922
rect 90528 64350 90848 64384
rect 90528 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 90848 64350
rect 90528 64226 90848 64294
rect 90528 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 90848 64226
rect 90528 64102 90848 64170
rect 90528 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 90848 64102
rect 90528 63978 90848 64046
rect 90528 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 90848 63978
rect 90528 63888 90848 63922
rect 121248 64350 121568 64384
rect 121248 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 121568 64350
rect 121248 64226 121568 64294
rect 121248 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 121568 64226
rect 121248 64102 121568 64170
rect 121248 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 121568 64102
rect 121248 63978 121568 64046
rect 121248 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 121568 63978
rect 121248 63888 121568 63922
rect 151968 64350 152288 64384
rect 151968 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 152288 64350
rect 151968 64226 152288 64294
rect 151968 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 152288 64226
rect 151968 64102 152288 64170
rect 151968 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 152288 64102
rect 151968 63978 152288 64046
rect 151968 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 152288 63978
rect 151968 63888 152288 63922
rect 182688 64350 183008 64384
rect 182688 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 183008 64350
rect 182688 64226 183008 64294
rect 182688 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 183008 64226
rect 182688 64102 183008 64170
rect 182688 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 183008 64102
rect 182688 63978 183008 64046
rect 182688 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 183008 63978
rect 182688 63888 183008 63922
rect 213408 64350 213728 64384
rect 213408 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 213728 64350
rect 213408 64226 213728 64294
rect 213408 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 213728 64226
rect 213408 64102 213728 64170
rect 213408 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 213728 64102
rect 213408 63978 213728 64046
rect 213408 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 213728 63978
rect 213408 63888 213728 63922
rect 244128 64350 244448 64384
rect 244128 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 244448 64350
rect 244128 64226 244448 64294
rect 244128 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 244448 64226
rect 244128 64102 244448 64170
rect 244128 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 244448 64102
rect 244128 63978 244448 64046
rect 244128 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 244448 63978
rect 244128 63888 244448 63922
rect 44448 58350 44768 58384
rect 44448 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 44768 58350
rect 44448 58226 44768 58294
rect 44448 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 44768 58226
rect 44448 58102 44768 58170
rect 44448 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 44768 58102
rect 44448 57978 44768 58046
rect 44448 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 44768 57978
rect 44448 57888 44768 57922
rect 75168 58350 75488 58384
rect 75168 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 75488 58350
rect 75168 58226 75488 58294
rect 75168 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 75488 58226
rect 75168 58102 75488 58170
rect 75168 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 75488 58102
rect 75168 57978 75488 58046
rect 75168 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 75488 57978
rect 75168 57888 75488 57922
rect 105888 58350 106208 58384
rect 105888 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 106208 58350
rect 105888 58226 106208 58294
rect 105888 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 106208 58226
rect 105888 58102 106208 58170
rect 105888 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 106208 58102
rect 105888 57978 106208 58046
rect 105888 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 106208 57978
rect 105888 57888 106208 57922
rect 136608 58350 136928 58384
rect 136608 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 136928 58350
rect 136608 58226 136928 58294
rect 136608 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 136928 58226
rect 136608 58102 136928 58170
rect 136608 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 136928 58102
rect 136608 57978 136928 58046
rect 136608 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 136928 57978
rect 136608 57888 136928 57922
rect 167328 58350 167648 58384
rect 167328 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 167648 58350
rect 167328 58226 167648 58294
rect 167328 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 167648 58226
rect 167328 58102 167648 58170
rect 167328 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 167648 58102
rect 167328 57978 167648 58046
rect 167328 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 167648 57978
rect 167328 57888 167648 57922
rect 198048 58350 198368 58384
rect 198048 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 198368 58350
rect 198048 58226 198368 58294
rect 198048 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 198368 58226
rect 198048 58102 198368 58170
rect 198048 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 198368 58102
rect 198048 57978 198368 58046
rect 198048 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 198368 57978
rect 198048 57888 198368 57922
rect 228768 58350 229088 58384
rect 228768 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 229088 58350
rect 228768 58226 229088 58294
rect 228768 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 229088 58226
rect 228768 58102 229088 58170
rect 228768 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 229088 58102
rect 228768 57978 229088 58046
rect 228768 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 229088 57978
rect 228768 57888 229088 57922
rect 259488 58350 259808 58384
rect 259488 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 259808 58350
rect 259488 58226 259808 58294
rect 259488 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 259808 58226
rect 259488 58102 259808 58170
rect 259488 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 259808 58102
rect 259488 57978 259808 58046
rect 259488 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 259808 57978
rect 259488 57888 259808 57922
rect 45612 50820 45668 50830
rect 45612 50372 45668 50764
rect 45612 50306 45668 50316
rect 41916 4386 41972 4396
rect 66858 40350 67478 53002
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 46350 71198 53002
rect 87500 51268 87556 51278
rect 87500 50596 87556 51212
rect 87500 50530 87556 50540
rect 89404 51268 89460 51278
rect 89404 50596 89460 51212
rect 89404 50530 89460 50540
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 70578 28350 71198 45922
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 40350 98198 53002
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 97578 22350 98198 39922
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 46350 101918 53002
rect 101298 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 101918 46350
rect 101298 46226 101918 46294
rect 101298 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 101918 46226
rect 101298 46102 101918 46170
rect 101298 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 101918 46102
rect 101298 45978 101918 46046
rect 101298 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 101918 45978
rect 101298 28350 101918 45922
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 40350 128918 53002
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 128298 22350 128918 39922
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 128298 4350 128918 21922
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 46350 132638 53002
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 132018 10350 132638 27922
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 40350 159638 53002
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 159018 4350 159638 21922
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 46350 163358 53002
rect 173180 51380 173236 51390
rect 173180 50596 173236 51324
rect 173180 50530 173236 50540
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 40350 190358 53002
rect 190428 51492 190484 51502
rect 190428 50372 190484 51436
rect 190428 50306 190484 50316
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 189738 4350 190358 21922
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 46350 194078 53002
rect 209356 51828 209412 51838
rect 201740 51716 201796 51726
rect 196028 51604 196084 51614
rect 196028 50372 196084 51548
rect 196028 50306 196084 50316
rect 201740 50372 201796 51660
rect 201740 50306 201796 50316
rect 209356 50372 209412 51772
rect 209356 50306 209412 50316
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 193458 10350 194078 27922
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 193458 -1120 194078 9922
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 40350 221078 53002
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 46350 224798 53002
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 40350 251798 53002
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 251178 4350 251798 21922
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 46350 255518 53002
rect 266924 51268 266980 235004
rect 267036 204958 267092 236908
rect 267036 204892 267092 204902
rect 266924 51202 266980 51212
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 254898 28350 255518 45922
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 254898 -1120 255518 9922
rect 267148 7588 267204 237122
rect 267372 236998 267428 237008
rect 267260 235172 267316 235182
rect 267260 42868 267316 235116
rect 267372 49812 267428 236942
rect 267484 231812 267540 231822
rect 267484 51380 267540 231756
rect 267708 211428 267764 211438
rect 267708 210980 267764 211372
rect 267708 210914 267764 210924
rect 267932 211316 267988 211326
rect 267932 210756 267988 211260
rect 267932 210690 267988 210700
rect 267932 205858 267988 205868
rect 267484 51314 267540 51324
rect 267596 204058 267652 204068
rect 267372 49746 267428 49756
rect 267596 46228 267652 204002
rect 267932 143398 267988 205802
rect 268044 201538 268100 239708
rect 275660 239652 275716 239662
rect 268828 238084 268884 238094
rect 268716 237076 268772 237086
rect 268044 201472 268100 201482
rect 268604 236964 268660 236974
rect 267932 143332 267988 143342
rect 268604 115138 268660 236908
rect 268716 115318 268772 237020
rect 268716 115252 268772 115262
rect 268604 115072 268660 115082
rect 267596 46162 267652 46172
rect 267260 42802 267316 42812
rect 268828 9268 268884 238028
rect 270396 237076 270452 237086
rect 270284 236964 270340 236974
rect 269500 233268 269556 233278
rect 268940 231028 268996 231038
rect 268940 42980 268996 230972
rect 269052 227556 269108 227566
rect 269052 43204 269108 227500
rect 269500 195412 269556 233212
rect 269612 209076 269668 209086
rect 269612 204820 269668 209020
rect 269612 204754 269668 204764
rect 269724 206578 269780 206588
rect 269612 201538 269668 201548
rect 269612 201460 269668 201482
rect 269612 201394 269668 201404
rect 269500 195346 269556 195356
rect 269724 191548 269780 206522
rect 269612 191492 269780 191548
rect 269836 204958 269892 204968
rect 269612 109738 269668 191492
rect 269836 114268 269892 204902
rect 270284 145124 270340 236908
rect 270284 145058 270340 145068
rect 270396 142212 270452 237020
rect 275324 237076 275380 237086
rect 272076 236964 272132 236974
rect 270508 227668 270564 227678
rect 270508 203364 270564 227612
rect 271292 226548 271348 226558
rect 270620 224980 270676 224990
rect 270620 220078 270676 224924
rect 270620 220022 270900 220078
rect 270844 215068 270900 220022
rect 270620 215012 270900 215068
rect 270620 211708 270676 215012
rect 270620 211652 271012 211708
rect 270508 203298 270564 203308
rect 270732 203140 270788 203150
rect 270732 197578 270788 203084
rect 270956 199948 271012 211652
rect 270396 142146 270452 142156
rect 270508 197522 270788 197578
rect 270844 199892 271012 199948
rect 269836 114212 270116 114268
rect 269612 109682 270004 109738
rect 269948 105364 270004 109682
rect 269948 105298 270004 105308
rect 270060 105028 270116 114212
rect 270060 104962 270116 104972
rect 269052 43138 269108 43148
rect 268940 42914 268996 42924
rect 270508 39508 270564 197522
rect 270844 197218 270900 199892
rect 270620 197162 270900 197218
rect 270620 157556 270676 197162
rect 270620 157490 270676 157500
rect 270620 143668 270676 143678
rect 270620 55378 270676 143612
rect 270620 55312 270676 55322
rect 270508 39442 270564 39452
rect 268828 9202 268884 9212
rect 267148 7522 267204 7532
rect 271292 5908 271348 226492
rect 271404 222598 271460 222608
rect 271404 7588 271460 222542
rect 271516 216356 271572 216366
rect 271516 27972 271572 216300
rect 271740 214788 271796 214798
rect 271628 206218 271684 206228
rect 271628 113428 271684 206162
rect 271740 160692 271796 214732
rect 271852 206038 271908 206048
rect 271852 176372 271908 205982
rect 271852 176306 271908 176316
rect 271740 160626 271796 160636
rect 272076 149044 272132 236908
rect 272300 231588 272356 231598
rect 272300 209860 272356 231532
rect 273308 229908 273364 229918
rect 272300 209794 272356 209804
rect 272524 219940 272580 219950
rect 272412 209748 272468 209758
rect 272300 204238 272356 204248
rect 272188 203252 272244 203262
rect 272188 192500 272244 203196
rect 272188 192434 272244 192444
rect 272076 148978 272132 148988
rect 272188 143398 272244 143408
rect 272188 142858 272244 143342
rect 272188 137172 272244 142802
rect 272188 137106 272244 137116
rect 271628 113362 271684 113372
rect 272300 36148 272356 204182
rect 272412 198324 272468 209692
rect 272412 198258 272468 198268
rect 272524 186676 272580 219884
rect 273196 218260 273252 218270
rect 272524 186610 272580 186620
rect 272636 216468 272692 216478
rect 272300 36082 272356 36092
rect 272412 186452 272468 186462
rect 271516 27906 271572 27916
rect 272412 19348 272468 186396
rect 272636 177940 272692 216412
rect 272860 216244 272916 216254
rect 272748 209636 272804 209646
rect 272748 197578 272804 209580
rect 272860 203252 272916 216188
rect 273084 207478 273140 207488
rect 272972 206398 273028 206426
rect 272972 206322 273028 206332
rect 272860 203186 272916 203196
rect 272748 197522 273028 197578
rect 272748 197428 272804 197438
rect 272748 180852 272804 197372
rect 272748 180786 272804 180796
rect 272860 190708 272916 190718
rect 272636 177874 272692 177884
rect 272636 145908 272692 145918
rect 272636 36820 272692 145852
rect 272860 39732 272916 190652
rect 272972 189588 273028 197522
rect 272972 189522 273028 189532
rect 272972 143938 273028 143948
rect 272972 125524 273028 143882
rect 272972 125458 273028 125468
rect 272860 39666 272916 39676
rect 272636 36754 272692 36764
rect 273084 36372 273140 207422
rect 273196 183764 273252 218204
rect 273308 209188 273364 229852
rect 273980 226324 274036 226334
rect 273868 221284 273924 221294
rect 273308 209122 273364 209132
rect 273420 211092 273476 211102
rect 273420 197428 273476 211036
rect 273420 197362 273476 197372
rect 273756 199220 273812 199230
rect 273196 183698 273252 183708
rect 273644 178500 273700 178510
rect 273644 146132 273700 178444
rect 273644 145908 273700 146076
rect 273644 145842 273700 145852
rect 273196 143578 273252 143588
rect 273196 131348 273252 143522
rect 273756 143578 273812 199164
rect 273868 151732 273924 221228
rect 273980 172116 274036 226268
rect 274988 222964 275044 222974
rect 274764 212518 274820 212528
rect 273980 172050 274036 172060
rect 274652 211078 274708 211088
rect 273868 151666 273924 151676
rect 273756 143512 273812 143522
rect 273196 131282 273252 131292
rect 273084 36306 273140 36316
rect 272412 19282 272468 19292
rect 271404 7522 271460 7532
rect 274652 7140 274708 211022
rect 274764 20356 274820 212462
rect 274876 204418 274932 204428
rect 274876 110068 274932 204362
rect 274988 161218 275044 222908
rect 274988 161152 275044 161162
rect 275324 150724 275380 237020
rect 275324 150658 275380 150668
rect 275436 236964 275492 236974
rect 275436 150388 275492 236908
rect 275436 150322 275492 150332
rect 275548 209748 275604 209758
rect 274876 110002 274932 110012
rect 274988 132598 275044 132608
rect 274988 99316 275044 132542
rect 274988 99250 275044 99260
rect 275548 48356 275604 209692
rect 275660 160468 275716 239596
rect 278124 239652 278180 239662
rect 277116 236964 277172 236974
rect 276556 236628 276612 236638
rect 275660 160402 275716 160412
rect 275772 223412 275828 223422
rect 275772 154644 275828 223356
rect 276444 220052 276500 220062
rect 275772 154578 275828 154588
rect 276332 211798 276388 211808
rect 275548 48290 275604 48300
rect 276332 35218 276388 211742
rect 276444 84868 276500 219996
rect 276556 161038 276612 236572
rect 276556 160972 276612 160982
rect 277116 150500 277172 236908
rect 277116 150434 277172 150444
rect 278012 226436 278068 226446
rect 276444 84802 276500 84812
rect 276332 35152 276388 35162
rect 274764 20290 274820 20300
rect 278012 7700 278068 226380
rect 278124 45220 278180 239596
rect 278348 239540 278404 239550
rect 278236 214900 278292 214910
rect 278236 139438 278292 214844
rect 278236 139372 278292 139382
rect 278348 47796 278404 239484
rect 286412 239518 286468 239528
rect 281898 238350 282518 239082
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 278796 237076 278852 237086
rect 278684 236964 278740 236974
rect 278684 155764 278740 236908
rect 278684 155698 278740 155708
rect 278796 150612 278852 237020
rect 278796 150546 278852 150556
rect 279692 236098 279748 236108
rect 278348 47730 278404 47740
rect 278124 45154 278180 45164
rect 279692 37940 279748 236042
rect 280140 235060 280196 235070
rect 279804 232820 279860 232830
rect 279804 47908 279860 232764
rect 279804 47842 279860 47852
rect 279916 227668 279972 227678
rect 279916 44884 279972 227612
rect 280028 212884 280084 212894
rect 280028 48468 280084 212828
rect 280140 143758 280196 235004
rect 281484 231058 281540 231068
rect 280252 214676 280308 214686
rect 280252 160468 280308 214620
rect 280252 160402 280308 160412
rect 281372 211540 281428 211550
rect 280140 128436 280196 143702
rect 280140 128370 280196 128380
rect 280252 131878 280308 131888
rect 280252 102228 280308 131822
rect 281372 104158 281428 211484
rect 281484 158676 281540 231002
rect 281898 220350 282518 237922
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 281708 216580 281764 216590
rect 281484 158610 281540 158620
rect 281596 212660 281652 212670
rect 281596 153748 281652 212604
rect 281708 159598 281764 216524
rect 281708 159532 281764 159542
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281596 153682 281652 153692
rect 281372 104092 281428 104102
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 282604 236740 282660 236750
rect 282604 132598 282660 236684
rect 284732 234500 284788 234510
rect 283276 218148 283332 218158
rect 283164 215938 283220 215948
rect 282604 132532 282660 132542
rect 283052 212436 283108 212446
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 280252 102162 280308 102172
rect 280028 48402 280084 48412
rect 281898 94350 282518 111922
rect 283052 103978 283108 212380
rect 283164 150418 283220 215882
rect 283276 159460 283332 218092
rect 283276 159394 283332 159404
rect 283164 150352 283220 150362
rect 283052 103912 283108 103922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 281898 76350 282518 93922
rect 281898 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 282518 76350
rect 281898 76226 282518 76294
rect 281898 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 282518 76226
rect 281898 76102 282518 76170
rect 281898 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 282518 76102
rect 281898 75978 282518 76046
rect 281898 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 282518 75978
rect 281898 58350 282518 75922
rect 281898 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 282518 58350
rect 281898 58226 282518 58294
rect 281898 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 282518 58226
rect 281898 58102 282518 58170
rect 281898 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 282518 58102
rect 281898 57978 282518 58046
rect 281898 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 282518 57978
rect 279916 44818 279972 44828
rect 279692 37874 279748 37884
rect 281898 40350 282518 57922
rect 284732 41524 284788 234444
rect 284844 231028 284900 231038
rect 284844 48132 284900 230972
rect 284844 48066 284900 48076
rect 284956 229348 285012 229358
rect 284956 44660 285012 229292
rect 285618 226350 286238 239082
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285180 219178 285236 219188
rect 285068 214564 285124 214574
rect 285068 48356 285124 214508
rect 285180 134398 285236 219122
rect 285292 215012 285348 215022
rect 285292 152038 285348 214956
rect 285292 151972 285348 151982
rect 285618 208350 286238 225922
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285180 134332 285236 134342
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285068 48290 285124 48300
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 285618 82350 286238 99922
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 64350 286238 81922
rect 285618 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 286238 64350
rect 285618 64226 286238 64294
rect 285618 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 286238 64226
rect 285618 64102 286238 64170
rect 285618 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 286238 64102
rect 285618 63978 286238 64046
rect 285618 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 286238 63978
rect 284956 44594 285012 44604
rect 285618 46350 286238 63922
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 284732 41458 284788 41468
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 278012 7634 278068 7644
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 274652 7074 274708 7084
rect 271292 5842 271348 5852
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 4350 282518 21922
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 28350 286238 45922
rect 286412 41748 286468 239462
rect 288876 237748 288932 237758
rect 288092 236628 288148 236638
rect 286412 41682 286468 41692
rect 286636 231700 286692 231710
rect 286636 41412 286692 231644
rect 286636 41346 286692 41356
rect 288092 29428 288148 236572
rect 288428 233380 288484 233390
rect 288204 231812 288260 231822
rect 288204 37828 288260 231756
rect 288316 231058 288372 231068
rect 288316 41300 288372 231002
rect 288428 48244 288484 233324
rect 288652 216132 288708 216142
rect 288652 48580 288708 216076
rect 288876 147364 288932 237692
rect 293916 237076 293972 237086
rect 290556 236964 290612 236974
rect 289772 236740 289828 236750
rect 289660 234948 289716 234958
rect 289660 197652 289716 234892
rect 289660 197586 289716 197596
rect 288876 147298 288932 147308
rect 288652 48514 288708 48524
rect 288428 48178 288484 48188
rect 288316 41234 288372 41244
rect 289772 41188 289828 236684
rect 290108 235172 290164 235182
rect 289884 234948 289940 234958
rect 289884 44996 289940 234892
rect 289996 230916 290052 230926
rect 289996 49588 290052 230860
rect 289996 49522 290052 49532
rect 289884 44930 289940 44940
rect 290108 44772 290164 235116
rect 290444 199108 290500 199118
rect 290444 140308 290500 199052
rect 290444 140242 290500 140252
rect 290556 138516 290612 236908
rect 293804 236964 293860 236974
rect 291452 234612 291508 234622
rect 290668 221396 290724 221406
rect 290668 144478 290724 221340
rect 290846 184350 291166 184384
rect 290846 184294 290916 184350
rect 290972 184294 291040 184350
rect 291096 184294 291166 184350
rect 290846 184226 291166 184294
rect 290846 184170 290916 184226
rect 290972 184170 291040 184226
rect 291096 184170 291166 184226
rect 290846 184102 291166 184170
rect 290846 184046 290916 184102
rect 290972 184046 291040 184102
rect 291096 184046 291166 184102
rect 290846 183978 291166 184046
rect 290846 183922 290916 183978
rect 290972 183922 291040 183978
rect 291096 183922 291166 183978
rect 290846 183888 291166 183922
rect 290846 166350 291166 166384
rect 290846 166294 290916 166350
rect 290972 166294 291040 166350
rect 291096 166294 291166 166350
rect 290846 166226 291166 166294
rect 290846 166170 290916 166226
rect 290972 166170 291040 166226
rect 291096 166170 291166 166226
rect 290846 166102 291166 166170
rect 290846 166046 290916 166102
rect 290972 166046 291040 166102
rect 291096 166046 291166 166102
rect 290846 165978 291166 166046
rect 290846 165922 290916 165978
rect 290972 165922 291040 165978
rect 291096 165922 291166 165978
rect 290846 165888 291166 165922
rect 290668 144412 290724 144422
rect 290556 138450 290612 138460
rect 290108 44706 290164 44716
rect 291452 44548 291508 234556
rect 291564 233492 291620 233502
rect 291564 47684 291620 233436
rect 292348 224218 292404 224228
rect 292236 198884 292292 198894
rect 292236 152068 292292 198828
rect 292236 152002 292292 152012
rect 292348 132418 292404 224162
rect 293356 222852 293412 222862
rect 293244 218372 293300 218382
rect 293132 212772 293188 212782
rect 293132 154532 293188 212716
rect 293244 159348 293300 218316
rect 293356 169858 293412 222796
rect 293356 169792 293412 169802
rect 293692 199892 293748 199902
rect 293244 159282 293300 159292
rect 293132 154466 293188 154476
rect 293692 140420 293748 199836
rect 293804 153972 293860 236908
rect 293804 153906 293860 153916
rect 293916 145348 293972 237020
rect 293916 145282 293972 145292
rect 293692 140354 293748 140364
rect 292348 132352 292404 132362
rect 293132 134578 293188 134588
rect 293132 110964 293188 134522
rect 293132 110898 293188 110908
rect 294812 98308 294868 240380
rect 321804 239876 321860 239886
rect 321692 239338 321748 239348
rect 312618 238350 313238 239082
rect 295260 238308 295316 238318
rect 294924 234298 294980 234308
rect 294924 152758 294980 234242
rect 294924 152692 294980 152702
rect 295036 214138 295092 214148
rect 295036 98420 295092 214082
rect 295148 202804 295204 202814
rect 295148 155428 295204 202748
rect 295260 170578 295316 238252
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 298284 238084 298340 238094
rect 298284 237860 298340 238028
rect 298284 237794 298340 237804
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 295260 170512 295316 170522
rect 295372 236964 295428 236974
rect 295148 155362 295204 155372
rect 295372 141092 295428 236908
rect 298956 236964 299012 236974
rect 298956 199018 299012 236908
rect 305676 236964 305732 236974
rect 298956 198952 299012 198962
rect 301196 200004 301252 200014
rect 301196 198660 301252 199948
rect 301420 200004 301476 200014
rect 301420 199108 301476 199948
rect 301420 199042 301476 199052
rect 301196 198594 301252 198604
rect 305676 197876 305732 236908
rect 308252 236516 308308 236526
rect 308252 202580 308308 236460
rect 308252 202514 308308 202524
rect 308476 234388 308532 234398
rect 308476 202468 308532 234332
rect 308476 202402 308532 202412
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 312618 202350 313238 219922
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 308588 199444 308644 199454
rect 308588 198884 308644 199388
rect 310828 199444 310884 199454
rect 310268 199332 310324 199342
rect 310268 199198 310324 199276
rect 310268 199142 310660 199198
rect 310604 199108 310660 199142
rect 310604 199042 310660 199052
rect 310828 198996 310884 199388
rect 310828 198930 310884 198940
rect 311836 199444 311892 199454
rect 308588 198818 308644 198828
rect 311836 198884 311892 199388
rect 311836 198818 311892 198828
rect 305676 197810 305732 197820
rect 312618 197430 313238 201922
rect 316338 226350 316958 239082
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 316338 208350 316958 225922
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 316338 197430 316958 207922
rect 321692 197398 321748 239282
rect 321804 197764 321860 239820
rect 324268 238308 324324 238318
rect 323372 236278 323428 236288
rect 323372 219268 323428 236222
rect 323372 219202 323428 219212
rect 323932 219604 323988 219614
rect 321804 197698 321860 197708
rect 323148 217588 323204 217598
rect 321692 197332 321748 197342
rect 323148 191458 323204 217532
rect 323372 214452 323428 214462
rect 323148 191392 323204 191402
rect 323260 198996 323316 199006
rect 295508 190350 295828 190384
rect 295508 190294 295578 190350
rect 295634 190294 295702 190350
rect 295758 190294 295828 190350
rect 295508 190226 295828 190294
rect 295508 190170 295578 190226
rect 295634 190170 295702 190226
rect 295758 190170 295828 190226
rect 295508 190102 295828 190170
rect 295508 190046 295578 190102
rect 295634 190046 295702 190102
rect 295758 190046 295828 190102
rect 295508 189978 295828 190046
rect 295508 189922 295578 189978
rect 295634 189922 295702 189978
rect 295758 189922 295828 189978
rect 295508 189888 295828 189922
rect 304832 190350 305152 190384
rect 304832 190294 304902 190350
rect 304958 190294 305026 190350
rect 305082 190294 305152 190350
rect 304832 190226 305152 190294
rect 304832 190170 304902 190226
rect 304958 190170 305026 190226
rect 305082 190170 305152 190226
rect 304832 190102 305152 190170
rect 304832 190046 304902 190102
rect 304958 190046 305026 190102
rect 305082 190046 305152 190102
rect 304832 189978 305152 190046
rect 304832 189922 304902 189978
rect 304958 189922 305026 189978
rect 305082 189922 305152 189978
rect 304832 189888 305152 189922
rect 314156 190350 314476 190384
rect 314156 190294 314226 190350
rect 314282 190294 314350 190350
rect 314406 190294 314476 190350
rect 314156 190226 314476 190294
rect 314156 190170 314226 190226
rect 314282 190170 314350 190226
rect 314406 190170 314476 190226
rect 314156 190102 314476 190170
rect 314156 190046 314226 190102
rect 314282 190046 314350 190102
rect 314406 190046 314476 190102
rect 314156 189978 314476 190046
rect 314156 189922 314226 189978
rect 314282 189922 314350 189978
rect 314406 189922 314476 189978
rect 314156 189888 314476 189922
rect 300170 184350 300490 184384
rect 300170 184294 300240 184350
rect 300296 184294 300364 184350
rect 300420 184294 300490 184350
rect 300170 184226 300490 184294
rect 300170 184170 300240 184226
rect 300296 184170 300364 184226
rect 300420 184170 300490 184226
rect 300170 184102 300490 184170
rect 300170 184046 300240 184102
rect 300296 184046 300364 184102
rect 300420 184046 300490 184102
rect 300170 183978 300490 184046
rect 300170 183922 300240 183978
rect 300296 183922 300364 183978
rect 300420 183922 300490 183978
rect 300170 183888 300490 183922
rect 309494 184350 309814 184384
rect 309494 184294 309564 184350
rect 309620 184294 309688 184350
rect 309744 184294 309814 184350
rect 309494 184226 309814 184294
rect 309494 184170 309564 184226
rect 309620 184170 309688 184226
rect 309744 184170 309814 184226
rect 309494 184102 309814 184170
rect 309494 184046 309564 184102
rect 309620 184046 309688 184102
rect 309744 184046 309814 184102
rect 309494 183978 309814 184046
rect 309494 183922 309564 183978
rect 309620 183922 309688 183978
rect 309744 183922 309814 183978
rect 309494 183888 309814 183922
rect 318818 184350 319138 184384
rect 318818 184294 318888 184350
rect 318944 184294 319012 184350
rect 319068 184294 319138 184350
rect 318818 184226 319138 184294
rect 318818 184170 318888 184226
rect 318944 184170 319012 184226
rect 319068 184170 319138 184226
rect 318818 184102 319138 184170
rect 318818 184046 318888 184102
rect 318944 184046 319012 184102
rect 319068 184046 319138 184102
rect 318818 183978 319138 184046
rect 318818 183922 318888 183978
rect 318944 183922 319012 183978
rect 319068 183922 319138 183978
rect 318818 183888 319138 183922
rect 295508 172350 295828 172384
rect 295508 172294 295578 172350
rect 295634 172294 295702 172350
rect 295758 172294 295828 172350
rect 295508 172226 295828 172294
rect 295508 172170 295578 172226
rect 295634 172170 295702 172226
rect 295758 172170 295828 172226
rect 295508 172102 295828 172170
rect 295508 172046 295578 172102
rect 295634 172046 295702 172102
rect 295758 172046 295828 172102
rect 295508 171978 295828 172046
rect 295508 171922 295578 171978
rect 295634 171922 295702 171978
rect 295758 171922 295828 171978
rect 295508 171888 295828 171922
rect 304832 172350 305152 172384
rect 304832 172294 304902 172350
rect 304958 172294 305026 172350
rect 305082 172294 305152 172350
rect 304832 172226 305152 172294
rect 304832 172170 304902 172226
rect 304958 172170 305026 172226
rect 305082 172170 305152 172226
rect 304832 172102 305152 172170
rect 304832 172046 304902 172102
rect 304958 172046 305026 172102
rect 305082 172046 305152 172102
rect 304832 171978 305152 172046
rect 304832 171922 304902 171978
rect 304958 171922 305026 171978
rect 305082 171922 305152 171978
rect 304832 171888 305152 171922
rect 314156 172350 314476 172384
rect 314156 172294 314226 172350
rect 314282 172294 314350 172350
rect 314406 172294 314476 172350
rect 314156 172226 314476 172294
rect 314156 172170 314226 172226
rect 314282 172170 314350 172226
rect 314406 172170 314476 172226
rect 314156 172102 314476 172170
rect 314156 172046 314226 172102
rect 314282 172046 314350 172102
rect 314406 172046 314476 172102
rect 314156 171978 314476 172046
rect 314156 171922 314226 171978
rect 314282 171922 314350 171978
rect 314406 171922 314476 171978
rect 314156 171888 314476 171922
rect 297500 170578 297556 170588
rect 295372 141026 295428 141036
rect 297388 169858 297444 169868
rect 297388 135658 297444 169802
rect 297500 160356 297556 170522
rect 300170 166350 300490 166384
rect 300170 166294 300240 166350
rect 300296 166294 300364 166350
rect 300420 166294 300490 166350
rect 300170 166226 300490 166294
rect 300170 166170 300240 166226
rect 300296 166170 300364 166226
rect 300420 166170 300490 166226
rect 300170 166102 300490 166170
rect 300170 166046 300240 166102
rect 300296 166046 300364 166102
rect 300420 166046 300490 166102
rect 300170 165978 300490 166046
rect 300170 165922 300240 165978
rect 300296 165922 300364 165978
rect 300420 165922 300490 165978
rect 300170 165888 300490 165922
rect 309494 166350 309814 166384
rect 309494 166294 309564 166350
rect 309620 166294 309688 166350
rect 309744 166294 309814 166350
rect 309494 166226 309814 166294
rect 309494 166170 309564 166226
rect 309620 166170 309688 166226
rect 309744 166170 309814 166226
rect 309494 166102 309814 166170
rect 309494 166046 309564 166102
rect 309620 166046 309688 166102
rect 309744 166046 309814 166102
rect 309494 165978 309814 166046
rect 309494 165922 309564 165978
rect 309620 165922 309688 165978
rect 309744 165922 309814 165978
rect 309494 165888 309814 165922
rect 312618 166350 313238 170618
rect 312618 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 313238 166350
rect 312618 166226 313238 166294
rect 312618 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 313238 166226
rect 312618 166102 313238 166170
rect 312618 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 313238 166102
rect 312618 165978 313238 166046
rect 312618 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 313238 165978
rect 297500 160290 297556 160300
rect 312618 148350 313238 165922
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 297388 134578 297444 135602
rect 297388 134512 297444 134522
rect 306572 136918 306628 136928
rect 304892 132778 304948 132788
rect 304892 116788 304948 132722
rect 304892 116722 304948 116732
rect 306572 113876 306628 136862
rect 306572 113810 306628 113820
rect 312618 130350 313238 147922
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 295036 98354 295092 98364
rect 312618 112350 313238 129922
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 294812 98242 294868 98252
rect 312618 94350 313238 111922
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 299500 82147 299820 82204
rect 299500 82091 299528 82147
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 299820 82147
rect 299500 82043 299820 82091
rect 299500 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 299820 82043
rect 299500 81939 299820 81987
rect 299500 81883 299528 81939
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 299820 81939
rect 299500 81826 299820 81883
rect 307816 82147 308136 82204
rect 307816 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 308136 82147
rect 307816 82043 308136 82091
rect 307816 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 308136 82043
rect 307816 81939 308136 81987
rect 307816 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 308136 81939
rect 307816 81826 308136 81883
rect 312618 77350 313238 93922
rect 316338 154350 316958 170618
rect 318818 166350 319138 166384
rect 318818 166294 318888 166350
rect 318944 166294 319012 166350
rect 319068 166294 319138 166350
rect 318818 166226 319138 166294
rect 318818 166170 318888 166226
rect 318944 166170 319012 166226
rect 319068 166170 319138 166226
rect 318818 166102 319138 166170
rect 318818 166046 318888 166102
rect 318944 166046 319012 166102
rect 319068 166046 319138 166102
rect 318818 165978 319138 166046
rect 318818 165922 318888 165978
rect 318944 165922 319012 165978
rect 319068 165922 319138 165978
rect 318818 165888 319138 165922
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 316338 136350 316958 153922
rect 323260 140532 323316 198940
rect 323372 197764 323428 214396
rect 323372 197698 323428 197708
rect 323480 190350 323800 190384
rect 323480 190294 323550 190350
rect 323606 190294 323674 190350
rect 323730 190294 323800 190350
rect 323480 190226 323800 190294
rect 323480 190170 323550 190226
rect 323606 190170 323674 190226
rect 323730 190170 323800 190226
rect 323480 190102 323800 190170
rect 323480 190046 323550 190102
rect 323606 190046 323674 190102
rect 323730 190046 323800 190102
rect 323480 189978 323800 190046
rect 323480 189922 323550 189978
rect 323606 189922 323674 189978
rect 323730 189922 323800 189978
rect 323480 189888 323800 189922
rect 323480 172350 323800 172384
rect 323480 172294 323550 172350
rect 323606 172294 323674 172350
rect 323730 172294 323800 172350
rect 323480 172226 323800 172294
rect 323480 172170 323550 172226
rect 323606 172170 323674 172226
rect 323730 172170 323800 172226
rect 323480 172102 323800 172170
rect 323480 172046 323550 172102
rect 323606 172046 323674 172102
rect 323730 172046 323800 172102
rect 323480 171978 323800 172046
rect 323480 171922 323550 171978
rect 323606 171922 323674 171978
rect 323730 171922 323800 171978
rect 323480 171888 323800 171922
rect 323260 140466 323316 140476
rect 323932 138628 323988 219548
rect 324044 199108 324100 199118
rect 324044 140756 324100 199052
rect 324268 158788 324324 238252
rect 325836 238308 325892 238318
rect 325724 238196 325780 238206
rect 324268 158722 324324 158732
rect 325052 236852 325108 236862
rect 324044 140690 324100 140700
rect 323932 138562 323988 138572
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 84316 316958 99922
rect 316132 82147 316452 82204
rect 316132 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 316452 82147
rect 316132 82043 316452 82091
rect 316132 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 316452 82043
rect 316132 81939 316452 81987
rect 316132 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 316452 81939
rect 316132 81826 316452 81883
rect 324448 82147 324768 82204
rect 324448 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82091 324768 82147
rect 324448 82043 324768 82091
rect 324448 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 324768 82043
rect 324448 81939 324768 81987
rect 324448 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81883 324768 81939
rect 324448 81826 324768 81883
rect 295342 76350 295662 76384
rect 295342 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 295662 76350
rect 295342 76226 295662 76294
rect 295342 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 295662 76226
rect 295342 76102 295662 76170
rect 295342 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 295662 76102
rect 295342 75978 295662 76046
rect 295342 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 295662 75978
rect 295342 75888 295662 75922
rect 303658 76350 303978 76384
rect 303658 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 303978 76350
rect 303658 76226 303978 76294
rect 303658 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 303978 76226
rect 303658 76102 303978 76170
rect 303658 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 303978 76102
rect 303658 75978 303978 76046
rect 303658 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 303978 75978
rect 303658 75888 303978 75922
rect 311974 76350 312294 76384
rect 311974 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 312294 76350
rect 311974 76226 312294 76294
rect 311974 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 312294 76226
rect 311974 76102 312294 76170
rect 311974 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 312294 76102
rect 311974 75978 312294 76046
rect 311974 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 312294 75978
rect 311974 75888 312294 75922
rect 320290 76350 320610 76384
rect 320290 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 320610 76350
rect 320290 76226 320610 76294
rect 320290 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 320610 76226
rect 320290 76102 320610 76170
rect 320290 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 320610 76102
rect 320290 75978 320610 76046
rect 320290 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 320610 75978
rect 320290 75888 320610 75922
rect 299500 64350 299820 64384
rect 299500 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 299820 64350
rect 299500 64226 299820 64294
rect 299500 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 299820 64226
rect 299500 64102 299820 64170
rect 299500 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 299820 64102
rect 299500 63978 299820 64046
rect 299500 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 299820 63978
rect 299500 63888 299820 63922
rect 307816 64350 308136 64384
rect 307816 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 308136 64350
rect 307816 64226 308136 64294
rect 307816 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 308136 64226
rect 307816 64102 308136 64170
rect 307816 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 308136 64102
rect 307816 63978 308136 64046
rect 307816 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 308136 63978
rect 307816 63888 308136 63922
rect 316132 64350 316452 64384
rect 316132 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 316452 64350
rect 316132 64226 316452 64294
rect 316132 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 316452 64226
rect 316132 64102 316452 64170
rect 316132 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 316452 64102
rect 316132 63978 316452 64046
rect 316132 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 316452 63978
rect 316132 63888 316452 63922
rect 324448 64350 324768 64384
rect 324448 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 324768 64350
rect 324448 64226 324768 64294
rect 324448 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 324768 64226
rect 324448 64102 324768 64170
rect 324448 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 324768 64102
rect 324448 63978 324768 64046
rect 324448 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 324768 63978
rect 324448 63888 324768 63922
rect 295342 58350 295662 58384
rect 295342 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 295662 58350
rect 295342 58226 295662 58294
rect 295342 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 295662 58226
rect 295342 58102 295662 58170
rect 295342 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 295662 58102
rect 295342 57978 295662 58046
rect 295342 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 295662 57978
rect 295342 57888 295662 57922
rect 303658 58350 303978 58384
rect 303658 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 303978 58350
rect 303658 58226 303978 58294
rect 303658 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 303978 58226
rect 303658 58102 303978 58170
rect 303658 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 303978 58102
rect 303658 57978 303978 58046
rect 303658 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 303978 57978
rect 303658 57888 303978 57922
rect 311974 58350 312294 58384
rect 311974 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 312294 58350
rect 311974 58226 312294 58294
rect 311974 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 312294 58226
rect 311974 58102 312294 58170
rect 311974 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 312294 58102
rect 311974 57978 312294 58046
rect 311974 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 312294 57978
rect 311974 57888 312294 57922
rect 320290 58350 320610 58384
rect 320290 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 320610 58350
rect 320290 58226 320610 58294
rect 320290 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 320610 58226
rect 320290 58102 320610 58170
rect 320290 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 320610 58102
rect 320290 57978 320610 58046
rect 320290 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 320610 57978
rect 320290 57888 320610 57922
rect 291564 47618 291620 47628
rect 291452 44482 291508 44492
rect 289772 41122 289828 41132
rect 288204 37762 288260 37772
rect 312618 40350 313238 53674
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 288092 29362 288148 29372
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 285618 -1120 286238 9922
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 22350 313238 39922
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 312618 4350 313238 21922
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 46350 316958 50964
rect 325052 50708 325108 236796
rect 325276 232932 325332 232942
rect 325164 229460 325220 229470
rect 325164 157798 325220 229404
rect 325276 210898 325332 232876
rect 325276 210832 325332 210842
rect 325388 202692 325444 202702
rect 325164 157732 325220 157742
rect 325276 199444 325332 199454
rect 325276 138740 325332 199388
rect 325388 153860 325444 202636
rect 325388 153794 325444 153804
rect 325276 138674 325332 138684
rect 325724 105252 325780 238140
rect 325724 105186 325780 105196
rect 325836 98644 325892 238252
rect 326508 235956 326564 240604
rect 326508 235890 326564 235900
rect 326620 230916 326676 240722
rect 326620 230850 326676 230860
rect 326732 227668 326788 240902
rect 326844 240598 326900 240608
rect 326844 235172 326900 240542
rect 326844 235106 326900 235116
rect 326956 240418 327012 240428
rect 326732 227602 326788 227612
rect 326732 221060 326788 221070
rect 326620 198660 326676 198670
rect 326620 162118 326676 198604
rect 326620 162052 326676 162062
rect 326732 98756 326788 221004
rect 326956 200004 327012 240362
rect 326956 199938 327012 199948
rect 327068 238618 327124 238628
rect 326844 199018 326900 199028
rect 326844 140338 326900 198962
rect 327068 188132 327124 238562
rect 327404 237718 327460 248102
rect 327068 188066 327124 188076
rect 327180 237662 327460 237718
rect 327516 240436 327572 240446
rect 327180 155458 327236 237662
rect 327516 237538 327572 240380
rect 327180 155392 327236 155402
rect 327292 237482 327572 237538
rect 327628 239338 327684 239348
rect 326844 140272 326900 140282
rect 327292 108612 327348 237482
rect 327628 237358 327684 239282
rect 327516 237302 327684 237358
rect 327292 108546 327348 108556
rect 327404 235956 327460 235966
rect 326732 98690 326788 98700
rect 325836 98578 325892 98588
rect 327404 51492 327460 235900
rect 327404 51426 327460 51436
rect 325052 50642 325108 50652
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 316338 10350 316958 27922
rect 327516 20132 327572 237302
rect 327628 210868 327684 210878
rect 327628 166068 327684 210812
rect 327628 166002 327684 166012
rect 327628 161924 327684 161934
rect 327628 146132 327684 161868
rect 327628 146066 327684 146076
rect 327964 134148 328020 260342
rect 328076 155876 328132 311642
rect 328412 282718 328468 379682
rect 328524 313318 328580 407596
rect 335132 407458 335188 407468
rect 333564 399028 333620 399038
rect 332780 397378 332836 397388
rect 330316 390292 330372 390302
rect 330204 389956 330260 389966
rect 329756 388836 329812 388846
rect 328636 380548 328692 380558
rect 328636 379652 328692 380492
rect 328636 379586 328692 379596
rect 329084 379652 329140 379662
rect 329084 369658 329140 379596
rect 329084 369592 329140 369602
rect 329420 372260 329476 372270
rect 329308 326564 329364 326574
rect 329308 326458 329364 326508
rect 328748 326402 329364 326458
rect 328524 313252 328580 313262
rect 328636 321058 328692 321068
rect 328412 282652 328468 282662
rect 328524 313138 328580 313148
rect 328412 258598 328468 258608
rect 328300 249238 328356 249248
rect 328300 231812 328356 249182
rect 328412 233268 328468 258542
rect 328524 240324 328580 313082
rect 328636 249598 328692 321002
rect 328748 283798 328804 326402
rect 329308 323876 329364 323886
rect 329308 323758 329364 323820
rect 328860 323702 329364 323758
rect 328860 308278 328916 323702
rect 329308 321188 329364 321198
rect 329308 321058 329364 321132
rect 329308 320992 329364 321002
rect 328860 308212 328916 308222
rect 328972 314020 329364 314038
rect 328972 313982 329308 314020
rect 328748 283732 328804 283742
rect 328860 296578 328916 296588
rect 328636 249532 328692 249542
rect 328748 283078 328804 283088
rect 328748 249418 328804 283022
rect 328748 249352 328804 249362
rect 328524 240258 328580 240268
rect 328636 248338 328692 248348
rect 328636 236852 328692 248282
rect 328636 236786 328692 236796
rect 328748 242218 328804 242228
rect 328748 233380 328804 242162
rect 328748 233314 328804 233324
rect 328412 233202 328468 233212
rect 328300 231746 328356 231756
rect 328636 204484 328692 204494
rect 328076 155810 328132 155820
rect 328412 202580 328468 202590
rect 327964 134082 328020 134092
rect 328412 110180 328468 202524
rect 328524 200004 328580 200014
rect 328524 150836 328580 199948
rect 328636 174692 328692 204428
rect 328636 174626 328692 174636
rect 328860 156212 328916 296522
rect 328972 158698 329028 313982
rect 329308 313954 329364 313964
rect 329308 313138 329364 313162
rect 329308 313058 329364 313068
rect 329084 300898 329140 300908
rect 329084 285778 329140 300842
rect 329084 285712 329140 285722
rect 329308 282718 329364 282728
rect 329308 282660 329364 282662
rect 329308 282594 329364 282604
rect 329084 272998 329140 273008
rect 329084 265618 329140 272942
rect 329308 265636 329364 265646
rect 329084 265580 329308 265618
rect 329084 265562 329364 265580
rect 329420 260398 329476 372204
rect 329420 260332 329476 260342
rect 329532 333732 329588 333742
rect 329196 253738 329252 253748
rect 329084 248518 329140 248528
rect 329084 242038 329140 248462
rect 329196 247978 329252 253682
rect 329196 247912 329252 247922
rect 329084 241972 329140 241982
rect 329532 240418 329588 333676
rect 329756 331940 329812 388780
rect 329756 331874 329812 331884
rect 330092 378756 330148 378766
rect 329756 329252 329812 329262
rect 329084 240362 329588 240418
rect 329644 296996 329700 297006
rect 329084 189028 329140 240362
rect 329084 188962 329140 188972
rect 328972 158632 329028 158642
rect 328860 156146 328916 156156
rect 328524 150770 328580 150780
rect 328412 110114 328468 110124
rect 329644 101892 329700 296940
rect 329756 253738 329812 329196
rect 329980 308278 330036 308288
rect 329868 297892 329924 297902
rect 329868 264292 329924 297836
rect 329868 264226 329924 264236
rect 329980 258692 330036 308222
rect 330092 279636 330148 378700
rect 330204 308868 330260 389900
rect 330204 308802 330260 308812
rect 330092 279570 330148 279580
rect 330204 285778 330260 285788
rect 330204 265524 330260 285722
rect 330316 285348 330372 390236
rect 331548 388052 331604 388062
rect 331548 386578 331604 387996
rect 331548 386512 331604 386522
rect 331772 383698 331828 383708
rect 330428 373156 330484 373166
rect 330428 296578 330484 373100
rect 330988 356132 331044 356142
rect 330428 296512 330484 296522
rect 330876 299348 330932 299358
rect 330316 285282 330372 285292
rect 330540 285796 330596 285806
rect 330540 272998 330596 285740
rect 330876 285684 330932 299292
rect 330876 285618 330932 285628
rect 330540 272932 330596 272942
rect 330652 275604 330708 275614
rect 330204 265458 330260 265468
rect 330540 264068 330596 264078
rect 330316 260372 330372 260382
rect 329980 258626 330036 258636
rect 330092 259924 330148 259934
rect 330092 255388 330148 259868
rect 329756 253672 329812 253682
rect 329868 255332 330148 255388
rect 329756 245364 329812 245374
rect 329756 236278 329812 245308
rect 329756 236212 329812 236222
rect 329644 101826 329700 101836
rect 329868 98532 329924 255332
rect 330092 252532 330148 252542
rect 329980 252420 330036 252430
rect 329980 240436 330036 252364
rect 329980 240370 330036 240380
rect 330092 235060 330148 252476
rect 330092 234994 330148 235004
rect 330204 240324 330260 240334
rect 330092 225988 330148 225998
rect 330092 98868 330148 225932
rect 330204 140980 330260 240268
rect 330316 238308 330372 260316
rect 330316 238242 330372 238252
rect 330428 249598 330484 249608
rect 330204 140914 330260 140924
rect 330316 236180 330372 236190
rect 330316 99988 330372 236124
rect 330428 136052 330484 249542
rect 330540 245028 330596 264012
rect 330540 244962 330596 244972
rect 330428 135986 330484 135996
rect 330540 236292 330596 236302
rect 330540 100100 330596 236236
rect 330652 132132 330708 275548
rect 330764 272692 330820 272702
rect 330764 250404 330820 272636
rect 330764 250338 330820 250348
rect 330876 258580 330932 258590
rect 330876 248158 330932 258524
rect 330988 248518 331044 356076
rect 330988 248452 331044 248462
rect 331100 331044 331156 331054
rect 330876 248092 330932 248102
rect 330988 247044 331044 247054
rect 330876 244916 330932 244926
rect 330876 238196 330932 244860
rect 330988 242116 331044 246988
rect 330988 242050 331044 242060
rect 331100 240418 331156 330988
rect 331772 301618 331828 383642
rect 332668 376498 332724 376508
rect 332668 343588 332724 376442
rect 332668 343522 332724 343532
rect 332108 334628 332164 334638
rect 331772 301552 331828 301562
rect 331996 320292 332052 320302
rect 331884 301476 331940 301486
rect 331772 300580 331828 300590
rect 331324 299684 331380 299694
rect 331212 298788 331268 298798
rect 331212 252420 331268 298732
rect 331324 264068 331380 299628
rect 331324 264002 331380 264012
rect 331660 264628 331716 264638
rect 331660 258580 331716 264572
rect 331660 258514 331716 258524
rect 331212 252354 331268 252364
rect 331212 248724 331268 248734
rect 331212 248338 331268 248668
rect 331212 248272 331268 248282
rect 331100 240352 331156 240362
rect 331660 242038 331716 242048
rect 331548 238644 331604 238654
rect 331548 238550 331604 238562
rect 330876 238130 330932 238140
rect 330652 132066 330708 132076
rect 330764 189812 330820 189822
rect 330540 100034 330596 100044
rect 330316 99922 330372 99932
rect 330092 98802 330148 98812
rect 329868 98466 329924 98476
rect 330764 31798 330820 189756
rect 331660 151172 331716 241982
rect 331660 151106 331716 151116
rect 331772 115332 331828 300524
rect 331884 118692 331940 301420
rect 331996 142678 332052 320236
rect 332108 287476 332164 334572
rect 332332 322084 332388 322094
rect 332220 308868 332276 308878
rect 332220 299124 332276 308812
rect 332220 299058 332276 299068
rect 332108 287410 332164 287420
rect 332108 282212 332164 282222
rect 332108 275604 332164 282156
rect 332108 275538 332164 275548
rect 332108 268772 332164 268782
rect 332108 245252 332164 268716
rect 332332 268100 332388 322028
rect 332556 316036 332612 316046
rect 332444 305732 332500 305742
rect 332444 297444 332500 305676
rect 332556 299236 332612 315980
rect 332556 299170 332612 299180
rect 332444 297378 332500 297388
rect 332668 299124 332724 299134
rect 332668 287140 332724 299068
rect 332780 296324 332836 397322
rect 333116 394884 333172 394894
rect 333004 389998 333060 390008
rect 332780 296258 332836 296268
rect 332892 389818 332948 389828
rect 332780 296100 332836 296110
rect 332780 293412 332836 296044
rect 332780 293346 332836 293356
rect 332668 287074 332724 287084
rect 332780 293188 332836 293198
rect 332668 281428 332724 281438
rect 332668 276388 332724 281372
rect 332668 276322 332724 276332
rect 332332 268034 332388 268044
rect 332556 273924 332612 273934
rect 332108 245186 332164 245196
rect 332220 253764 332276 253774
rect 331996 142612 332052 142622
rect 332108 245028 332164 245038
rect 331884 118626 331940 118636
rect 331772 115266 331828 115276
rect 332108 111972 332164 244972
rect 332220 240660 332276 253708
rect 332444 250404 332500 250414
rect 332332 249508 332388 249518
rect 332332 240778 332388 249452
rect 332444 246932 332500 250348
rect 332444 246866 332500 246876
rect 332332 240712 332388 240722
rect 332444 240772 332500 240782
rect 332220 240594 332276 240604
rect 332332 238644 332388 238654
rect 332108 111906 332164 111916
rect 332220 227638 332276 227648
rect 332220 101668 332276 227582
rect 332332 146998 332388 238588
rect 332332 146932 332388 146942
rect 332444 141958 332500 240716
rect 332444 141892 332500 141902
rect 332556 125412 332612 273868
rect 332668 266532 332724 266542
rect 332668 258598 332724 266476
rect 332668 258532 332724 258542
rect 332668 253204 332724 253214
rect 332668 249238 332724 253148
rect 332780 250404 332836 293132
rect 332892 289828 332948 389762
rect 333004 291620 333060 389942
rect 333116 308084 333172 394828
rect 333452 394212 333508 394222
rect 333228 391618 333284 391628
rect 333228 308308 333284 391562
rect 333340 370468 333396 370478
rect 333340 317044 333396 370412
rect 333452 344484 333508 394156
rect 333452 344418 333508 344428
rect 333340 316978 333396 316988
rect 333228 308242 333284 308252
rect 333116 308018 333172 308028
rect 333004 291554 333060 291564
rect 333116 305060 333172 305070
rect 332892 289762 332948 289772
rect 332892 283798 332948 283808
rect 332892 272692 332948 283742
rect 333116 282212 333172 305004
rect 333228 302372 333284 302382
rect 333228 293748 333284 302316
rect 333228 293682 333284 293692
rect 333340 296324 333396 296334
rect 333340 293188 333396 296268
rect 333340 293122 333396 293132
rect 333116 282146 333172 282156
rect 333564 292516 333620 398972
rect 334460 393316 334516 393326
rect 334348 393204 334404 393214
rect 333788 315812 333844 315822
rect 333676 308644 333732 308654
rect 333676 300916 333732 308588
rect 333788 305732 333844 315756
rect 333788 305666 333844 305676
rect 334012 306852 334068 306862
rect 334012 302148 334068 306796
rect 334348 305758 334404 393148
rect 334460 328356 334516 393260
rect 334572 384778 334628 384788
rect 334572 334404 334628 384722
rect 334572 334338 334628 334348
rect 334460 328290 334516 328300
rect 334572 332836 334628 332846
rect 334012 302082 334068 302092
rect 334124 305702 334404 305758
rect 334460 318500 334516 318510
rect 333676 300850 333732 300860
rect 333116 279972 333172 279982
rect 333116 275940 333172 279916
rect 333564 278908 333620 292460
rect 334124 290668 334180 305702
rect 334348 303268 334404 303278
rect 333900 290612 334180 290668
rect 334236 293972 334292 293982
rect 333900 284452 333956 290612
rect 333900 284386 333956 284396
rect 333116 275874 333172 275884
rect 333228 278852 333620 278908
rect 332892 272626 332948 272636
rect 332780 250338 332836 250348
rect 332892 271908 332948 271918
rect 332668 249172 332724 249182
rect 332668 243460 332724 243470
rect 332668 236740 332724 243404
rect 332892 242004 332948 271852
rect 333004 264292 333060 264302
rect 333004 256228 333060 264236
rect 333228 260372 333284 278852
rect 333452 275716 333508 275726
rect 333228 260306 333284 260316
rect 333340 261156 333396 261166
rect 333004 256162 333060 256172
rect 333116 255780 333172 255790
rect 332892 241938 332948 241948
rect 333004 248948 333060 248958
rect 332668 236674 332724 236684
rect 332668 236068 332724 236078
rect 332668 198212 332724 236012
rect 333004 231058 333060 248892
rect 333116 242218 333172 255724
rect 333228 254884 333284 254894
rect 333228 245476 333284 254828
rect 333228 245410 333284 245420
rect 333116 242152 333172 242162
rect 333340 240598 333396 261100
rect 333452 252084 333508 275660
rect 334124 275604 334180 275614
rect 334124 263732 334180 275548
rect 334236 266308 334292 293916
rect 334348 273924 334404 303212
rect 334460 293860 334516 318444
rect 334460 293794 334516 293804
rect 334348 273858 334404 273868
rect 334460 281764 334516 281774
rect 334236 266242 334292 266252
rect 334124 263666 334180 263676
rect 333788 262948 333844 262958
rect 333452 252018 333508 252028
rect 333676 257124 333732 257134
rect 333340 240532 333396 240542
rect 333452 250628 333508 250638
rect 333452 238588 333508 250572
rect 333228 238532 333508 238588
rect 333564 247978 333620 247988
rect 333228 231700 333284 238532
rect 333228 231634 333284 231644
rect 333004 230992 333060 231002
rect 332668 197540 332724 198156
rect 332668 197474 332724 197484
rect 333452 217558 333508 217568
rect 333340 135298 333396 135308
rect 332556 125346 332612 125356
rect 332668 134372 332724 134382
rect 332220 101602 332276 101612
rect 332668 83188 332724 134316
rect 333340 134372 333396 135242
rect 333340 134306 333396 134316
rect 333452 98980 333508 217502
rect 333564 152180 333620 247922
rect 333676 245364 333732 257068
rect 333788 253652 333844 262892
rect 334236 260372 334292 260382
rect 334236 255332 334292 260316
rect 334236 255266 334292 255276
rect 334348 256228 334404 256238
rect 333788 253586 333844 253596
rect 333676 245298 333732 245308
rect 333788 251300 333844 251310
rect 333676 243460 333732 243470
rect 333676 235844 333732 243404
rect 333676 152964 333732 235788
rect 333788 234500 333844 251244
rect 334348 250348 334404 256172
rect 334236 250292 334404 250348
rect 334124 246932 334180 246942
rect 333788 234434 333844 234444
rect 333900 243572 333956 243582
rect 333900 229258 333956 243516
rect 334124 243236 334180 246876
rect 334236 244916 334292 250292
rect 334236 244850 334292 244860
rect 334124 243170 334180 243180
rect 334236 243796 334292 243806
rect 333900 229192 333956 229202
rect 333788 226100 333844 226110
rect 333788 155638 333844 226044
rect 333900 198212 333956 198222
rect 333900 178500 333956 198156
rect 333900 173068 333956 178444
rect 334124 188132 334180 188142
rect 334124 184996 334180 188076
rect 333900 173012 334068 173068
rect 333788 155572 333844 155582
rect 333676 152898 333732 152908
rect 333564 152114 333620 152124
rect 333900 127558 333956 127568
rect 333900 121828 333956 127502
rect 333900 121762 333956 121772
rect 334012 100212 334068 173012
rect 334124 107044 334180 184940
rect 334124 106978 334180 106988
rect 334012 100146 334068 100156
rect 333452 98914 333508 98924
rect 332668 83122 332724 83132
rect 334236 33598 334292 243740
rect 334460 240100 334516 281708
rect 334572 280868 334628 332780
rect 334684 319396 334740 319406
rect 334684 297220 334740 319340
rect 334796 314916 334852 314926
rect 334796 304052 334852 314860
rect 334796 303986 334852 303996
rect 335020 305956 335076 305966
rect 334684 297154 334740 297164
rect 334572 280802 334628 280812
rect 334684 293412 334740 293422
rect 334572 275940 334628 275950
rect 334572 240212 334628 275884
rect 334684 259924 334740 293356
rect 335020 290388 335076 305900
rect 335020 290322 335076 290332
rect 334684 259858 334740 259868
rect 334796 287476 334852 287486
rect 334796 257124 334852 287420
rect 334796 257058 334852 257068
rect 334908 283556 334964 283566
rect 334908 253764 334964 283500
rect 334908 253698 334964 253708
rect 335020 280644 335076 280654
rect 334572 240146 334628 240156
rect 334684 253652 334740 253662
rect 334460 240034 334516 240044
rect 334460 239428 334516 239438
rect 334460 188132 334516 239372
rect 334684 238532 334740 253596
rect 334684 238466 334740 238476
rect 334796 245364 334852 245374
rect 334796 189812 334852 245308
rect 335020 240100 335076 280588
rect 335132 277396 335188 407402
rect 336028 407278 336084 407288
rect 335916 383572 335972 383582
rect 335916 383452 335972 383462
rect 335356 369658 335412 369668
rect 335132 277330 335188 277340
rect 335244 293748 335300 293758
rect 335132 263844 335188 263854
rect 335132 243478 335188 263788
rect 335132 243412 335188 243422
rect 335020 240034 335076 240044
rect 335132 240212 335188 240222
rect 334796 189746 334852 189756
rect 335132 238868 335188 240156
rect 334460 188066 334516 188076
rect 335020 142660 335076 142670
rect 335020 137638 335076 142604
rect 335020 137572 335076 137582
rect 335132 42868 335188 238812
rect 335244 122052 335300 293692
rect 335356 291060 335412 369602
rect 335580 322980 335636 322990
rect 335356 290994 335412 291004
rect 335468 304164 335524 304174
rect 335356 286804 335412 286814
rect 335356 282212 335412 286748
rect 335356 282146 335412 282156
rect 335468 260372 335524 304108
rect 335580 294756 335636 322924
rect 336028 300898 336084 407222
rect 336140 402164 336196 402174
rect 336140 401604 336196 402108
rect 336140 401538 336196 401548
rect 336924 392868 336980 410462
rect 354620 410518 354676 410528
rect 359996 410518 360052 410528
rect 352828 410158 352884 410168
rect 352828 409780 352884 410102
rect 352828 409714 352884 409724
rect 340844 408898 340900 408908
rect 339612 407278 339668 407288
rect 336924 392802 336980 392812
rect 337484 406738 337540 406748
rect 337484 392868 337540 406682
rect 338604 406084 338660 406094
rect 338492 404758 338548 404768
rect 337596 402164 337652 402174
rect 337596 399364 337652 402108
rect 337596 399298 337652 399308
rect 337708 399718 337764 399728
rect 337708 396340 337764 399662
rect 337708 396274 337764 396284
rect 337484 392802 337540 392812
rect 337820 388388 337876 388398
rect 336028 300832 336084 300842
rect 336140 384958 336196 384968
rect 335580 294690 335636 294700
rect 335692 296548 335748 296558
rect 335580 285572 335636 285582
rect 335580 283978 335636 285516
rect 335580 283912 335636 283922
rect 335692 283078 335748 296492
rect 336140 286244 336196 384902
rect 336252 380098 336308 380108
rect 336252 289156 336308 380042
rect 337708 378118 337764 378128
rect 336364 360838 336420 360848
rect 336364 360388 336420 360782
rect 336364 360322 336420 360332
rect 336812 327684 336868 327694
rect 336476 317604 336532 317614
rect 336252 289090 336308 289100
rect 336364 315812 336420 315822
rect 336364 314916 336420 315756
rect 336140 286178 336196 286188
rect 335692 283012 335748 283022
rect 336140 283892 336196 283902
rect 336028 263956 336084 263966
rect 335468 260306 335524 260316
rect 335916 260484 335972 260494
rect 335692 255332 335748 255342
rect 335244 121986 335300 121996
rect 335356 240100 335412 240110
rect 335356 239316 335412 240044
rect 335356 44548 335412 239260
rect 335580 239988 335636 239998
rect 335468 232708 335524 232718
rect 335468 106708 335524 232652
rect 335468 106642 335524 106652
rect 335580 47908 335636 239932
rect 335692 128772 335748 255276
rect 335916 248836 335972 260428
rect 336028 257236 336084 263900
rect 336028 257170 336084 257180
rect 336140 257124 336196 283836
rect 336140 257058 336196 257068
rect 336252 257572 336308 257582
rect 336252 256978 336308 257516
rect 336140 256922 336308 256978
rect 335916 248770 335972 248780
rect 336028 252196 336084 252206
rect 336028 248698 336084 252140
rect 335804 248642 336084 248698
rect 335804 231028 335860 248642
rect 336028 245252 336084 245262
rect 336028 243572 336084 245196
rect 336028 243506 336084 243516
rect 336140 234612 336196 256922
rect 336252 253988 336308 253998
rect 336252 239518 336308 253932
rect 336364 240324 336420 314860
rect 336476 299348 336532 317548
rect 336476 299282 336532 299292
rect 336588 302148 336644 302158
rect 336476 259364 336532 259374
rect 336476 253540 336532 259308
rect 336476 253474 336532 253484
rect 336476 250292 336532 250302
rect 336476 244132 336532 250236
rect 336588 247044 336644 302092
rect 336700 287812 336756 287822
rect 336700 277284 336756 287756
rect 336700 277218 336756 277228
rect 336588 246978 336644 246988
rect 336476 244066 336532 244076
rect 336364 240258 336420 240268
rect 336252 239452 336308 239462
rect 336140 234546 336196 234556
rect 335804 230962 335860 230972
rect 335692 128706 335748 128716
rect 335804 202468 335860 202478
rect 335804 110404 335860 202412
rect 336140 198100 336196 198110
rect 336140 197428 336196 198044
rect 336028 191492 336084 191502
rect 336028 191392 336084 191402
rect 336028 174692 336084 174702
rect 336028 173098 336084 174636
rect 336028 173032 336084 173042
rect 336140 171220 336196 197372
rect 336028 168308 336084 168318
rect 336028 168058 336084 168252
rect 336028 167992 336084 168002
rect 336140 162298 336196 171164
rect 336140 162232 336196 162242
rect 336028 147924 336084 147934
rect 336028 142548 336084 147868
rect 336028 142482 336084 142492
rect 336140 143938 336196 143948
rect 335916 142324 335972 142334
rect 335916 134038 335972 142268
rect 336140 140084 336196 143882
rect 336140 140018 336196 140028
rect 336812 136918 336868 327628
rect 336924 313318 336980 313328
rect 336924 262948 336980 313262
rect 337596 308420 337652 308430
rect 337036 300804 337092 300814
rect 337036 288036 337092 300748
rect 337036 287970 337092 287980
rect 336924 262882 336980 262892
rect 337484 262948 337540 262958
rect 337372 247044 337428 247054
rect 337260 246932 337316 246942
rect 336812 136852 336868 136862
rect 336924 243236 336980 243246
rect 336812 134372 336868 134382
rect 335916 133972 335972 133982
rect 336028 134218 336084 134228
rect 336028 132778 336084 134162
rect 336812 134218 336868 134316
rect 336812 134152 336868 134162
rect 336028 132712 336084 132722
rect 335804 110338 335860 110348
rect 336812 132238 336868 132248
rect 336812 99092 336868 132182
rect 336924 101780 336980 243180
rect 337148 214004 337204 214014
rect 337148 213444 337204 213948
rect 336924 101714 336980 101724
rect 337036 197398 337092 197408
rect 336812 99026 336868 99036
rect 337036 99092 337092 197342
rect 337148 143938 337204 213388
rect 337260 198324 337316 246876
rect 337260 198258 337316 198268
rect 337372 183764 337428 246988
rect 337372 183698 337428 183708
rect 337372 182308 337428 182318
rect 337260 179732 337316 179742
rect 337260 155652 337316 179676
rect 337372 156100 337428 182252
rect 337372 156034 337428 156044
rect 337260 155586 337316 155596
rect 337484 149604 337540 262892
rect 337148 143872 337204 143882
rect 337260 149492 337540 149548
rect 337260 139188 337316 149492
rect 337596 147924 337652 308364
rect 337708 277844 337764 378062
rect 337820 300804 337876 388332
rect 338492 379652 338548 404702
rect 338604 382452 338660 406028
rect 338828 405972 338884 405982
rect 338716 402958 338772 402968
rect 338716 392338 338772 402902
rect 338828 396004 338884 405916
rect 339500 404218 339556 404228
rect 338828 395938 338884 395948
rect 339052 402598 339108 402608
rect 338716 392272 338772 392282
rect 339052 382564 339108 402542
rect 339500 397572 339556 404162
rect 339612 399700 339668 407222
rect 340172 404938 340228 404948
rect 340172 402276 340228 404882
rect 340172 402210 340228 402220
rect 339612 399634 339668 399644
rect 339500 397506 339556 397516
rect 340844 396508 340900 408842
rect 354508 408660 354564 408670
rect 354508 408178 354564 408604
rect 354508 408112 354564 408122
rect 342636 407764 342692 407774
rect 340956 406196 341012 406206
rect 340956 403318 341012 406140
rect 342524 404852 342580 404862
rect 342524 404068 342580 404796
rect 342524 404002 342580 404012
rect 340956 403252 341012 403262
rect 341516 403498 341572 403508
rect 341180 402836 341236 402846
rect 341180 399718 341236 402780
rect 341516 400618 341572 403442
rect 342636 402724 342692 407708
rect 350476 407540 350532 407550
rect 347900 405412 347956 405422
rect 347788 405300 347844 405310
rect 342748 404852 342804 404862
rect 342748 402948 342804 404796
rect 342748 402882 342804 402892
rect 346108 404398 346164 404408
rect 342636 402658 342692 402668
rect 346108 401158 346164 404342
rect 346892 403956 346948 403966
rect 346892 403732 346948 403900
rect 346892 403666 346948 403676
rect 347788 403060 347844 405244
rect 347900 403498 347956 405356
rect 350476 404758 350532 407484
rect 352156 406756 352212 406766
rect 352156 406662 352212 406682
rect 354620 406420 354676 410462
rect 359884 410452 359940 410462
rect 359772 410158 359828 410168
rect 359548 410116 359604 410126
rect 354620 406354 354676 406364
rect 354732 409978 354788 409988
rect 354732 405412 354788 409922
rect 359548 409618 359604 410060
rect 359660 409978 359716 409988
rect 359660 409780 359716 409922
rect 359660 409714 359716 409724
rect 359548 409552 359604 409562
rect 356188 408898 356244 408908
rect 356188 408548 356244 408842
rect 356188 408482 356244 408492
rect 356636 408538 356692 408548
rect 354732 405346 354788 405356
rect 354508 405188 354564 405198
rect 350588 405062 351092 405118
rect 350588 404964 350644 405062
rect 350588 404898 350644 404908
rect 350924 404964 350980 404974
rect 350700 404852 350756 404862
rect 350476 404702 350644 404758
rect 347900 403432 347956 403442
rect 347788 402994 347844 403004
rect 350476 403396 350532 403406
rect 350476 402958 350532 403340
rect 350476 402892 350532 402902
rect 350588 402500 350644 404702
rect 350700 402958 350756 404796
rect 350700 402892 350756 402902
rect 350812 404404 350868 404414
rect 350812 402778 350868 404348
rect 350924 403138 350980 404908
rect 351036 403172 351092 405062
rect 354508 404398 354564 405132
rect 354508 404332 354564 404342
rect 356188 405076 356244 405086
rect 351036 403106 351092 403116
rect 351484 404292 351540 404302
rect 350924 403072 350980 403082
rect 350812 402712 350868 402722
rect 351484 402612 351540 404236
rect 356188 403620 356244 405020
rect 356188 403554 356244 403564
rect 351484 402546 351540 402556
rect 352716 403508 352772 403518
rect 350588 402434 350644 402444
rect 352716 401518 352772 403452
rect 356636 403060 356692 408482
rect 358540 407652 358596 407662
rect 357308 405412 357364 405422
rect 357308 404938 357364 405356
rect 357308 404872 357364 404882
rect 357868 404292 357924 404302
rect 357868 403172 357924 404236
rect 357868 403106 357924 403116
rect 356636 402994 356692 403004
rect 352716 401452 352772 401462
rect 358540 401518 358596 407596
rect 359772 403508 359828 410102
rect 359772 403442 359828 403452
rect 359884 402948 359940 410396
rect 359996 403396 360052 410462
rect 365932 410518 365988 410528
rect 362796 407764 362852 407774
rect 362796 407540 362852 407708
rect 362796 407474 362852 407484
rect 362796 406532 362852 406542
rect 362796 406378 362852 406476
rect 362796 406322 362964 406378
rect 362908 404852 362964 406322
rect 362908 404786 362964 404796
rect 364812 404852 364868 404862
rect 359996 403330 360052 403340
rect 363020 404404 363076 404414
rect 359884 402882 359940 402892
rect 361228 403172 361284 403182
rect 358540 401452 358596 401462
rect 361228 401518 361284 403116
rect 363020 403060 363076 404348
rect 364700 404404 364756 404414
rect 364700 403732 364756 404348
rect 364700 403666 364756 403676
rect 364812 403138 364868 404796
rect 365932 403858 365988 410462
rect 366268 410158 366324 410168
rect 366268 409780 366324 410102
rect 371308 410158 371364 410168
rect 366268 409714 366324 409724
rect 369628 409978 369684 409988
rect 366044 408996 366100 409006
rect 366044 404758 366100 408940
rect 369628 408996 369684 409922
rect 369628 408930 369684 408940
rect 366156 408718 366212 408728
rect 366156 408212 366212 408662
rect 366156 408146 366212 408156
rect 371308 405636 371364 410102
rect 386204 410158 386260 410168
rect 386092 409978 386148 409988
rect 386092 409108 386148 409922
rect 386204 409892 386260 410102
rect 386204 409826 386260 409836
rect 404908 410158 404964 410168
rect 404908 409892 404964 410102
rect 404908 409826 404964 409836
rect 478828 409332 478884 575148
rect 480620 575092 480676 575102
rect 478940 573860 478996 573870
rect 478940 410116 478996 573804
rect 480508 573748 480564 573758
rect 478940 410050 478996 410060
rect 479052 572180 479108 572190
rect 478828 409266 478884 409276
rect 479052 409220 479108 572124
rect 479164 570388 479220 570398
rect 479164 410228 479220 570332
rect 479164 410162 479220 410172
rect 479276 567364 479332 567374
rect 479052 409154 479108 409164
rect 386092 409042 386148 409052
rect 374668 408660 374724 408670
rect 371308 405570 371364 405580
rect 372764 406644 372820 406654
rect 367948 405188 368004 405198
rect 366044 404692 366100 404702
rect 367612 404964 367668 404974
rect 366156 404404 366212 404414
rect 366156 404038 366212 404348
rect 366156 403972 366212 403982
rect 365932 403792 365988 403802
rect 367612 403844 367668 404908
rect 367836 404964 367892 404974
rect 367836 404292 367892 404908
rect 367836 404226 367892 404236
rect 367612 403778 367668 403788
rect 364812 403072 364868 403082
rect 363020 402994 363076 403004
rect 366156 402958 366212 402968
rect 366156 402612 366212 402902
rect 367948 402778 368004 405132
rect 366156 402546 366212 402556
rect 367836 402724 367892 402734
rect 367948 402712 368004 402722
rect 361228 401452 361284 401462
rect 367836 401518 367892 402668
rect 372764 402388 372820 406588
rect 373660 404292 373716 404302
rect 373660 402948 373716 404236
rect 374556 404068 374612 404078
rect 374556 403508 374612 404012
rect 374556 403442 374612 403452
rect 374668 403060 374724 408604
rect 384860 408548 384916 408558
rect 383068 406756 383124 406766
rect 383068 405658 383124 406700
rect 383068 405592 383124 405602
rect 383180 404516 383236 404526
rect 374668 402994 374724 403004
rect 383068 403318 383124 403328
rect 383068 403060 383124 403262
rect 383068 402994 383124 403004
rect 373660 402882 373716 402892
rect 383180 402724 383236 404460
rect 384860 403172 384916 408492
rect 393484 408324 393540 408334
rect 393148 405300 393204 405310
rect 391468 404964 391524 404974
rect 389676 404516 389732 404526
rect 384860 403106 384916 403116
rect 389452 404180 389508 404190
rect 383180 402658 383236 402668
rect 389452 402612 389508 404124
rect 389676 402948 389732 404460
rect 389900 404516 389956 404526
rect 389676 402882 389732 402892
rect 389788 403620 389844 403630
rect 389788 402724 389844 403564
rect 389900 403172 389956 404460
rect 390572 404404 390628 404414
rect 390572 403732 390628 404348
rect 390572 403666 390628 403676
rect 389900 403106 389956 403116
rect 391468 403060 391524 404908
rect 391468 402994 391524 403004
rect 393148 403060 393204 405244
rect 393484 403172 393540 408268
rect 479276 408100 479332 567308
rect 480508 410564 480564 573692
rect 480508 410498 480564 410508
rect 480620 410452 480676 575036
rect 496938 562350 497558 579922
rect 496938 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 497558 562350
rect 496938 562226 497558 562294
rect 496938 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 497558 562226
rect 496938 562102 497558 562170
rect 496938 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 497558 562102
rect 496938 561978 497558 562046
rect 496938 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 497558 561978
rect 486288 550350 486608 550384
rect 486288 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 486608 550350
rect 486288 550226 486608 550294
rect 486288 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 486608 550226
rect 486288 550102 486608 550170
rect 486288 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 486608 550102
rect 486288 549978 486608 550046
rect 486288 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 486608 549978
rect 486288 549888 486608 549922
rect 496938 544350 497558 561922
rect 496938 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 497558 544350
rect 496938 544226 497558 544294
rect 496938 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 497558 544226
rect 496938 544102 497558 544170
rect 496938 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 497558 544102
rect 496938 543978 497558 544046
rect 496938 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 497558 543978
rect 486288 532350 486608 532384
rect 486288 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 486608 532350
rect 486288 532226 486608 532294
rect 486288 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 486608 532226
rect 486288 532102 486608 532170
rect 486288 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 486608 532102
rect 486288 531978 486608 532046
rect 486288 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 486608 531978
rect 486288 531888 486608 531922
rect 496938 526350 497558 543922
rect 496938 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 497558 526350
rect 496938 526226 497558 526294
rect 496938 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 497558 526226
rect 496938 526102 497558 526170
rect 496938 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 497558 526102
rect 496938 525978 497558 526046
rect 496938 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 497558 525978
rect 486288 514350 486608 514384
rect 486288 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 486608 514350
rect 486288 514226 486608 514294
rect 486288 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 486608 514226
rect 486288 514102 486608 514170
rect 486288 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 486608 514102
rect 486288 513978 486608 514046
rect 486288 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 486608 513978
rect 486288 513888 486608 513922
rect 496938 508350 497558 525922
rect 496938 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 497558 508350
rect 496938 508226 497558 508294
rect 496938 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 497558 508226
rect 496938 508102 497558 508170
rect 496938 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 497558 508102
rect 496938 507978 497558 508046
rect 496938 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 497558 507978
rect 486288 496350 486608 496384
rect 486288 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 486608 496350
rect 486288 496226 486608 496294
rect 486288 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 486608 496226
rect 486288 496102 486608 496170
rect 486288 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 486608 496102
rect 486288 495978 486608 496046
rect 486288 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 486608 495978
rect 486288 495888 486608 495922
rect 496938 490350 497558 507922
rect 496938 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 497558 490350
rect 496938 490226 497558 490294
rect 496938 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 497558 490226
rect 496938 490102 497558 490170
rect 496938 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 497558 490102
rect 496938 489978 497558 490046
rect 496938 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 497558 489978
rect 486288 478350 486608 478384
rect 486288 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 486608 478350
rect 486288 478226 486608 478294
rect 486288 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 486608 478226
rect 486288 478102 486608 478170
rect 486288 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 486608 478102
rect 486288 477978 486608 478046
rect 486288 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 486608 477978
rect 486288 477888 486608 477922
rect 496938 472350 497558 489922
rect 496938 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 497558 472350
rect 496938 472226 497558 472294
rect 496938 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 497558 472226
rect 496938 472102 497558 472170
rect 496938 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 497558 472102
rect 496938 471978 497558 472046
rect 496938 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 497558 471978
rect 486288 460350 486608 460384
rect 486288 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 486608 460350
rect 486288 460226 486608 460294
rect 486288 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 486608 460226
rect 486288 460102 486608 460170
rect 486288 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 486608 460102
rect 486288 459978 486608 460046
rect 486288 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 486608 459978
rect 486288 459888 486608 459922
rect 496938 454350 497558 471922
rect 496938 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 497558 454350
rect 496938 454226 497558 454294
rect 496938 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 497558 454226
rect 496938 454102 497558 454170
rect 496938 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 497558 454102
rect 496938 453978 497558 454046
rect 496938 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 497558 453978
rect 486288 442350 486608 442384
rect 486288 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 486608 442350
rect 486288 442226 486608 442294
rect 486288 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 486608 442226
rect 486288 442102 486608 442170
rect 486288 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 486608 442102
rect 486288 441978 486608 442046
rect 486288 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 486608 441978
rect 486288 441888 486608 441922
rect 496938 436350 497558 453922
rect 496938 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 497558 436350
rect 496938 436226 497558 436294
rect 496938 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 497558 436226
rect 496938 436102 497558 436170
rect 496938 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 497558 436102
rect 496938 435978 497558 436046
rect 496938 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 497558 435978
rect 486288 424350 486608 424384
rect 486288 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 486608 424350
rect 486288 424226 486608 424294
rect 486288 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 486608 424226
rect 486288 424102 486608 424170
rect 486288 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 486608 424102
rect 486288 423978 486608 424046
rect 486288 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 486608 423978
rect 486288 423888 486608 423922
rect 480620 410386 480676 410396
rect 496938 418350 497558 435922
rect 496938 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 497558 418350
rect 496938 418226 497558 418294
rect 496938 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 497558 418226
rect 496938 418102 497558 418170
rect 496938 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 497558 418102
rect 496938 417978 497558 418046
rect 496938 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 497558 417978
rect 496412 409332 496468 409342
rect 496412 408538 496468 409276
rect 496412 408472 496468 408482
rect 479276 408034 479332 408044
rect 434588 406644 434644 406654
rect 403228 406196 403284 406206
rect 398188 405076 398244 405086
rect 393484 403106 393540 403116
rect 395836 404404 395892 404414
rect 393148 402994 393204 403004
rect 395836 402836 395892 404348
rect 398188 403732 398244 405020
rect 398300 404522 398692 404578
rect 398300 404516 398356 404522
rect 398300 404450 398356 404460
rect 398412 404404 398468 404414
rect 398412 404180 398468 404348
rect 398636 404404 398692 404522
rect 398636 404338 398692 404348
rect 398412 404114 398468 404124
rect 398188 403666 398244 403676
rect 403228 403172 403284 406140
rect 403228 403106 403284 403116
rect 434588 402948 434644 406588
rect 439068 404740 439124 404750
rect 439068 403956 439124 404684
rect 439068 403890 439124 403900
rect 447580 404292 447636 404302
rect 447580 403732 447636 404236
rect 447580 403666 447636 403676
rect 454972 404292 455028 404302
rect 454972 403060 455028 404236
rect 454972 402994 455028 403004
rect 496938 402950 497558 417922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 568350 501278 585922
rect 500658 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 501278 568350
rect 500658 568226 501278 568294
rect 500658 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 501278 568226
rect 500658 568102 501278 568170
rect 500658 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 501278 568102
rect 500658 567978 501278 568046
rect 500658 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 501278 567978
rect 500658 550350 501278 567922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 501648 562350 501968 562384
rect 501648 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 501968 562350
rect 501648 562226 501968 562294
rect 501648 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 501968 562226
rect 501648 562102 501968 562170
rect 501648 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 501968 562102
rect 501648 561978 501968 562046
rect 501648 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 501968 561978
rect 501648 561888 501968 561922
rect 527658 562350 528278 579922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 529676 576548 529732 576558
rect 529452 573300 529508 573310
rect 527658 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 528278 562350
rect 527658 562226 528278 562294
rect 527658 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 528278 562226
rect 527658 562102 528278 562170
rect 527658 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 528278 562102
rect 527658 561978 528278 562046
rect 527658 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 528278 561978
rect 500658 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 501278 550350
rect 500658 550226 501278 550294
rect 500658 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 501278 550226
rect 500658 550102 501278 550170
rect 500658 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 501278 550102
rect 500658 549978 501278 550046
rect 500658 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 501278 549978
rect 500658 532350 501278 549922
rect 517008 550350 517328 550384
rect 517008 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 517328 550350
rect 517008 550226 517328 550294
rect 517008 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 517328 550226
rect 517008 550102 517328 550170
rect 517008 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 517328 550102
rect 517008 549978 517328 550046
rect 517008 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 517328 549978
rect 517008 549888 517328 549922
rect 501648 544350 501968 544384
rect 501648 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 501968 544350
rect 501648 544226 501968 544294
rect 501648 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 501968 544226
rect 501648 544102 501968 544170
rect 501648 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 501968 544102
rect 501648 543978 501968 544046
rect 501648 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 501968 543978
rect 501648 543888 501968 543922
rect 527658 544350 528278 561922
rect 527658 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 528278 544350
rect 527658 544226 528278 544294
rect 527658 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 528278 544226
rect 527658 544102 528278 544170
rect 527658 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 528278 544102
rect 527658 543978 528278 544046
rect 527658 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 528278 543978
rect 500658 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 501278 532350
rect 500658 532226 501278 532294
rect 500658 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 501278 532226
rect 500658 532102 501278 532170
rect 500658 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 501278 532102
rect 500658 531978 501278 532046
rect 500658 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 501278 531978
rect 500658 514350 501278 531922
rect 517008 532350 517328 532384
rect 517008 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 517328 532350
rect 517008 532226 517328 532294
rect 517008 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 517328 532226
rect 517008 532102 517328 532170
rect 517008 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 517328 532102
rect 517008 531978 517328 532046
rect 517008 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 517328 531978
rect 517008 531888 517328 531922
rect 501648 526350 501968 526384
rect 501648 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 501968 526350
rect 501648 526226 501968 526294
rect 501648 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 501968 526226
rect 501648 526102 501968 526170
rect 501648 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 501968 526102
rect 501648 525978 501968 526046
rect 501648 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 501968 525978
rect 501648 525888 501968 525922
rect 527658 526350 528278 543922
rect 527658 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 528278 526350
rect 527658 526226 528278 526294
rect 527658 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 528278 526226
rect 527658 526102 528278 526170
rect 527658 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 528278 526102
rect 527658 525978 528278 526046
rect 527658 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 528278 525978
rect 500658 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 501278 514350
rect 500658 514226 501278 514294
rect 500658 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 501278 514226
rect 500658 514102 501278 514170
rect 500658 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 501278 514102
rect 500658 513978 501278 514046
rect 500658 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 501278 513978
rect 500658 496350 501278 513922
rect 517008 514350 517328 514384
rect 517008 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 517328 514350
rect 517008 514226 517328 514294
rect 517008 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 517328 514226
rect 517008 514102 517328 514170
rect 517008 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 517328 514102
rect 517008 513978 517328 514046
rect 517008 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 517328 513978
rect 517008 513888 517328 513922
rect 501648 508350 501968 508384
rect 501648 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 501968 508350
rect 501648 508226 501968 508294
rect 501648 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 501968 508226
rect 501648 508102 501968 508170
rect 501648 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 501968 508102
rect 501648 507978 501968 508046
rect 501648 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 501968 507978
rect 501648 507888 501968 507922
rect 527658 508350 528278 525922
rect 527658 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 528278 508350
rect 527658 508226 528278 508294
rect 527658 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 528278 508226
rect 527658 508102 528278 508170
rect 527658 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 528278 508102
rect 527658 507978 528278 508046
rect 527658 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 528278 507978
rect 500658 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 501278 496350
rect 500658 496226 501278 496294
rect 500658 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 501278 496226
rect 500658 496102 501278 496170
rect 500658 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 501278 496102
rect 500658 495978 501278 496046
rect 500658 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 501278 495978
rect 500658 478350 501278 495922
rect 517008 496350 517328 496384
rect 517008 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 517328 496350
rect 517008 496226 517328 496294
rect 517008 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 517328 496226
rect 517008 496102 517328 496170
rect 517008 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 517328 496102
rect 517008 495978 517328 496046
rect 517008 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 517328 495978
rect 517008 495888 517328 495922
rect 501648 490350 501968 490384
rect 501648 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 501968 490350
rect 501648 490226 501968 490294
rect 501648 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 501968 490226
rect 501648 490102 501968 490170
rect 501648 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 501968 490102
rect 501648 489978 501968 490046
rect 501648 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 501968 489978
rect 501648 489888 501968 489922
rect 527658 490350 528278 507922
rect 529340 568484 529396 568494
rect 529340 494564 529396 568428
rect 529452 508676 529508 573244
rect 529564 572068 529620 572078
rect 529564 532196 529620 572012
rect 529564 532130 529620 532140
rect 529452 508610 529508 508620
rect 529340 494498 529396 494508
rect 527658 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 528278 490350
rect 527658 490226 528278 490294
rect 527658 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 528278 490226
rect 527658 490102 528278 490170
rect 527658 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 528278 490102
rect 527658 489978 528278 490046
rect 527658 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 528278 489978
rect 500658 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 501278 478350
rect 500658 478226 501278 478294
rect 500658 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 501278 478226
rect 500658 478102 501278 478170
rect 500658 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 501278 478102
rect 500658 477978 501278 478046
rect 500658 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 501278 477978
rect 500658 460350 501278 477922
rect 517008 478350 517328 478384
rect 517008 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 517328 478350
rect 517008 478226 517328 478294
rect 517008 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 517328 478226
rect 517008 478102 517328 478170
rect 517008 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 517328 478102
rect 517008 477978 517328 478046
rect 517008 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 517328 477978
rect 517008 477888 517328 477922
rect 501648 472350 501968 472384
rect 501648 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 501968 472350
rect 501648 472226 501968 472294
rect 501648 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 501968 472226
rect 501648 472102 501968 472170
rect 501648 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 501968 472102
rect 501648 471978 501968 472046
rect 501648 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 501968 471978
rect 501648 471888 501968 471922
rect 527658 472350 528278 489922
rect 529676 489860 529732 576492
rect 529676 489794 529732 489804
rect 531378 568350 531998 585922
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 531378 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 531998 568350
rect 531378 568226 531998 568294
rect 531378 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 531998 568226
rect 531378 568102 531998 568170
rect 531378 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 531998 568102
rect 531378 567978 531998 568046
rect 531378 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 531998 567978
rect 531378 550350 531998 567922
rect 532588 576436 532644 576446
rect 532588 560420 532644 576380
rect 532812 574868 532868 574878
rect 532588 560354 532644 560364
rect 532700 570164 532756 570174
rect 531378 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 531998 550350
rect 531378 550226 531998 550294
rect 531378 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 531998 550226
rect 531378 550102 531998 550170
rect 531378 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 531998 550102
rect 531378 549978 531998 550046
rect 531378 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 531998 549978
rect 531378 532350 531998 549922
rect 532700 541604 532756 570108
rect 532812 565124 532868 574812
rect 533260 571844 533316 571854
rect 533036 570276 533092 570286
rect 532812 565058 532868 565068
rect 532924 568596 532980 568606
rect 532812 564900 532868 564910
rect 532812 546308 532868 564844
rect 532924 551012 532980 568540
rect 533036 555716 533092 570220
rect 533036 555650 533092 555660
rect 533148 566218 533204 566228
rect 532924 550946 532980 550956
rect 532812 546242 532868 546252
rect 532700 541538 532756 541548
rect 531378 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 531998 532350
rect 531378 532226 531998 532294
rect 531378 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 531998 532226
rect 531378 532102 531998 532170
rect 531378 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 531998 532102
rect 531378 531978 531998 532046
rect 531378 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 531998 531978
rect 531378 514350 531998 531922
rect 531378 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 531998 514350
rect 531378 514226 531998 514294
rect 531378 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 531998 514226
rect 531378 514102 531998 514170
rect 531378 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 531998 514102
rect 531378 513978 531998 514046
rect 531378 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 531998 513978
rect 531378 496350 531998 513922
rect 531378 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 531998 496350
rect 531378 496226 531998 496294
rect 531378 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 531998 496226
rect 531378 496102 531998 496170
rect 531378 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 531998 496102
rect 531378 495978 531998 496046
rect 531378 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 531998 495978
rect 527658 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 528278 472350
rect 527658 472226 528278 472294
rect 527658 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 528278 472226
rect 527658 472102 528278 472170
rect 527658 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 528278 472102
rect 527658 471978 528278 472046
rect 527658 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 528278 471978
rect 500658 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 501278 460350
rect 500658 460226 501278 460294
rect 500658 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 501278 460226
rect 500658 460102 501278 460170
rect 500658 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 501278 460102
rect 500658 459978 501278 460046
rect 500658 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 501278 459978
rect 500658 442350 501278 459922
rect 517008 460350 517328 460384
rect 517008 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 517328 460350
rect 517008 460226 517328 460294
rect 517008 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 517328 460226
rect 517008 460102 517328 460170
rect 517008 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 517328 460102
rect 517008 459978 517328 460046
rect 517008 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 517328 459978
rect 517008 459888 517328 459922
rect 501648 454350 501968 454384
rect 501648 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 501968 454350
rect 501648 454226 501968 454294
rect 501648 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 501968 454226
rect 501648 454102 501968 454170
rect 501648 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 501968 454102
rect 501648 453978 501968 454046
rect 501648 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 501968 453978
rect 501648 453888 501968 453922
rect 527658 454350 528278 471922
rect 527658 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 528278 454350
rect 527658 454226 528278 454294
rect 527658 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 528278 454226
rect 527658 454102 528278 454170
rect 527658 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 528278 454102
rect 527658 453978 528278 454046
rect 527658 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 528278 453978
rect 500658 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 501278 442350
rect 500658 442226 501278 442294
rect 500658 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 501278 442226
rect 500658 442102 501278 442170
rect 500658 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 501278 442102
rect 500658 441978 501278 442046
rect 500658 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 501278 441978
rect 500658 424350 501278 441922
rect 517008 442350 517328 442384
rect 517008 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 517328 442350
rect 517008 442226 517328 442294
rect 517008 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 517328 442226
rect 517008 442102 517328 442170
rect 517008 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 517328 442102
rect 517008 441978 517328 442046
rect 517008 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 517328 441978
rect 517008 441888 517328 441922
rect 501648 436350 501968 436384
rect 501648 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 501968 436350
rect 501648 436226 501968 436294
rect 501648 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 501968 436226
rect 501648 436102 501968 436170
rect 501648 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 501968 436102
rect 501648 435978 501968 436046
rect 501648 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 501968 435978
rect 501648 435888 501968 435922
rect 527658 436350 528278 453922
rect 527658 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 528278 436350
rect 527658 436226 528278 436294
rect 527658 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 528278 436226
rect 527658 436102 528278 436170
rect 527658 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 528278 436102
rect 527658 435978 528278 436046
rect 527658 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 528278 435978
rect 500658 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 501278 424350
rect 500658 424226 501278 424294
rect 500658 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 501278 424226
rect 500658 424102 501278 424170
rect 500658 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 501278 424102
rect 500658 423978 501278 424046
rect 500658 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 501278 423978
rect 499324 410338 499380 410348
rect 499324 406644 499380 410282
rect 499324 406578 499380 406588
rect 500658 406350 501278 423922
rect 517008 424350 517328 424384
rect 517008 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 517328 424350
rect 517008 424226 517328 424294
rect 517008 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 517328 424226
rect 517008 424102 517328 424170
rect 517008 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 517328 424102
rect 517008 423978 517328 424046
rect 517008 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 517328 423978
rect 517008 423888 517328 423922
rect 501648 418350 501968 418384
rect 501648 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 501968 418350
rect 501648 418226 501968 418294
rect 501648 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 501968 418226
rect 501648 418102 501968 418170
rect 501648 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 501968 418102
rect 501648 417978 501968 418046
rect 501648 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 501968 417978
rect 501648 417888 501968 417922
rect 527658 418350 528278 435922
rect 527658 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 528278 418350
rect 527658 418226 528278 418294
rect 527658 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 528278 418226
rect 527658 418102 528278 418170
rect 527658 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 528278 418102
rect 527658 417978 528278 418046
rect 527658 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 528278 417978
rect 514108 408358 514164 408368
rect 500658 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 501278 406350
rect 500658 406226 501278 406294
rect 500658 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 501278 406226
rect 500658 406102 501278 406170
rect 500658 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 501278 406102
rect 500658 405978 501278 406046
rect 500658 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 501278 405978
rect 500658 402950 501278 405922
rect 501564 406644 501620 406654
rect 434588 402882 434644 402892
rect 395836 402770 395892 402780
rect 389788 402658 389844 402668
rect 501564 402724 501620 406588
rect 501564 402658 501620 402668
rect 511868 406644 511924 406654
rect 389452 402546 389508 402556
rect 511868 402598 511924 406588
rect 514108 406644 514164 408302
rect 514108 406578 514164 406588
rect 517020 406644 517076 406654
rect 511868 402532 511924 402542
rect 517020 402418 517076 406588
rect 522172 406644 522228 406654
rect 522172 404218 522228 406588
rect 522172 404152 522228 404162
rect 527436 404852 527492 404862
rect 517020 402352 517076 402362
rect 527436 402388 527492 404796
rect 527658 402950 528278 417922
rect 531378 478350 531998 495922
rect 531378 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 531998 478350
rect 531378 478226 531998 478294
rect 531378 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 531998 478226
rect 531378 478102 531998 478170
rect 531378 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 531998 478102
rect 531378 477978 531998 478046
rect 531378 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 531998 477978
rect 531378 460350 531998 477922
rect 533148 466340 533204 566162
rect 533260 564900 533316 571788
rect 533260 564834 533316 564844
rect 533148 466274 533204 466284
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 531378 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 531998 460350
rect 531378 460226 531998 460294
rect 531378 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 531998 460226
rect 531378 460102 531998 460170
rect 531378 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 531998 460102
rect 531378 459978 531998 460046
rect 531378 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 531998 459978
rect 531378 442350 531998 459922
rect 531378 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 531998 442350
rect 531378 442226 531998 442294
rect 531378 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 531998 442226
rect 531378 442102 531998 442170
rect 531378 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 531998 442102
rect 531378 441978 531998 442046
rect 531378 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 531998 441978
rect 531378 424350 531998 441922
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 531378 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 531998 424350
rect 531378 424226 531998 424294
rect 531378 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 531998 424226
rect 531378 424102 531998 424170
rect 531378 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 531998 424102
rect 531378 423978 531998 424046
rect 531378 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 531998 423978
rect 528892 407278 528948 407288
rect 528892 406644 528948 407222
rect 528892 406578 528948 406588
rect 531378 406350 531998 423922
rect 532588 428708 532644 428718
rect 532588 409078 532644 428652
rect 532588 409012 532644 409022
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 558236 408178 558292 408188
rect 543676 407098 543732 407108
rect 543676 406644 543732 407042
rect 543676 406578 543732 406588
rect 551068 406918 551124 406928
rect 551068 406644 551124 406862
rect 551068 406578 551124 406588
rect 558236 406644 558292 408122
rect 558236 406578 558292 406588
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 402950 531998 405922
rect 558378 402950 558998 417922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 589098 580350 589718 596784
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 590492 588644 590548 588654
rect 590492 573778 590548 588588
rect 590492 573712 590548 573722
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 590604 571258 590660 571268
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 590492 569818 590548 569828
rect 590492 469924 590548 569762
rect 590604 496356 590660 571202
rect 590828 569638 590884 569648
rect 590716 568148 590772 568158
rect 590716 509572 590772 568092
rect 590828 549220 590884 569582
rect 590828 549154 590884 549164
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 590716 509506 590772 509516
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 590604 496290 590660 496300
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 590492 469858 590548 469868
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 580636 407638 580692 407648
rect 580636 406644 580692 407582
rect 580636 406578 580692 406588
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 402950 562718 405922
rect 565852 404292 565908 404302
rect 565852 403138 565908 404236
rect 565852 403072 565908 403082
rect 582092 404038 582148 404048
rect 372764 402322 372820 402332
rect 527436 402322 527492 402332
rect 367836 401452 367892 401462
rect 346108 401092 346164 401102
rect 341516 400552 341572 400562
rect 344448 400350 344768 400384
rect 344448 400294 344518 400350
rect 344574 400294 344642 400350
rect 344698 400294 344768 400350
rect 344448 400226 344768 400294
rect 344448 400170 344518 400226
rect 344574 400170 344642 400226
rect 344698 400170 344768 400226
rect 344448 400102 344768 400170
rect 344448 400046 344518 400102
rect 344574 400046 344642 400102
rect 344698 400046 344768 400102
rect 344448 399978 344768 400046
rect 344448 399922 344518 399978
rect 344574 399922 344642 399978
rect 344698 399922 344768 399978
rect 344448 399888 344768 399922
rect 375168 400350 375488 400384
rect 375168 400294 375238 400350
rect 375294 400294 375362 400350
rect 375418 400294 375488 400350
rect 375168 400226 375488 400294
rect 375168 400170 375238 400226
rect 375294 400170 375362 400226
rect 375418 400170 375488 400226
rect 375168 400102 375488 400170
rect 375168 400046 375238 400102
rect 375294 400046 375362 400102
rect 375418 400046 375488 400102
rect 375168 399978 375488 400046
rect 375168 399922 375238 399978
rect 375294 399922 375362 399978
rect 375418 399922 375488 399978
rect 375168 399888 375488 399922
rect 405888 400350 406208 400384
rect 405888 400294 405958 400350
rect 406014 400294 406082 400350
rect 406138 400294 406208 400350
rect 405888 400226 406208 400294
rect 405888 400170 405958 400226
rect 406014 400170 406082 400226
rect 406138 400170 406208 400226
rect 405888 400102 406208 400170
rect 405888 400046 405958 400102
rect 406014 400046 406082 400102
rect 406138 400046 406208 400102
rect 405888 399978 406208 400046
rect 405888 399922 405958 399978
rect 406014 399922 406082 399978
rect 406138 399922 406208 399978
rect 405888 399888 406208 399922
rect 436608 400350 436928 400384
rect 436608 400294 436678 400350
rect 436734 400294 436802 400350
rect 436858 400294 436928 400350
rect 436608 400226 436928 400294
rect 436608 400170 436678 400226
rect 436734 400170 436802 400226
rect 436858 400170 436928 400226
rect 436608 400102 436928 400170
rect 436608 400046 436678 400102
rect 436734 400046 436802 400102
rect 436858 400046 436928 400102
rect 436608 399978 436928 400046
rect 436608 399922 436678 399978
rect 436734 399922 436802 399978
rect 436858 399922 436928 399978
rect 436608 399888 436928 399922
rect 467328 400350 467648 400384
rect 467328 400294 467398 400350
rect 467454 400294 467522 400350
rect 467578 400294 467648 400350
rect 467328 400226 467648 400294
rect 467328 400170 467398 400226
rect 467454 400170 467522 400226
rect 467578 400170 467648 400226
rect 467328 400102 467648 400170
rect 467328 400046 467398 400102
rect 467454 400046 467522 400102
rect 467578 400046 467648 400102
rect 467328 399978 467648 400046
rect 467328 399922 467398 399978
rect 467454 399922 467522 399978
rect 467578 399922 467648 399978
rect 467328 399888 467648 399922
rect 498048 400350 498368 400384
rect 498048 400294 498118 400350
rect 498174 400294 498242 400350
rect 498298 400294 498368 400350
rect 498048 400226 498368 400294
rect 498048 400170 498118 400226
rect 498174 400170 498242 400226
rect 498298 400170 498368 400226
rect 498048 400102 498368 400170
rect 498048 400046 498118 400102
rect 498174 400046 498242 400102
rect 498298 400046 498368 400102
rect 498048 399978 498368 400046
rect 498048 399922 498118 399978
rect 498174 399922 498242 399978
rect 498298 399922 498368 399978
rect 498048 399888 498368 399922
rect 528768 400350 529088 400384
rect 528768 400294 528838 400350
rect 528894 400294 528962 400350
rect 529018 400294 529088 400350
rect 528768 400226 529088 400294
rect 528768 400170 528838 400226
rect 528894 400170 528962 400226
rect 529018 400170 529088 400226
rect 528768 400102 529088 400170
rect 528768 400046 528838 400102
rect 528894 400046 528962 400102
rect 529018 400046 529088 400102
rect 528768 399978 529088 400046
rect 528768 399922 528838 399978
rect 528894 399922 528962 399978
rect 529018 399922 529088 399978
rect 528768 399888 529088 399922
rect 559488 400350 559808 400384
rect 559488 400294 559558 400350
rect 559614 400294 559682 400350
rect 559738 400294 559808 400350
rect 559488 400226 559808 400294
rect 559488 400170 559558 400226
rect 559614 400170 559682 400226
rect 559738 400170 559808 400226
rect 559488 400102 559808 400170
rect 559488 400046 559558 400102
rect 559614 400046 559682 400102
rect 559738 400046 559808 400102
rect 559488 399978 559808 400046
rect 559488 399922 559558 399978
rect 559614 399922 559682 399978
rect 559738 399922 559808 399978
rect 559488 399888 559808 399922
rect 341180 399652 341236 399662
rect 340620 396452 340900 396508
rect 340620 395668 340676 396452
rect 340620 395602 340676 395612
rect 582092 391438 582148 403982
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 582092 391372 582148 391382
rect 587132 391438 587188 391448
rect 359808 388350 360128 388384
rect 359808 388294 359878 388350
rect 359934 388294 360002 388350
rect 360058 388294 360128 388350
rect 359808 388226 360128 388294
rect 359808 388170 359878 388226
rect 359934 388170 360002 388226
rect 360058 388170 360128 388226
rect 359808 388102 360128 388170
rect 359808 388046 359878 388102
rect 359934 388046 360002 388102
rect 360058 388046 360128 388102
rect 359808 387978 360128 388046
rect 359808 387922 359878 387978
rect 359934 387922 360002 387978
rect 360058 387922 360128 387978
rect 359808 387888 360128 387922
rect 390528 388350 390848 388384
rect 390528 388294 390598 388350
rect 390654 388294 390722 388350
rect 390778 388294 390848 388350
rect 390528 388226 390848 388294
rect 390528 388170 390598 388226
rect 390654 388170 390722 388226
rect 390778 388170 390848 388226
rect 390528 388102 390848 388170
rect 390528 388046 390598 388102
rect 390654 388046 390722 388102
rect 390778 388046 390848 388102
rect 390528 387978 390848 388046
rect 390528 387922 390598 387978
rect 390654 387922 390722 387978
rect 390778 387922 390848 387978
rect 390528 387888 390848 387922
rect 421248 388350 421568 388384
rect 421248 388294 421318 388350
rect 421374 388294 421442 388350
rect 421498 388294 421568 388350
rect 421248 388226 421568 388294
rect 421248 388170 421318 388226
rect 421374 388170 421442 388226
rect 421498 388170 421568 388226
rect 421248 388102 421568 388170
rect 421248 388046 421318 388102
rect 421374 388046 421442 388102
rect 421498 388046 421568 388102
rect 421248 387978 421568 388046
rect 421248 387922 421318 387978
rect 421374 387922 421442 387978
rect 421498 387922 421568 387978
rect 421248 387888 421568 387922
rect 451968 388350 452288 388384
rect 451968 388294 452038 388350
rect 452094 388294 452162 388350
rect 452218 388294 452288 388350
rect 451968 388226 452288 388294
rect 451968 388170 452038 388226
rect 452094 388170 452162 388226
rect 452218 388170 452288 388226
rect 451968 388102 452288 388170
rect 451968 388046 452038 388102
rect 452094 388046 452162 388102
rect 452218 388046 452288 388102
rect 451968 387978 452288 388046
rect 451968 387922 452038 387978
rect 452094 387922 452162 387978
rect 452218 387922 452288 387978
rect 451968 387888 452288 387922
rect 482688 388350 483008 388384
rect 482688 388294 482758 388350
rect 482814 388294 482882 388350
rect 482938 388294 483008 388350
rect 482688 388226 483008 388294
rect 482688 388170 482758 388226
rect 482814 388170 482882 388226
rect 482938 388170 483008 388226
rect 482688 388102 483008 388170
rect 482688 388046 482758 388102
rect 482814 388046 482882 388102
rect 482938 388046 483008 388102
rect 482688 387978 483008 388046
rect 482688 387922 482758 387978
rect 482814 387922 482882 387978
rect 482938 387922 483008 387978
rect 482688 387888 483008 387922
rect 513408 388350 513728 388384
rect 513408 388294 513478 388350
rect 513534 388294 513602 388350
rect 513658 388294 513728 388350
rect 513408 388226 513728 388294
rect 513408 388170 513478 388226
rect 513534 388170 513602 388226
rect 513658 388170 513728 388226
rect 513408 388102 513728 388170
rect 513408 388046 513478 388102
rect 513534 388046 513602 388102
rect 513658 388046 513728 388102
rect 513408 387978 513728 388046
rect 513408 387922 513478 387978
rect 513534 387922 513602 387978
rect 513658 387922 513728 387978
rect 513408 387888 513728 387922
rect 544128 388350 544448 388384
rect 544128 388294 544198 388350
rect 544254 388294 544322 388350
rect 544378 388294 544448 388350
rect 544128 388226 544448 388294
rect 544128 388170 544198 388226
rect 544254 388170 544322 388226
rect 544378 388170 544448 388226
rect 544128 388102 544448 388170
rect 544128 388046 544198 388102
rect 544254 388046 544322 388102
rect 544378 388046 544448 388102
rect 544128 387978 544448 388046
rect 544128 387922 544198 387978
rect 544254 387922 544322 387978
rect 544378 387922 544448 387978
rect 544128 387888 544448 387922
rect 574848 388350 575168 388384
rect 574848 388294 574918 388350
rect 574974 388294 575042 388350
rect 575098 388294 575168 388350
rect 574848 388226 575168 388294
rect 574848 388170 574918 388226
rect 574974 388170 575042 388226
rect 575098 388170 575168 388226
rect 574848 388102 575168 388170
rect 574848 388046 574918 388102
rect 574974 388046 575042 388102
rect 575098 388046 575168 388102
rect 574848 387978 575168 388046
rect 574848 387922 574918 387978
rect 574974 387922 575042 387978
rect 575098 387922 575168 387978
rect 574848 387888 575168 387922
rect 339052 382498 339108 382508
rect 339500 386820 339556 386830
rect 338604 382386 338660 382396
rect 338492 379586 338548 379596
rect 338044 362404 338100 362414
rect 337820 300738 337876 300748
rect 337932 330148 337988 330158
rect 337708 277778 337764 277788
rect 337820 300580 337876 300590
rect 337708 254660 337764 254670
rect 337708 243796 337764 254604
rect 337820 253652 337876 300524
rect 337932 264628 337988 330092
rect 338044 311698 338100 362348
rect 338604 327460 338660 327470
rect 338044 311632 338100 311642
rect 338492 325668 338548 325678
rect 338156 311332 338212 311342
rect 337932 264562 337988 264572
rect 338044 307748 338100 307758
rect 338044 254996 338100 307692
rect 338156 286804 338212 311276
rect 338156 286738 338212 286748
rect 338268 290388 338324 290398
rect 338044 254930 338100 254940
rect 338156 268100 338212 268110
rect 337820 253586 337876 253596
rect 337708 243730 337764 243740
rect 337932 248724 337988 248734
rect 337820 243572 337876 243582
rect 337596 147858 337652 147868
rect 337708 198324 337764 198334
rect 337260 139122 337316 139132
rect 337708 132238 337764 198268
rect 337820 179732 337876 243516
rect 337932 189812 337988 248668
rect 338156 240772 338212 268044
rect 338268 248724 338324 290332
rect 338268 248658 338324 248668
rect 338380 259700 338436 259710
rect 338380 240958 338436 259644
rect 338380 240892 338436 240902
rect 338156 240706 338212 240716
rect 337932 189746 337988 189756
rect 337820 179666 337876 179676
rect 338492 139076 338548 325612
rect 338604 142498 338660 327404
rect 338716 324772 338772 324782
rect 338716 145378 338772 324716
rect 339388 309540 339444 309550
rect 338940 267652 338996 267662
rect 338828 249418 338884 249428
rect 338828 152852 338884 249362
rect 338940 242004 338996 267596
rect 338940 241938 338996 241948
rect 339276 247044 339332 247054
rect 338828 152786 338884 152796
rect 338940 189028 338996 189038
rect 338716 145312 338772 145322
rect 338604 142432 338660 142442
rect 338940 142324 338996 188972
rect 338940 142258 338996 142268
rect 338492 139010 338548 139020
rect 337708 132172 337764 132182
rect 337148 127652 337204 127662
rect 337148 127558 337204 127596
rect 337148 127492 337204 127502
rect 337036 99026 337092 99036
rect 335580 47842 335636 47852
rect 335356 44482 335412 44492
rect 335132 42802 335188 42812
rect 334236 33532 334292 33542
rect 330764 31732 330820 31742
rect 339276 30178 339332 246988
rect 339388 208348 339444 309484
rect 339500 278180 339556 386764
rect 344448 382350 344768 382384
rect 344448 382294 344518 382350
rect 344574 382294 344642 382350
rect 344698 382294 344768 382350
rect 344448 382226 344768 382294
rect 344448 382170 344518 382226
rect 344574 382170 344642 382226
rect 344698 382170 344768 382226
rect 344448 382102 344768 382170
rect 344448 382046 344518 382102
rect 344574 382046 344642 382102
rect 344698 382046 344768 382102
rect 344448 381978 344768 382046
rect 344448 381922 344518 381978
rect 344574 381922 344642 381978
rect 344698 381922 344768 381978
rect 344448 381888 344768 381922
rect 375168 382350 375488 382384
rect 375168 382294 375238 382350
rect 375294 382294 375362 382350
rect 375418 382294 375488 382350
rect 375168 382226 375488 382294
rect 375168 382170 375238 382226
rect 375294 382170 375362 382226
rect 375418 382170 375488 382226
rect 375168 382102 375488 382170
rect 375168 382046 375238 382102
rect 375294 382046 375362 382102
rect 375418 382046 375488 382102
rect 375168 381978 375488 382046
rect 375168 381922 375238 381978
rect 375294 381922 375362 381978
rect 375418 381922 375488 381978
rect 375168 381888 375488 381922
rect 405888 382350 406208 382384
rect 405888 382294 405958 382350
rect 406014 382294 406082 382350
rect 406138 382294 406208 382350
rect 405888 382226 406208 382294
rect 405888 382170 405958 382226
rect 406014 382170 406082 382226
rect 406138 382170 406208 382226
rect 405888 382102 406208 382170
rect 405888 382046 405958 382102
rect 406014 382046 406082 382102
rect 406138 382046 406208 382102
rect 405888 381978 406208 382046
rect 405888 381922 405958 381978
rect 406014 381922 406082 381978
rect 406138 381922 406208 381978
rect 405888 381888 406208 381922
rect 436608 382350 436928 382384
rect 436608 382294 436678 382350
rect 436734 382294 436802 382350
rect 436858 382294 436928 382350
rect 436608 382226 436928 382294
rect 436608 382170 436678 382226
rect 436734 382170 436802 382226
rect 436858 382170 436928 382226
rect 436608 382102 436928 382170
rect 436608 382046 436678 382102
rect 436734 382046 436802 382102
rect 436858 382046 436928 382102
rect 436608 381978 436928 382046
rect 436608 381922 436678 381978
rect 436734 381922 436802 381978
rect 436858 381922 436928 381978
rect 436608 381888 436928 381922
rect 467328 382350 467648 382384
rect 467328 382294 467398 382350
rect 467454 382294 467522 382350
rect 467578 382294 467648 382350
rect 467328 382226 467648 382294
rect 467328 382170 467398 382226
rect 467454 382170 467522 382226
rect 467578 382170 467648 382226
rect 467328 382102 467648 382170
rect 467328 382046 467398 382102
rect 467454 382046 467522 382102
rect 467578 382046 467648 382102
rect 467328 381978 467648 382046
rect 467328 381922 467398 381978
rect 467454 381922 467522 381978
rect 467578 381922 467648 381978
rect 467328 381888 467648 381922
rect 498048 382350 498368 382384
rect 498048 382294 498118 382350
rect 498174 382294 498242 382350
rect 498298 382294 498368 382350
rect 498048 382226 498368 382294
rect 498048 382170 498118 382226
rect 498174 382170 498242 382226
rect 498298 382170 498368 382226
rect 498048 382102 498368 382170
rect 498048 382046 498118 382102
rect 498174 382046 498242 382102
rect 498298 382046 498368 382102
rect 498048 381978 498368 382046
rect 498048 381922 498118 381978
rect 498174 381922 498242 381978
rect 498298 381922 498368 381978
rect 498048 381888 498368 381922
rect 528768 382350 529088 382384
rect 528768 382294 528838 382350
rect 528894 382294 528962 382350
rect 529018 382294 529088 382350
rect 528768 382226 529088 382294
rect 528768 382170 528838 382226
rect 528894 382170 528962 382226
rect 529018 382170 529088 382226
rect 528768 382102 529088 382170
rect 528768 382046 528838 382102
rect 528894 382046 528962 382102
rect 529018 382046 529088 382102
rect 528768 381978 529088 382046
rect 528768 381922 528838 381978
rect 528894 381922 528962 381978
rect 529018 381922 529088 381978
rect 528768 381888 529088 381922
rect 559488 382350 559808 382384
rect 559488 382294 559558 382350
rect 559614 382294 559682 382350
rect 559738 382294 559808 382350
rect 559488 382226 559808 382294
rect 559488 382170 559558 382226
rect 559614 382170 559682 382226
rect 559738 382170 559808 382226
rect 559488 382102 559808 382170
rect 559488 382046 559558 382102
rect 559614 382046 559682 382102
rect 559738 382046 559808 382102
rect 559488 381978 559808 382046
rect 559488 381922 559558 381978
rect 559614 381922 559682 381978
rect 559738 381922 559808 381978
rect 559488 381888 559808 381922
rect 587132 377412 587188 391382
rect 587132 377346 587188 377356
rect 589098 382350 589718 399922
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 340508 371364 340564 371374
rect 339500 278114 339556 278124
rect 340172 312228 340228 312238
rect 339500 257124 339556 257134
rect 339500 246932 339556 257068
rect 339500 246866 339556 246876
rect 339948 248612 340004 248622
rect 339388 208292 339556 208348
rect 339388 197652 339444 197662
rect 339388 197316 339444 197596
rect 339388 197250 339444 197260
rect 339500 197204 339556 208292
rect 339500 197138 339556 197148
rect 339948 135492 340004 248556
rect 340060 197316 340116 197326
rect 340060 160858 340116 197260
rect 340060 160792 340116 160802
rect 339948 135426 340004 135436
rect 339276 30112 339332 30122
rect 340172 21588 340228 312172
rect 340284 310436 340340 310446
rect 340284 22820 340340 310380
rect 340396 294756 340452 294766
rect 340396 294598 340452 294700
rect 340396 294532 340452 294542
rect 340396 283798 340452 283808
rect 340396 275268 340452 283742
rect 340396 275202 340452 275212
rect 340284 22754 340340 22764
rect 340396 264740 340452 264750
rect 340172 21522 340228 21532
rect 340396 21476 340452 264684
rect 340508 157618 340564 371308
rect 359808 370350 360128 370384
rect 359808 370294 359878 370350
rect 359934 370294 360002 370350
rect 360058 370294 360128 370350
rect 359808 370226 360128 370294
rect 359808 370170 359878 370226
rect 359934 370170 360002 370226
rect 360058 370170 360128 370226
rect 359808 370102 360128 370170
rect 359808 370046 359878 370102
rect 359934 370046 360002 370102
rect 360058 370046 360128 370102
rect 359808 369978 360128 370046
rect 359808 369922 359878 369978
rect 359934 369922 360002 369978
rect 360058 369922 360128 369978
rect 359808 369888 360128 369922
rect 390528 370350 390848 370384
rect 390528 370294 390598 370350
rect 390654 370294 390722 370350
rect 390778 370294 390848 370350
rect 390528 370226 390848 370294
rect 390528 370170 390598 370226
rect 390654 370170 390722 370226
rect 390778 370170 390848 370226
rect 390528 370102 390848 370170
rect 390528 370046 390598 370102
rect 390654 370046 390722 370102
rect 390778 370046 390848 370102
rect 390528 369978 390848 370046
rect 390528 369922 390598 369978
rect 390654 369922 390722 369978
rect 390778 369922 390848 369978
rect 390528 369888 390848 369922
rect 421248 370350 421568 370384
rect 421248 370294 421318 370350
rect 421374 370294 421442 370350
rect 421498 370294 421568 370350
rect 421248 370226 421568 370294
rect 421248 370170 421318 370226
rect 421374 370170 421442 370226
rect 421498 370170 421568 370226
rect 421248 370102 421568 370170
rect 421248 370046 421318 370102
rect 421374 370046 421442 370102
rect 421498 370046 421568 370102
rect 421248 369978 421568 370046
rect 421248 369922 421318 369978
rect 421374 369922 421442 369978
rect 421498 369922 421568 369978
rect 421248 369888 421568 369922
rect 451968 370350 452288 370384
rect 451968 370294 452038 370350
rect 452094 370294 452162 370350
rect 452218 370294 452288 370350
rect 451968 370226 452288 370294
rect 451968 370170 452038 370226
rect 452094 370170 452162 370226
rect 452218 370170 452288 370226
rect 451968 370102 452288 370170
rect 451968 370046 452038 370102
rect 452094 370046 452162 370102
rect 452218 370046 452288 370102
rect 451968 369978 452288 370046
rect 451968 369922 452038 369978
rect 452094 369922 452162 369978
rect 452218 369922 452288 369978
rect 451968 369888 452288 369922
rect 482688 370350 483008 370384
rect 482688 370294 482758 370350
rect 482814 370294 482882 370350
rect 482938 370294 483008 370350
rect 482688 370226 483008 370294
rect 482688 370170 482758 370226
rect 482814 370170 482882 370226
rect 482938 370170 483008 370226
rect 482688 370102 483008 370170
rect 482688 370046 482758 370102
rect 482814 370046 482882 370102
rect 482938 370046 483008 370102
rect 482688 369978 483008 370046
rect 482688 369922 482758 369978
rect 482814 369922 482882 369978
rect 482938 369922 483008 369978
rect 482688 369888 483008 369922
rect 513408 370350 513728 370384
rect 513408 370294 513478 370350
rect 513534 370294 513602 370350
rect 513658 370294 513728 370350
rect 513408 370226 513728 370294
rect 513408 370170 513478 370226
rect 513534 370170 513602 370226
rect 513658 370170 513728 370226
rect 513408 370102 513728 370170
rect 513408 370046 513478 370102
rect 513534 370046 513602 370102
rect 513658 370046 513728 370102
rect 513408 369978 513728 370046
rect 513408 369922 513478 369978
rect 513534 369922 513602 369978
rect 513658 369922 513728 369978
rect 513408 369888 513728 369922
rect 544128 370350 544448 370384
rect 544128 370294 544198 370350
rect 544254 370294 544322 370350
rect 544378 370294 544448 370350
rect 544128 370226 544448 370294
rect 544128 370170 544198 370226
rect 544254 370170 544322 370226
rect 544378 370170 544448 370226
rect 544128 370102 544448 370170
rect 544128 370046 544198 370102
rect 544254 370046 544322 370102
rect 544378 370046 544448 370102
rect 544128 369978 544448 370046
rect 544128 369922 544198 369978
rect 544254 369922 544322 369978
rect 544378 369922 544448 369978
rect 544128 369888 544448 369922
rect 574848 370350 575168 370384
rect 574848 370294 574918 370350
rect 574974 370294 575042 370350
rect 575098 370294 575168 370350
rect 574848 370226 575168 370294
rect 574848 370170 574918 370226
rect 574974 370170 575042 370226
rect 575098 370170 575168 370226
rect 574848 370102 575168 370170
rect 574848 370046 574918 370102
rect 574974 370046 575042 370102
rect 575098 370046 575168 370102
rect 574848 369978 575168 370046
rect 574848 369922 574918 369978
rect 574974 369922 575042 369978
rect 575098 369922 575168 369978
rect 574848 369888 575168 369922
rect 340620 365988 340676 365998
rect 340620 361228 340676 365932
rect 344448 364350 344768 364384
rect 344448 364294 344518 364350
rect 344574 364294 344642 364350
rect 344698 364294 344768 364350
rect 344448 364226 344768 364294
rect 344448 364170 344518 364226
rect 344574 364170 344642 364226
rect 344698 364170 344768 364226
rect 344448 364102 344768 364170
rect 344448 364046 344518 364102
rect 344574 364046 344642 364102
rect 344698 364046 344768 364102
rect 344448 363978 344768 364046
rect 344448 363922 344518 363978
rect 344574 363922 344642 363978
rect 344698 363922 344768 363978
rect 344448 363888 344768 363922
rect 375168 364350 375488 364384
rect 375168 364294 375238 364350
rect 375294 364294 375362 364350
rect 375418 364294 375488 364350
rect 375168 364226 375488 364294
rect 375168 364170 375238 364226
rect 375294 364170 375362 364226
rect 375418 364170 375488 364226
rect 375168 364102 375488 364170
rect 375168 364046 375238 364102
rect 375294 364046 375362 364102
rect 375418 364046 375488 364102
rect 375168 363978 375488 364046
rect 375168 363922 375238 363978
rect 375294 363922 375362 363978
rect 375418 363922 375488 363978
rect 375168 363888 375488 363922
rect 405888 364350 406208 364384
rect 405888 364294 405958 364350
rect 406014 364294 406082 364350
rect 406138 364294 406208 364350
rect 405888 364226 406208 364294
rect 405888 364170 405958 364226
rect 406014 364170 406082 364226
rect 406138 364170 406208 364226
rect 405888 364102 406208 364170
rect 405888 364046 405958 364102
rect 406014 364046 406082 364102
rect 406138 364046 406208 364102
rect 405888 363978 406208 364046
rect 405888 363922 405958 363978
rect 406014 363922 406082 363978
rect 406138 363922 406208 363978
rect 405888 363888 406208 363922
rect 436608 364350 436928 364384
rect 436608 364294 436678 364350
rect 436734 364294 436802 364350
rect 436858 364294 436928 364350
rect 436608 364226 436928 364294
rect 436608 364170 436678 364226
rect 436734 364170 436802 364226
rect 436858 364170 436928 364226
rect 436608 364102 436928 364170
rect 436608 364046 436678 364102
rect 436734 364046 436802 364102
rect 436858 364046 436928 364102
rect 436608 363978 436928 364046
rect 436608 363922 436678 363978
rect 436734 363922 436802 363978
rect 436858 363922 436928 363978
rect 436608 363888 436928 363922
rect 467328 364350 467648 364384
rect 467328 364294 467398 364350
rect 467454 364294 467522 364350
rect 467578 364294 467648 364350
rect 467328 364226 467648 364294
rect 467328 364170 467398 364226
rect 467454 364170 467522 364226
rect 467578 364170 467648 364226
rect 467328 364102 467648 364170
rect 467328 364046 467398 364102
rect 467454 364046 467522 364102
rect 467578 364046 467648 364102
rect 467328 363978 467648 364046
rect 467328 363922 467398 363978
rect 467454 363922 467522 363978
rect 467578 363922 467648 363978
rect 467328 363888 467648 363922
rect 498048 364350 498368 364384
rect 498048 364294 498118 364350
rect 498174 364294 498242 364350
rect 498298 364294 498368 364350
rect 498048 364226 498368 364294
rect 498048 364170 498118 364226
rect 498174 364170 498242 364226
rect 498298 364170 498368 364226
rect 498048 364102 498368 364170
rect 498048 364046 498118 364102
rect 498174 364046 498242 364102
rect 498298 364046 498368 364102
rect 498048 363978 498368 364046
rect 498048 363922 498118 363978
rect 498174 363922 498242 363978
rect 498298 363922 498368 363978
rect 498048 363888 498368 363922
rect 528768 364350 529088 364384
rect 528768 364294 528838 364350
rect 528894 364294 528962 364350
rect 529018 364294 529088 364350
rect 528768 364226 529088 364294
rect 528768 364170 528838 364226
rect 528894 364170 528962 364226
rect 529018 364170 529088 364226
rect 528768 364102 529088 364170
rect 528768 364046 528838 364102
rect 528894 364046 528962 364102
rect 529018 364046 529088 364102
rect 528768 363978 529088 364046
rect 528768 363922 528838 363978
rect 528894 363922 528962 363978
rect 529018 363922 529088 363978
rect 528768 363888 529088 363922
rect 559488 364350 559808 364384
rect 559488 364294 559558 364350
rect 559614 364294 559682 364350
rect 559738 364294 559808 364350
rect 559488 364226 559808 364294
rect 559488 364170 559558 364226
rect 559614 364170 559682 364226
rect 559738 364170 559808 364226
rect 559488 364102 559808 364170
rect 559488 364046 559558 364102
rect 559614 364046 559682 364102
rect 559738 364046 559808 364102
rect 559488 363978 559808 364046
rect 559488 363922 559558 363978
rect 559614 363922 559682 363978
rect 559738 363922 559808 363978
rect 559488 363888 559808 363922
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 340620 361172 340900 361228
rect 340508 157552 340564 157562
rect 340620 335524 340676 335534
rect 340620 142660 340676 335468
rect 340844 157438 340900 361172
rect 359808 352350 360128 352384
rect 359808 352294 359878 352350
rect 359934 352294 360002 352350
rect 360058 352294 360128 352350
rect 359808 352226 360128 352294
rect 359808 352170 359878 352226
rect 359934 352170 360002 352226
rect 360058 352170 360128 352226
rect 359808 352102 360128 352170
rect 359808 352046 359878 352102
rect 359934 352046 360002 352102
rect 360058 352046 360128 352102
rect 359808 351978 360128 352046
rect 359808 351922 359878 351978
rect 359934 351922 360002 351978
rect 360058 351922 360128 351978
rect 359808 351888 360128 351922
rect 390528 352350 390848 352384
rect 390528 352294 390598 352350
rect 390654 352294 390722 352350
rect 390778 352294 390848 352350
rect 390528 352226 390848 352294
rect 390528 352170 390598 352226
rect 390654 352170 390722 352226
rect 390778 352170 390848 352226
rect 390528 352102 390848 352170
rect 390528 352046 390598 352102
rect 390654 352046 390722 352102
rect 390778 352046 390848 352102
rect 390528 351978 390848 352046
rect 390528 351922 390598 351978
rect 390654 351922 390722 351978
rect 390778 351922 390848 351978
rect 390528 351888 390848 351922
rect 421248 352350 421568 352384
rect 421248 352294 421318 352350
rect 421374 352294 421442 352350
rect 421498 352294 421568 352350
rect 421248 352226 421568 352294
rect 421248 352170 421318 352226
rect 421374 352170 421442 352226
rect 421498 352170 421568 352226
rect 421248 352102 421568 352170
rect 421248 352046 421318 352102
rect 421374 352046 421442 352102
rect 421498 352046 421568 352102
rect 421248 351978 421568 352046
rect 421248 351922 421318 351978
rect 421374 351922 421442 351978
rect 421498 351922 421568 351978
rect 421248 351888 421568 351922
rect 451968 352350 452288 352384
rect 451968 352294 452038 352350
rect 452094 352294 452162 352350
rect 452218 352294 452288 352350
rect 451968 352226 452288 352294
rect 451968 352170 452038 352226
rect 452094 352170 452162 352226
rect 452218 352170 452288 352226
rect 451968 352102 452288 352170
rect 451968 352046 452038 352102
rect 452094 352046 452162 352102
rect 452218 352046 452288 352102
rect 451968 351978 452288 352046
rect 451968 351922 452038 351978
rect 452094 351922 452162 351978
rect 452218 351922 452288 351978
rect 451968 351888 452288 351922
rect 482688 352350 483008 352384
rect 482688 352294 482758 352350
rect 482814 352294 482882 352350
rect 482938 352294 483008 352350
rect 482688 352226 483008 352294
rect 482688 352170 482758 352226
rect 482814 352170 482882 352226
rect 482938 352170 483008 352226
rect 482688 352102 483008 352170
rect 482688 352046 482758 352102
rect 482814 352046 482882 352102
rect 482938 352046 483008 352102
rect 482688 351978 483008 352046
rect 482688 351922 482758 351978
rect 482814 351922 482882 351978
rect 482938 351922 483008 351978
rect 482688 351888 483008 351922
rect 513408 352350 513728 352384
rect 513408 352294 513478 352350
rect 513534 352294 513602 352350
rect 513658 352294 513728 352350
rect 513408 352226 513728 352294
rect 513408 352170 513478 352226
rect 513534 352170 513602 352226
rect 513658 352170 513728 352226
rect 513408 352102 513728 352170
rect 513408 352046 513478 352102
rect 513534 352046 513602 352102
rect 513658 352046 513728 352102
rect 513408 351978 513728 352046
rect 513408 351922 513478 351978
rect 513534 351922 513602 351978
rect 513658 351922 513728 351978
rect 513408 351888 513728 351922
rect 544128 352350 544448 352384
rect 544128 352294 544198 352350
rect 544254 352294 544322 352350
rect 544378 352294 544448 352350
rect 544128 352226 544448 352294
rect 544128 352170 544198 352226
rect 544254 352170 544322 352226
rect 544378 352170 544448 352226
rect 544128 352102 544448 352170
rect 544128 352046 544198 352102
rect 544254 352046 544322 352102
rect 544378 352046 544448 352102
rect 544128 351978 544448 352046
rect 544128 351922 544198 351978
rect 544254 351922 544322 351978
rect 544378 351922 544448 351978
rect 544128 351888 544448 351922
rect 574848 352350 575168 352384
rect 574848 352294 574918 352350
rect 574974 352294 575042 352350
rect 575098 352294 575168 352350
rect 574848 352226 575168 352294
rect 574848 352170 574918 352226
rect 574974 352170 575042 352226
rect 575098 352170 575168 352226
rect 574848 352102 575168 352170
rect 574848 352046 574918 352102
rect 574974 352046 575042 352102
rect 575098 352046 575168 352102
rect 574848 351978 575168 352046
rect 574848 351922 574918 351978
rect 574974 351922 575042 351978
rect 575098 351922 575168 351978
rect 574848 351888 575168 351922
rect 344448 346350 344768 346384
rect 344448 346294 344518 346350
rect 344574 346294 344642 346350
rect 344698 346294 344768 346350
rect 344448 346226 344768 346294
rect 344448 346170 344518 346226
rect 344574 346170 344642 346226
rect 344698 346170 344768 346226
rect 344448 346102 344768 346170
rect 344448 346046 344518 346102
rect 344574 346046 344642 346102
rect 344698 346046 344768 346102
rect 344448 345978 344768 346046
rect 344448 345922 344518 345978
rect 344574 345922 344642 345978
rect 344698 345922 344768 345978
rect 344448 345888 344768 345922
rect 375168 346350 375488 346384
rect 375168 346294 375238 346350
rect 375294 346294 375362 346350
rect 375418 346294 375488 346350
rect 375168 346226 375488 346294
rect 375168 346170 375238 346226
rect 375294 346170 375362 346226
rect 375418 346170 375488 346226
rect 375168 346102 375488 346170
rect 375168 346046 375238 346102
rect 375294 346046 375362 346102
rect 375418 346046 375488 346102
rect 375168 345978 375488 346046
rect 375168 345922 375238 345978
rect 375294 345922 375362 345978
rect 375418 345922 375488 345978
rect 375168 345888 375488 345922
rect 405888 346350 406208 346384
rect 405888 346294 405958 346350
rect 406014 346294 406082 346350
rect 406138 346294 406208 346350
rect 405888 346226 406208 346294
rect 405888 346170 405958 346226
rect 406014 346170 406082 346226
rect 406138 346170 406208 346226
rect 405888 346102 406208 346170
rect 405888 346046 405958 346102
rect 406014 346046 406082 346102
rect 406138 346046 406208 346102
rect 405888 345978 406208 346046
rect 405888 345922 405958 345978
rect 406014 345922 406082 345978
rect 406138 345922 406208 345978
rect 405888 345888 406208 345922
rect 436608 346350 436928 346384
rect 436608 346294 436678 346350
rect 436734 346294 436802 346350
rect 436858 346294 436928 346350
rect 436608 346226 436928 346294
rect 436608 346170 436678 346226
rect 436734 346170 436802 346226
rect 436858 346170 436928 346226
rect 436608 346102 436928 346170
rect 436608 346046 436678 346102
rect 436734 346046 436802 346102
rect 436858 346046 436928 346102
rect 436608 345978 436928 346046
rect 436608 345922 436678 345978
rect 436734 345922 436802 345978
rect 436858 345922 436928 345978
rect 436608 345888 436928 345922
rect 467328 346350 467648 346384
rect 467328 346294 467398 346350
rect 467454 346294 467522 346350
rect 467578 346294 467648 346350
rect 467328 346226 467648 346294
rect 467328 346170 467398 346226
rect 467454 346170 467522 346226
rect 467578 346170 467648 346226
rect 467328 346102 467648 346170
rect 467328 346046 467398 346102
rect 467454 346046 467522 346102
rect 467578 346046 467648 346102
rect 467328 345978 467648 346046
rect 467328 345922 467398 345978
rect 467454 345922 467522 345978
rect 467578 345922 467648 345978
rect 467328 345888 467648 345922
rect 498048 346350 498368 346384
rect 498048 346294 498118 346350
rect 498174 346294 498242 346350
rect 498298 346294 498368 346350
rect 498048 346226 498368 346294
rect 498048 346170 498118 346226
rect 498174 346170 498242 346226
rect 498298 346170 498368 346226
rect 498048 346102 498368 346170
rect 498048 346046 498118 346102
rect 498174 346046 498242 346102
rect 498298 346046 498368 346102
rect 498048 345978 498368 346046
rect 498048 345922 498118 345978
rect 498174 345922 498242 345978
rect 498298 345922 498368 345978
rect 498048 345888 498368 345922
rect 528768 346350 529088 346384
rect 528768 346294 528838 346350
rect 528894 346294 528962 346350
rect 529018 346294 529088 346350
rect 528768 346226 529088 346294
rect 528768 346170 528838 346226
rect 528894 346170 528962 346226
rect 529018 346170 529088 346226
rect 528768 346102 529088 346170
rect 528768 346046 528838 346102
rect 528894 346046 528962 346102
rect 529018 346046 529088 346102
rect 528768 345978 529088 346046
rect 528768 345922 528838 345978
rect 528894 345922 528962 345978
rect 529018 345922 529088 345978
rect 528768 345888 529088 345922
rect 559488 346350 559808 346384
rect 559488 346294 559558 346350
rect 559614 346294 559682 346350
rect 559738 346294 559808 346350
rect 559488 346226 559808 346294
rect 559488 346170 559558 346226
rect 559614 346170 559682 346226
rect 559738 346170 559808 346226
rect 559488 346102 559808 346170
rect 559488 346046 559558 346102
rect 559614 346046 559682 346102
rect 559738 346046 559808 346102
rect 559488 345978 559808 346046
rect 559488 345922 559558 345978
rect 559614 345922 559682 345978
rect 559738 345922 559808 345978
rect 559488 345888 559808 345922
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 359808 334350 360128 334384
rect 359808 334294 359878 334350
rect 359934 334294 360002 334350
rect 360058 334294 360128 334350
rect 359808 334226 360128 334294
rect 359808 334170 359878 334226
rect 359934 334170 360002 334226
rect 360058 334170 360128 334226
rect 359808 334102 360128 334170
rect 359808 334046 359878 334102
rect 359934 334046 360002 334102
rect 360058 334046 360128 334102
rect 359808 333978 360128 334046
rect 359808 333922 359878 333978
rect 359934 333922 360002 333978
rect 360058 333922 360128 333978
rect 359808 333888 360128 333922
rect 390528 334350 390848 334384
rect 390528 334294 390598 334350
rect 390654 334294 390722 334350
rect 390778 334294 390848 334350
rect 390528 334226 390848 334294
rect 390528 334170 390598 334226
rect 390654 334170 390722 334226
rect 390778 334170 390848 334226
rect 390528 334102 390848 334170
rect 390528 334046 390598 334102
rect 390654 334046 390722 334102
rect 390778 334046 390848 334102
rect 390528 333978 390848 334046
rect 390528 333922 390598 333978
rect 390654 333922 390722 333978
rect 390778 333922 390848 333978
rect 390528 333888 390848 333922
rect 421248 334350 421568 334384
rect 421248 334294 421318 334350
rect 421374 334294 421442 334350
rect 421498 334294 421568 334350
rect 421248 334226 421568 334294
rect 421248 334170 421318 334226
rect 421374 334170 421442 334226
rect 421498 334170 421568 334226
rect 421248 334102 421568 334170
rect 421248 334046 421318 334102
rect 421374 334046 421442 334102
rect 421498 334046 421568 334102
rect 421248 333978 421568 334046
rect 421248 333922 421318 333978
rect 421374 333922 421442 333978
rect 421498 333922 421568 333978
rect 421248 333888 421568 333922
rect 451968 334350 452288 334384
rect 451968 334294 452038 334350
rect 452094 334294 452162 334350
rect 452218 334294 452288 334350
rect 451968 334226 452288 334294
rect 451968 334170 452038 334226
rect 452094 334170 452162 334226
rect 452218 334170 452288 334226
rect 451968 334102 452288 334170
rect 451968 334046 452038 334102
rect 452094 334046 452162 334102
rect 452218 334046 452288 334102
rect 451968 333978 452288 334046
rect 451968 333922 452038 333978
rect 452094 333922 452162 333978
rect 452218 333922 452288 333978
rect 451968 333888 452288 333922
rect 482688 334350 483008 334384
rect 482688 334294 482758 334350
rect 482814 334294 482882 334350
rect 482938 334294 483008 334350
rect 482688 334226 483008 334294
rect 482688 334170 482758 334226
rect 482814 334170 482882 334226
rect 482938 334170 483008 334226
rect 482688 334102 483008 334170
rect 482688 334046 482758 334102
rect 482814 334046 482882 334102
rect 482938 334046 483008 334102
rect 482688 333978 483008 334046
rect 482688 333922 482758 333978
rect 482814 333922 482882 333978
rect 482938 333922 483008 333978
rect 482688 333888 483008 333922
rect 513408 334350 513728 334384
rect 513408 334294 513478 334350
rect 513534 334294 513602 334350
rect 513658 334294 513728 334350
rect 513408 334226 513728 334294
rect 513408 334170 513478 334226
rect 513534 334170 513602 334226
rect 513658 334170 513728 334226
rect 513408 334102 513728 334170
rect 513408 334046 513478 334102
rect 513534 334046 513602 334102
rect 513658 334046 513728 334102
rect 513408 333978 513728 334046
rect 513408 333922 513478 333978
rect 513534 333922 513602 333978
rect 513658 333922 513728 333978
rect 513408 333888 513728 333922
rect 544128 334350 544448 334384
rect 544128 334294 544198 334350
rect 544254 334294 544322 334350
rect 544378 334294 544448 334350
rect 544128 334226 544448 334294
rect 544128 334170 544198 334226
rect 544254 334170 544322 334226
rect 544378 334170 544448 334226
rect 544128 334102 544448 334170
rect 544128 334046 544198 334102
rect 544254 334046 544322 334102
rect 544378 334046 544448 334102
rect 544128 333978 544448 334046
rect 544128 333922 544198 333978
rect 544254 333922 544322 333978
rect 544378 333922 544448 333978
rect 544128 333888 544448 333922
rect 574848 334350 575168 334384
rect 574848 334294 574918 334350
rect 574974 334294 575042 334350
rect 575098 334294 575168 334350
rect 574848 334226 575168 334294
rect 574848 334170 574918 334226
rect 574974 334170 575042 334226
rect 575098 334170 575168 334226
rect 574848 334102 575168 334170
rect 574848 334046 574918 334102
rect 574974 334046 575042 334102
rect 575098 334046 575168 334102
rect 574848 333978 575168 334046
rect 574848 333922 574918 333978
rect 574974 333922 575042 333978
rect 575098 333922 575168 333978
rect 574848 333888 575168 333922
rect 344448 328350 344768 328384
rect 344448 328294 344518 328350
rect 344574 328294 344642 328350
rect 344698 328294 344768 328350
rect 344448 328226 344768 328294
rect 344448 328170 344518 328226
rect 344574 328170 344642 328226
rect 344698 328170 344768 328226
rect 344448 328102 344768 328170
rect 344448 328046 344518 328102
rect 344574 328046 344642 328102
rect 344698 328046 344768 328102
rect 344448 327978 344768 328046
rect 344448 327922 344518 327978
rect 344574 327922 344642 327978
rect 344698 327922 344768 327978
rect 344448 327888 344768 327922
rect 375168 328350 375488 328384
rect 375168 328294 375238 328350
rect 375294 328294 375362 328350
rect 375418 328294 375488 328350
rect 375168 328226 375488 328294
rect 375168 328170 375238 328226
rect 375294 328170 375362 328226
rect 375418 328170 375488 328226
rect 375168 328102 375488 328170
rect 375168 328046 375238 328102
rect 375294 328046 375362 328102
rect 375418 328046 375488 328102
rect 375168 327978 375488 328046
rect 375168 327922 375238 327978
rect 375294 327922 375362 327978
rect 375418 327922 375488 327978
rect 375168 327888 375488 327922
rect 405888 328350 406208 328384
rect 405888 328294 405958 328350
rect 406014 328294 406082 328350
rect 406138 328294 406208 328350
rect 405888 328226 406208 328294
rect 405888 328170 405958 328226
rect 406014 328170 406082 328226
rect 406138 328170 406208 328226
rect 405888 328102 406208 328170
rect 405888 328046 405958 328102
rect 406014 328046 406082 328102
rect 406138 328046 406208 328102
rect 405888 327978 406208 328046
rect 405888 327922 405958 327978
rect 406014 327922 406082 327978
rect 406138 327922 406208 327978
rect 405888 327888 406208 327922
rect 436608 328350 436928 328384
rect 436608 328294 436678 328350
rect 436734 328294 436802 328350
rect 436858 328294 436928 328350
rect 436608 328226 436928 328294
rect 436608 328170 436678 328226
rect 436734 328170 436802 328226
rect 436858 328170 436928 328226
rect 436608 328102 436928 328170
rect 436608 328046 436678 328102
rect 436734 328046 436802 328102
rect 436858 328046 436928 328102
rect 436608 327978 436928 328046
rect 436608 327922 436678 327978
rect 436734 327922 436802 327978
rect 436858 327922 436928 327978
rect 436608 327888 436928 327922
rect 467328 328350 467648 328384
rect 467328 328294 467398 328350
rect 467454 328294 467522 328350
rect 467578 328294 467648 328350
rect 467328 328226 467648 328294
rect 467328 328170 467398 328226
rect 467454 328170 467522 328226
rect 467578 328170 467648 328226
rect 467328 328102 467648 328170
rect 467328 328046 467398 328102
rect 467454 328046 467522 328102
rect 467578 328046 467648 328102
rect 467328 327978 467648 328046
rect 467328 327922 467398 327978
rect 467454 327922 467522 327978
rect 467578 327922 467648 327978
rect 467328 327888 467648 327922
rect 498048 328350 498368 328384
rect 498048 328294 498118 328350
rect 498174 328294 498242 328350
rect 498298 328294 498368 328350
rect 498048 328226 498368 328294
rect 498048 328170 498118 328226
rect 498174 328170 498242 328226
rect 498298 328170 498368 328226
rect 498048 328102 498368 328170
rect 498048 328046 498118 328102
rect 498174 328046 498242 328102
rect 498298 328046 498368 328102
rect 498048 327978 498368 328046
rect 498048 327922 498118 327978
rect 498174 327922 498242 327978
rect 498298 327922 498368 327978
rect 498048 327888 498368 327922
rect 528768 328350 529088 328384
rect 528768 328294 528838 328350
rect 528894 328294 528962 328350
rect 529018 328294 529088 328350
rect 528768 328226 529088 328294
rect 528768 328170 528838 328226
rect 528894 328170 528962 328226
rect 529018 328170 529088 328226
rect 528768 328102 529088 328170
rect 528768 328046 528838 328102
rect 528894 328046 528962 328102
rect 529018 328046 529088 328102
rect 528768 327978 529088 328046
rect 528768 327922 528838 327978
rect 528894 327922 528962 327978
rect 529018 327922 529088 327978
rect 528768 327888 529088 327922
rect 559488 328350 559808 328384
rect 559488 328294 559558 328350
rect 559614 328294 559682 328350
rect 559738 328294 559808 328350
rect 559488 328226 559808 328294
rect 559488 328170 559558 328226
rect 559614 328170 559682 328226
rect 559738 328170 559808 328226
rect 559488 328102 559808 328170
rect 559488 328046 559558 328102
rect 559614 328046 559682 328102
rect 559738 328046 559808 328102
rect 559488 327978 559808 328046
rect 559488 327922 559558 327978
rect 559614 327922 559682 327978
rect 559738 327922 559808 327978
rect 559488 327888 559808 327922
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 359808 316350 360128 316384
rect 359808 316294 359878 316350
rect 359934 316294 360002 316350
rect 360058 316294 360128 316350
rect 359808 316226 360128 316294
rect 359808 316170 359878 316226
rect 359934 316170 360002 316226
rect 360058 316170 360128 316226
rect 359808 316102 360128 316170
rect 359808 316046 359878 316102
rect 359934 316046 360002 316102
rect 360058 316046 360128 316102
rect 359808 315978 360128 316046
rect 359808 315922 359878 315978
rect 359934 315922 360002 315978
rect 360058 315922 360128 315978
rect 359808 315888 360128 315922
rect 390528 316350 390848 316384
rect 390528 316294 390598 316350
rect 390654 316294 390722 316350
rect 390778 316294 390848 316350
rect 390528 316226 390848 316294
rect 390528 316170 390598 316226
rect 390654 316170 390722 316226
rect 390778 316170 390848 316226
rect 390528 316102 390848 316170
rect 390528 316046 390598 316102
rect 390654 316046 390722 316102
rect 390778 316046 390848 316102
rect 390528 315978 390848 316046
rect 390528 315922 390598 315978
rect 390654 315922 390722 315978
rect 390778 315922 390848 315978
rect 390528 315888 390848 315922
rect 421248 316350 421568 316384
rect 421248 316294 421318 316350
rect 421374 316294 421442 316350
rect 421498 316294 421568 316350
rect 421248 316226 421568 316294
rect 421248 316170 421318 316226
rect 421374 316170 421442 316226
rect 421498 316170 421568 316226
rect 421248 316102 421568 316170
rect 421248 316046 421318 316102
rect 421374 316046 421442 316102
rect 421498 316046 421568 316102
rect 421248 315978 421568 316046
rect 421248 315922 421318 315978
rect 421374 315922 421442 315978
rect 421498 315922 421568 315978
rect 421248 315888 421568 315922
rect 451968 316350 452288 316384
rect 451968 316294 452038 316350
rect 452094 316294 452162 316350
rect 452218 316294 452288 316350
rect 451968 316226 452288 316294
rect 451968 316170 452038 316226
rect 452094 316170 452162 316226
rect 452218 316170 452288 316226
rect 451968 316102 452288 316170
rect 451968 316046 452038 316102
rect 452094 316046 452162 316102
rect 452218 316046 452288 316102
rect 451968 315978 452288 316046
rect 451968 315922 452038 315978
rect 452094 315922 452162 315978
rect 452218 315922 452288 315978
rect 451968 315888 452288 315922
rect 482688 316350 483008 316384
rect 482688 316294 482758 316350
rect 482814 316294 482882 316350
rect 482938 316294 483008 316350
rect 482688 316226 483008 316294
rect 482688 316170 482758 316226
rect 482814 316170 482882 316226
rect 482938 316170 483008 316226
rect 482688 316102 483008 316170
rect 482688 316046 482758 316102
rect 482814 316046 482882 316102
rect 482938 316046 483008 316102
rect 482688 315978 483008 316046
rect 482688 315922 482758 315978
rect 482814 315922 482882 315978
rect 482938 315922 483008 315978
rect 482688 315888 483008 315922
rect 513408 316350 513728 316384
rect 513408 316294 513478 316350
rect 513534 316294 513602 316350
rect 513658 316294 513728 316350
rect 513408 316226 513728 316294
rect 513408 316170 513478 316226
rect 513534 316170 513602 316226
rect 513658 316170 513728 316226
rect 513408 316102 513728 316170
rect 513408 316046 513478 316102
rect 513534 316046 513602 316102
rect 513658 316046 513728 316102
rect 513408 315978 513728 316046
rect 513408 315922 513478 315978
rect 513534 315922 513602 315978
rect 513658 315922 513728 315978
rect 513408 315888 513728 315922
rect 544128 316350 544448 316384
rect 544128 316294 544198 316350
rect 544254 316294 544322 316350
rect 544378 316294 544448 316350
rect 544128 316226 544448 316294
rect 544128 316170 544198 316226
rect 544254 316170 544322 316226
rect 544378 316170 544448 316226
rect 544128 316102 544448 316170
rect 544128 316046 544198 316102
rect 544254 316046 544322 316102
rect 544378 316046 544448 316102
rect 544128 315978 544448 316046
rect 544128 315922 544198 315978
rect 544254 315922 544322 315978
rect 544378 315922 544448 315978
rect 544128 315888 544448 315922
rect 574848 316350 575168 316384
rect 574848 316294 574918 316350
rect 574974 316294 575042 316350
rect 575098 316294 575168 316350
rect 574848 316226 575168 316294
rect 574848 316170 574918 316226
rect 574974 316170 575042 316226
rect 575098 316170 575168 316226
rect 574848 316102 575168 316170
rect 574848 316046 574918 316102
rect 574974 316046 575042 316102
rect 575098 316046 575168 316102
rect 574848 315978 575168 316046
rect 574848 315922 574918 315978
rect 574974 315922 575042 315978
rect 575098 315922 575168 315978
rect 574848 315888 575168 315922
rect 344448 310350 344768 310384
rect 344448 310294 344518 310350
rect 344574 310294 344642 310350
rect 344698 310294 344768 310350
rect 344448 310226 344768 310294
rect 344448 310170 344518 310226
rect 344574 310170 344642 310226
rect 344698 310170 344768 310226
rect 344448 310102 344768 310170
rect 344448 310046 344518 310102
rect 344574 310046 344642 310102
rect 344698 310046 344768 310102
rect 344448 309978 344768 310046
rect 344448 309922 344518 309978
rect 344574 309922 344642 309978
rect 344698 309922 344768 309978
rect 344448 309888 344768 309922
rect 375168 310350 375488 310384
rect 375168 310294 375238 310350
rect 375294 310294 375362 310350
rect 375418 310294 375488 310350
rect 375168 310226 375488 310294
rect 375168 310170 375238 310226
rect 375294 310170 375362 310226
rect 375418 310170 375488 310226
rect 375168 310102 375488 310170
rect 375168 310046 375238 310102
rect 375294 310046 375362 310102
rect 375418 310046 375488 310102
rect 375168 309978 375488 310046
rect 375168 309922 375238 309978
rect 375294 309922 375362 309978
rect 375418 309922 375488 309978
rect 375168 309888 375488 309922
rect 405888 310350 406208 310384
rect 405888 310294 405958 310350
rect 406014 310294 406082 310350
rect 406138 310294 406208 310350
rect 405888 310226 406208 310294
rect 405888 310170 405958 310226
rect 406014 310170 406082 310226
rect 406138 310170 406208 310226
rect 405888 310102 406208 310170
rect 405888 310046 405958 310102
rect 406014 310046 406082 310102
rect 406138 310046 406208 310102
rect 405888 309978 406208 310046
rect 405888 309922 405958 309978
rect 406014 309922 406082 309978
rect 406138 309922 406208 309978
rect 405888 309888 406208 309922
rect 436608 310350 436928 310384
rect 436608 310294 436678 310350
rect 436734 310294 436802 310350
rect 436858 310294 436928 310350
rect 436608 310226 436928 310294
rect 436608 310170 436678 310226
rect 436734 310170 436802 310226
rect 436858 310170 436928 310226
rect 436608 310102 436928 310170
rect 436608 310046 436678 310102
rect 436734 310046 436802 310102
rect 436858 310046 436928 310102
rect 436608 309978 436928 310046
rect 436608 309922 436678 309978
rect 436734 309922 436802 309978
rect 436858 309922 436928 309978
rect 436608 309888 436928 309922
rect 467328 310350 467648 310384
rect 467328 310294 467398 310350
rect 467454 310294 467522 310350
rect 467578 310294 467648 310350
rect 467328 310226 467648 310294
rect 467328 310170 467398 310226
rect 467454 310170 467522 310226
rect 467578 310170 467648 310226
rect 467328 310102 467648 310170
rect 467328 310046 467398 310102
rect 467454 310046 467522 310102
rect 467578 310046 467648 310102
rect 467328 309978 467648 310046
rect 467328 309922 467398 309978
rect 467454 309922 467522 309978
rect 467578 309922 467648 309978
rect 467328 309888 467648 309922
rect 498048 310350 498368 310384
rect 498048 310294 498118 310350
rect 498174 310294 498242 310350
rect 498298 310294 498368 310350
rect 498048 310226 498368 310294
rect 498048 310170 498118 310226
rect 498174 310170 498242 310226
rect 498298 310170 498368 310226
rect 498048 310102 498368 310170
rect 498048 310046 498118 310102
rect 498174 310046 498242 310102
rect 498298 310046 498368 310102
rect 498048 309978 498368 310046
rect 498048 309922 498118 309978
rect 498174 309922 498242 309978
rect 498298 309922 498368 309978
rect 498048 309888 498368 309922
rect 528768 310350 529088 310384
rect 528768 310294 528838 310350
rect 528894 310294 528962 310350
rect 529018 310294 529088 310350
rect 528768 310226 529088 310294
rect 528768 310170 528838 310226
rect 528894 310170 528962 310226
rect 529018 310170 529088 310226
rect 528768 310102 529088 310170
rect 528768 310046 528838 310102
rect 528894 310046 528962 310102
rect 529018 310046 529088 310102
rect 528768 309978 529088 310046
rect 528768 309922 528838 309978
rect 528894 309922 528962 309978
rect 529018 309922 529088 309978
rect 528768 309888 529088 309922
rect 559488 310350 559808 310384
rect 559488 310294 559558 310350
rect 559614 310294 559682 310350
rect 559738 310294 559808 310350
rect 559488 310226 559808 310294
rect 559488 310170 559558 310226
rect 559614 310170 559682 310226
rect 559738 310170 559808 310226
rect 559488 310102 559808 310170
rect 559488 310046 559558 310102
rect 559614 310046 559682 310102
rect 559738 310046 559808 310102
rect 559488 309978 559808 310046
rect 559488 309922 559558 309978
rect 559614 309922 559682 309978
rect 559738 309922 559808 309978
rect 559488 309888 559808 309922
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 341068 301618 341124 301628
rect 340844 157372 340900 157382
rect 340956 294598 341012 294608
rect 340620 142594 340676 142604
rect 340956 138538 341012 294542
rect 341068 283798 341124 301562
rect 359808 298350 360128 298384
rect 359808 298294 359878 298350
rect 359934 298294 360002 298350
rect 360058 298294 360128 298350
rect 359808 298226 360128 298294
rect 359808 298170 359878 298226
rect 359934 298170 360002 298226
rect 360058 298170 360128 298226
rect 359808 298102 360128 298170
rect 359808 298046 359878 298102
rect 359934 298046 360002 298102
rect 360058 298046 360128 298102
rect 359808 297978 360128 298046
rect 359808 297922 359878 297978
rect 359934 297922 360002 297978
rect 360058 297922 360128 297978
rect 359808 297888 360128 297922
rect 390528 298350 390848 298384
rect 390528 298294 390598 298350
rect 390654 298294 390722 298350
rect 390778 298294 390848 298350
rect 390528 298226 390848 298294
rect 390528 298170 390598 298226
rect 390654 298170 390722 298226
rect 390778 298170 390848 298226
rect 390528 298102 390848 298170
rect 390528 298046 390598 298102
rect 390654 298046 390722 298102
rect 390778 298046 390848 298102
rect 390528 297978 390848 298046
rect 390528 297922 390598 297978
rect 390654 297922 390722 297978
rect 390778 297922 390848 297978
rect 390528 297888 390848 297922
rect 421248 298350 421568 298384
rect 421248 298294 421318 298350
rect 421374 298294 421442 298350
rect 421498 298294 421568 298350
rect 421248 298226 421568 298294
rect 421248 298170 421318 298226
rect 421374 298170 421442 298226
rect 421498 298170 421568 298226
rect 421248 298102 421568 298170
rect 421248 298046 421318 298102
rect 421374 298046 421442 298102
rect 421498 298046 421568 298102
rect 421248 297978 421568 298046
rect 421248 297922 421318 297978
rect 421374 297922 421442 297978
rect 421498 297922 421568 297978
rect 421248 297888 421568 297922
rect 451968 298350 452288 298384
rect 451968 298294 452038 298350
rect 452094 298294 452162 298350
rect 452218 298294 452288 298350
rect 451968 298226 452288 298294
rect 451968 298170 452038 298226
rect 452094 298170 452162 298226
rect 452218 298170 452288 298226
rect 451968 298102 452288 298170
rect 451968 298046 452038 298102
rect 452094 298046 452162 298102
rect 452218 298046 452288 298102
rect 451968 297978 452288 298046
rect 451968 297922 452038 297978
rect 452094 297922 452162 297978
rect 452218 297922 452288 297978
rect 451968 297888 452288 297922
rect 482688 298350 483008 298384
rect 482688 298294 482758 298350
rect 482814 298294 482882 298350
rect 482938 298294 483008 298350
rect 482688 298226 483008 298294
rect 482688 298170 482758 298226
rect 482814 298170 482882 298226
rect 482938 298170 483008 298226
rect 482688 298102 483008 298170
rect 482688 298046 482758 298102
rect 482814 298046 482882 298102
rect 482938 298046 483008 298102
rect 482688 297978 483008 298046
rect 482688 297922 482758 297978
rect 482814 297922 482882 297978
rect 482938 297922 483008 297978
rect 482688 297888 483008 297922
rect 513408 298350 513728 298384
rect 513408 298294 513478 298350
rect 513534 298294 513602 298350
rect 513658 298294 513728 298350
rect 513408 298226 513728 298294
rect 513408 298170 513478 298226
rect 513534 298170 513602 298226
rect 513658 298170 513728 298226
rect 513408 298102 513728 298170
rect 513408 298046 513478 298102
rect 513534 298046 513602 298102
rect 513658 298046 513728 298102
rect 513408 297978 513728 298046
rect 513408 297922 513478 297978
rect 513534 297922 513602 297978
rect 513658 297922 513728 297978
rect 513408 297888 513728 297922
rect 544128 298350 544448 298384
rect 544128 298294 544198 298350
rect 544254 298294 544322 298350
rect 544378 298294 544448 298350
rect 544128 298226 544448 298294
rect 544128 298170 544198 298226
rect 544254 298170 544322 298226
rect 544378 298170 544448 298226
rect 544128 298102 544448 298170
rect 544128 298046 544198 298102
rect 544254 298046 544322 298102
rect 544378 298046 544448 298102
rect 544128 297978 544448 298046
rect 544128 297922 544198 297978
rect 544254 297922 544322 297978
rect 544378 297922 544448 297978
rect 544128 297888 544448 297922
rect 574848 298350 575168 298384
rect 574848 298294 574918 298350
rect 574974 298294 575042 298350
rect 575098 298294 575168 298350
rect 574848 298226 575168 298294
rect 574848 298170 574918 298226
rect 574974 298170 575042 298226
rect 575098 298170 575168 298226
rect 574848 298102 575168 298170
rect 574848 298046 574918 298102
rect 574974 298046 575042 298102
rect 575098 298046 575168 298102
rect 574848 297978 575168 298046
rect 574848 297922 574918 297978
rect 574974 297922 575042 297978
rect 575098 297922 575168 297978
rect 574848 297888 575168 297922
rect 344448 292350 344768 292384
rect 344448 292294 344518 292350
rect 344574 292294 344642 292350
rect 344698 292294 344768 292350
rect 344448 292226 344768 292294
rect 344448 292170 344518 292226
rect 344574 292170 344642 292226
rect 344698 292170 344768 292226
rect 344448 292102 344768 292170
rect 344448 292046 344518 292102
rect 344574 292046 344642 292102
rect 344698 292046 344768 292102
rect 344448 291978 344768 292046
rect 344448 291922 344518 291978
rect 344574 291922 344642 291978
rect 344698 291922 344768 291978
rect 344448 291888 344768 291922
rect 375168 292350 375488 292384
rect 375168 292294 375238 292350
rect 375294 292294 375362 292350
rect 375418 292294 375488 292350
rect 375168 292226 375488 292294
rect 375168 292170 375238 292226
rect 375294 292170 375362 292226
rect 375418 292170 375488 292226
rect 375168 292102 375488 292170
rect 375168 292046 375238 292102
rect 375294 292046 375362 292102
rect 375418 292046 375488 292102
rect 375168 291978 375488 292046
rect 375168 291922 375238 291978
rect 375294 291922 375362 291978
rect 375418 291922 375488 291978
rect 375168 291888 375488 291922
rect 405888 292350 406208 292384
rect 405888 292294 405958 292350
rect 406014 292294 406082 292350
rect 406138 292294 406208 292350
rect 405888 292226 406208 292294
rect 405888 292170 405958 292226
rect 406014 292170 406082 292226
rect 406138 292170 406208 292226
rect 405888 292102 406208 292170
rect 405888 292046 405958 292102
rect 406014 292046 406082 292102
rect 406138 292046 406208 292102
rect 405888 291978 406208 292046
rect 405888 291922 405958 291978
rect 406014 291922 406082 291978
rect 406138 291922 406208 291978
rect 405888 291888 406208 291922
rect 436608 292350 436928 292384
rect 436608 292294 436678 292350
rect 436734 292294 436802 292350
rect 436858 292294 436928 292350
rect 436608 292226 436928 292294
rect 436608 292170 436678 292226
rect 436734 292170 436802 292226
rect 436858 292170 436928 292226
rect 436608 292102 436928 292170
rect 436608 292046 436678 292102
rect 436734 292046 436802 292102
rect 436858 292046 436928 292102
rect 436608 291978 436928 292046
rect 436608 291922 436678 291978
rect 436734 291922 436802 291978
rect 436858 291922 436928 291978
rect 436608 291888 436928 291922
rect 467328 292350 467648 292384
rect 467328 292294 467398 292350
rect 467454 292294 467522 292350
rect 467578 292294 467648 292350
rect 467328 292226 467648 292294
rect 467328 292170 467398 292226
rect 467454 292170 467522 292226
rect 467578 292170 467648 292226
rect 467328 292102 467648 292170
rect 467328 292046 467398 292102
rect 467454 292046 467522 292102
rect 467578 292046 467648 292102
rect 467328 291978 467648 292046
rect 467328 291922 467398 291978
rect 467454 291922 467522 291978
rect 467578 291922 467648 291978
rect 467328 291888 467648 291922
rect 498048 292350 498368 292384
rect 498048 292294 498118 292350
rect 498174 292294 498242 292350
rect 498298 292294 498368 292350
rect 498048 292226 498368 292294
rect 498048 292170 498118 292226
rect 498174 292170 498242 292226
rect 498298 292170 498368 292226
rect 498048 292102 498368 292170
rect 498048 292046 498118 292102
rect 498174 292046 498242 292102
rect 498298 292046 498368 292102
rect 498048 291978 498368 292046
rect 498048 291922 498118 291978
rect 498174 291922 498242 291978
rect 498298 291922 498368 291978
rect 498048 291888 498368 291922
rect 528768 292350 529088 292384
rect 528768 292294 528838 292350
rect 528894 292294 528962 292350
rect 529018 292294 529088 292350
rect 528768 292226 529088 292294
rect 528768 292170 528838 292226
rect 528894 292170 528962 292226
rect 529018 292170 529088 292226
rect 528768 292102 529088 292170
rect 528768 292046 528838 292102
rect 528894 292046 528962 292102
rect 529018 292046 529088 292102
rect 528768 291978 529088 292046
rect 528768 291922 528838 291978
rect 528894 291922 528962 291978
rect 529018 291922 529088 291978
rect 528768 291888 529088 291922
rect 559488 292350 559808 292384
rect 559488 292294 559558 292350
rect 559614 292294 559682 292350
rect 559738 292294 559808 292350
rect 559488 292226 559808 292294
rect 559488 292170 559558 292226
rect 559614 292170 559682 292226
rect 559738 292170 559808 292226
rect 559488 292102 559808 292170
rect 559488 292046 559558 292102
rect 559614 292046 559682 292102
rect 559738 292046 559808 292102
rect 559488 291978 559808 292046
rect 559488 291922 559558 291978
rect 559614 291922 559682 291978
rect 559738 291922 559808 291978
rect 559488 291888 559808 291922
rect 589098 292350 589718 309922
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 341068 283732 341124 283742
rect 341292 283978 341348 283988
rect 341068 243478 341124 243488
rect 341068 236098 341124 243422
rect 341292 239338 341348 283922
rect 359808 280350 360128 280384
rect 359808 280294 359878 280350
rect 359934 280294 360002 280350
rect 360058 280294 360128 280350
rect 359808 280226 360128 280294
rect 359808 280170 359878 280226
rect 359934 280170 360002 280226
rect 360058 280170 360128 280226
rect 359808 280102 360128 280170
rect 359808 280046 359878 280102
rect 359934 280046 360002 280102
rect 360058 280046 360128 280102
rect 359808 279978 360128 280046
rect 359808 279922 359878 279978
rect 359934 279922 360002 279978
rect 360058 279922 360128 279978
rect 359808 279888 360128 279922
rect 390528 280350 390848 280384
rect 390528 280294 390598 280350
rect 390654 280294 390722 280350
rect 390778 280294 390848 280350
rect 390528 280226 390848 280294
rect 390528 280170 390598 280226
rect 390654 280170 390722 280226
rect 390778 280170 390848 280226
rect 390528 280102 390848 280170
rect 390528 280046 390598 280102
rect 390654 280046 390722 280102
rect 390778 280046 390848 280102
rect 390528 279978 390848 280046
rect 390528 279922 390598 279978
rect 390654 279922 390722 279978
rect 390778 279922 390848 279978
rect 390528 279888 390848 279922
rect 421248 280350 421568 280384
rect 421248 280294 421318 280350
rect 421374 280294 421442 280350
rect 421498 280294 421568 280350
rect 421248 280226 421568 280294
rect 421248 280170 421318 280226
rect 421374 280170 421442 280226
rect 421498 280170 421568 280226
rect 421248 280102 421568 280170
rect 421248 280046 421318 280102
rect 421374 280046 421442 280102
rect 421498 280046 421568 280102
rect 421248 279978 421568 280046
rect 421248 279922 421318 279978
rect 421374 279922 421442 279978
rect 421498 279922 421568 279978
rect 421248 279888 421568 279922
rect 451968 280350 452288 280384
rect 451968 280294 452038 280350
rect 452094 280294 452162 280350
rect 452218 280294 452288 280350
rect 451968 280226 452288 280294
rect 451968 280170 452038 280226
rect 452094 280170 452162 280226
rect 452218 280170 452288 280226
rect 451968 280102 452288 280170
rect 451968 280046 452038 280102
rect 452094 280046 452162 280102
rect 452218 280046 452288 280102
rect 451968 279978 452288 280046
rect 451968 279922 452038 279978
rect 452094 279922 452162 279978
rect 452218 279922 452288 279978
rect 451968 279888 452288 279922
rect 482688 280350 483008 280384
rect 482688 280294 482758 280350
rect 482814 280294 482882 280350
rect 482938 280294 483008 280350
rect 482688 280226 483008 280294
rect 482688 280170 482758 280226
rect 482814 280170 482882 280226
rect 482938 280170 483008 280226
rect 482688 280102 483008 280170
rect 482688 280046 482758 280102
rect 482814 280046 482882 280102
rect 482938 280046 483008 280102
rect 482688 279978 483008 280046
rect 482688 279922 482758 279978
rect 482814 279922 482882 279978
rect 482938 279922 483008 279978
rect 482688 279888 483008 279922
rect 513408 280350 513728 280384
rect 513408 280294 513478 280350
rect 513534 280294 513602 280350
rect 513658 280294 513728 280350
rect 513408 280226 513728 280294
rect 513408 280170 513478 280226
rect 513534 280170 513602 280226
rect 513658 280170 513728 280226
rect 513408 280102 513728 280170
rect 513408 280046 513478 280102
rect 513534 280046 513602 280102
rect 513658 280046 513728 280102
rect 513408 279978 513728 280046
rect 513408 279922 513478 279978
rect 513534 279922 513602 279978
rect 513658 279922 513728 279978
rect 513408 279888 513728 279922
rect 544128 280350 544448 280384
rect 544128 280294 544198 280350
rect 544254 280294 544322 280350
rect 544378 280294 544448 280350
rect 544128 280226 544448 280294
rect 544128 280170 544198 280226
rect 544254 280170 544322 280226
rect 544378 280170 544448 280226
rect 544128 280102 544448 280170
rect 544128 280046 544198 280102
rect 544254 280046 544322 280102
rect 544378 280046 544448 280102
rect 544128 279978 544448 280046
rect 544128 279922 544198 279978
rect 544254 279922 544322 279978
rect 544378 279922 544448 279978
rect 544128 279888 544448 279922
rect 574848 280350 575168 280384
rect 574848 280294 574918 280350
rect 574974 280294 575042 280350
rect 575098 280294 575168 280350
rect 574848 280226 575168 280294
rect 574848 280170 574918 280226
rect 574974 280170 575042 280226
rect 575098 280170 575168 280226
rect 574848 280102 575168 280170
rect 574848 280046 574918 280102
rect 574974 280046 575042 280102
rect 575098 280046 575168 280102
rect 574848 279978 575168 280046
rect 574848 279922 574918 279978
rect 574974 279922 575042 279978
rect 575098 279922 575168 279978
rect 574848 279888 575168 279922
rect 344448 274350 344768 274384
rect 344448 274294 344518 274350
rect 344574 274294 344642 274350
rect 344698 274294 344768 274350
rect 344448 274226 344768 274294
rect 344448 274170 344518 274226
rect 344574 274170 344642 274226
rect 344698 274170 344768 274226
rect 344448 274102 344768 274170
rect 344448 274046 344518 274102
rect 344574 274046 344642 274102
rect 344698 274046 344768 274102
rect 344448 273978 344768 274046
rect 344448 273922 344518 273978
rect 344574 273922 344642 273978
rect 344698 273922 344768 273978
rect 344448 273888 344768 273922
rect 375168 274350 375488 274384
rect 375168 274294 375238 274350
rect 375294 274294 375362 274350
rect 375418 274294 375488 274350
rect 375168 274226 375488 274294
rect 375168 274170 375238 274226
rect 375294 274170 375362 274226
rect 375418 274170 375488 274226
rect 375168 274102 375488 274170
rect 375168 274046 375238 274102
rect 375294 274046 375362 274102
rect 375418 274046 375488 274102
rect 375168 273978 375488 274046
rect 375168 273922 375238 273978
rect 375294 273922 375362 273978
rect 375418 273922 375488 273978
rect 375168 273888 375488 273922
rect 405888 274350 406208 274384
rect 405888 274294 405958 274350
rect 406014 274294 406082 274350
rect 406138 274294 406208 274350
rect 405888 274226 406208 274294
rect 405888 274170 405958 274226
rect 406014 274170 406082 274226
rect 406138 274170 406208 274226
rect 405888 274102 406208 274170
rect 405888 274046 405958 274102
rect 406014 274046 406082 274102
rect 406138 274046 406208 274102
rect 405888 273978 406208 274046
rect 405888 273922 405958 273978
rect 406014 273922 406082 273978
rect 406138 273922 406208 273978
rect 405888 273888 406208 273922
rect 436608 274350 436928 274384
rect 436608 274294 436678 274350
rect 436734 274294 436802 274350
rect 436858 274294 436928 274350
rect 436608 274226 436928 274294
rect 436608 274170 436678 274226
rect 436734 274170 436802 274226
rect 436858 274170 436928 274226
rect 436608 274102 436928 274170
rect 436608 274046 436678 274102
rect 436734 274046 436802 274102
rect 436858 274046 436928 274102
rect 436608 273978 436928 274046
rect 436608 273922 436678 273978
rect 436734 273922 436802 273978
rect 436858 273922 436928 273978
rect 436608 273888 436928 273922
rect 467328 274350 467648 274384
rect 467328 274294 467398 274350
rect 467454 274294 467522 274350
rect 467578 274294 467648 274350
rect 467328 274226 467648 274294
rect 467328 274170 467398 274226
rect 467454 274170 467522 274226
rect 467578 274170 467648 274226
rect 467328 274102 467648 274170
rect 467328 274046 467398 274102
rect 467454 274046 467522 274102
rect 467578 274046 467648 274102
rect 467328 273978 467648 274046
rect 467328 273922 467398 273978
rect 467454 273922 467522 273978
rect 467578 273922 467648 273978
rect 467328 273888 467648 273922
rect 498048 274350 498368 274384
rect 498048 274294 498118 274350
rect 498174 274294 498242 274350
rect 498298 274294 498368 274350
rect 498048 274226 498368 274294
rect 498048 274170 498118 274226
rect 498174 274170 498242 274226
rect 498298 274170 498368 274226
rect 498048 274102 498368 274170
rect 498048 274046 498118 274102
rect 498174 274046 498242 274102
rect 498298 274046 498368 274102
rect 498048 273978 498368 274046
rect 498048 273922 498118 273978
rect 498174 273922 498242 273978
rect 498298 273922 498368 273978
rect 498048 273888 498368 273922
rect 528768 274350 529088 274384
rect 528768 274294 528838 274350
rect 528894 274294 528962 274350
rect 529018 274294 529088 274350
rect 528768 274226 529088 274294
rect 528768 274170 528838 274226
rect 528894 274170 528962 274226
rect 529018 274170 529088 274226
rect 528768 274102 529088 274170
rect 528768 274046 528838 274102
rect 528894 274046 528962 274102
rect 529018 274046 529088 274102
rect 528768 273978 529088 274046
rect 528768 273922 528838 273978
rect 528894 273922 528962 273978
rect 529018 273922 529088 273978
rect 528768 273888 529088 273922
rect 559488 274350 559808 274384
rect 559488 274294 559558 274350
rect 559614 274294 559682 274350
rect 559738 274294 559808 274350
rect 559488 274226 559808 274294
rect 559488 274170 559558 274226
rect 559614 274170 559682 274226
rect 559738 274170 559808 274226
rect 559488 274102 559808 274170
rect 559488 274046 559558 274102
rect 559614 274046 559682 274102
rect 559738 274046 559808 274102
rect 559488 273978 559808 274046
rect 559488 273922 559558 273978
rect 559614 273922 559682 273978
rect 559738 273922 559808 273978
rect 559488 273888 559808 273922
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 359808 262350 360128 262384
rect 359808 262294 359878 262350
rect 359934 262294 360002 262350
rect 360058 262294 360128 262350
rect 359808 262226 360128 262294
rect 359808 262170 359878 262226
rect 359934 262170 360002 262226
rect 360058 262170 360128 262226
rect 359808 262102 360128 262170
rect 359808 262046 359878 262102
rect 359934 262046 360002 262102
rect 360058 262046 360128 262102
rect 359808 261978 360128 262046
rect 359808 261922 359878 261978
rect 359934 261922 360002 261978
rect 360058 261922 360128 261978
rect 359808 261888 360128 261922
rect 390528 262350 390848 262384
rect 390528 262294 390598 262350
rect 390654 262294 390722 262350
rect 390778 262294 390848 262350
rect 390528 262226 390848 262294
rect 390528 262170 390598 262226
rect 390654 262170 390722 262226
rect 390778 262170 390848 262226
rect 390528 262102 390848 262170
rect 390528 262046 390598 262102
rect 390654 262046 390722 262102
rect 390778 262046 390848 262102
rect 390528 261978 390848 262046
rect 390528 261922 390598 261978
rect 390654 261922 390722 261978
rect 390778 261922 390848 261978
rect 390528 261888 390848 261922
rect 421248 262350 421568 262384
rect 421248 262294 421318 262350
rect 421374 262294 421442 262350
rect 421498 262294 421568 262350
rect 421248 262226 421568 262294
rect 421248 262170 421318 262226
rect 421374 262170 421442 262226
rect 421498 262170 421568 262226
rect 421248 262102 421568 262170
rect 421248 262046 421318 262102
rect 421374 262046 421442 262102
rect 421498 262046 421568 262102
rect 421248 261978 421568 262046
rect 421248 261922 421318 261978
rect 421374 261922 421442 261978
rect 421498 261922 421568 261978
rect 421248 261888 421568 261922
rect 451968 262350 452288 262384
rect 451968 262294 452038 262350
rect 452094 262294 452162 262350
rect 452218 262294 452288 262350
rect 451968 262226 452288 262294
rect 451968 262170 452038 262226
rect 452094 262170 452162 262226
rect 452218 262170 452288 262226
rect 451968 262102 452288 262170
rect 451968 262046 452038 262102
rect 452094 262046 452162 262102
rect 452218 262046 452288 262102
rect 451968 261978 452288 262046
rect 451968 261922 452038 261978
rect 452094 261922 452162 261978
rect 452218 261922 452288 261978
rect 451968 261888 452288 261922
rect 482688 262350 483008 262384
rect 482688 262294 482758 262350
rect 482814 262294 482882 262350
rect 482938 262294 483008 262350
rect 482688 262226 483008 262294
rect 482688 262170 482758 262226
rect 482814 262170 482882 262226
rect 482938 262170 483008 262226
rect 482688 262102 483008 262170
rect 482688 262046 482758 262102
rect 482814 262046 482882 262102
rect 482938 262046 483008 262102
rect 482688 261978 483008 262046
rect 482688 261922 482758 261978
rect 482814 261922 482882 261978
rect 482938 261922 483008 261978
rect 482688 261888 483008 261922
rect 513408 262350 513728 262384
rect 513408 262294 513478 262350
rect 513534 262294 513602 262350
rect 513658 262294 513728 262350
rect 513408 262226 513728 262294
rect 513408 262170 513478 262226
rect 513534 262170 513602 262226
rect 513658 262170 513728 262226
rect 513408 262102 513728 262170
rect 513408 262046 513478 262102
rect 513534 262046 513602 262102
rect 513658 262046 513728 262102
rect 513408 261978 513728 262046
rect 513408 261922 513478 261978
rect 513534 261922 513602 261978
rect 513658 261922 513728 261978
rect 513408 261888 513728 261922
rect 544128 262350 544448 262384
rect 544128 262294 544198 262350
rect 544254 262294 544322 262350
rect 544378 262294 544448 262350
rect 544128 262226 544448 262294
rect 544128 262170 544198 262226
rect 544254 262170 544322 262226
rect 544378 262170 544448 262226
rect 544128 262102 544448 262170
rect 544128 262046 544198 262102
rect 544254 262046 544322 262102
rect 544378 262046 544448 262102
rect 544128 261978 544448 262046
rect 544128 261922 544198 261978
rect 544254 261922 544322 261978
rect 544378 261922 544448 261978
rect 544128 261888 544448 261922
rect 574848 262350 575168 262384
rect 574848 262294 574918 262350
rect 574974 262294 575042 262350
rect 575098 262294 575168 262350
rect 574848 262226 575168 262294
rect 574848 262170 574918 262226
rect 574974 262170 575042 262226
rect 575098 262170 575168 262226
rect 574848 262102 575168 262170
rect 574848 262046 574918 262102
rect 574974 262046 575042 262102
rect 575098 262046 575168 262102
rect 574848 261978 575168 262046
rect 574848 261922 574918 261978
rect 574974 261922 575042 261978
rect 575098 261922 575168 261978
rect 574848 261888 575168 261922
rect 344448 256350 344768 256384
rect 344448 256294 344518 256350
rect 344574 256294 344642 256350
rect 344698 256294 344768 256350
rect 344448 256226 344768 256294
rect 344448 256170 344518 256226
rect 344574 256170 344642 256226
rect 344698 256170 344768 256226
rect 344448 256102 344768 256170
rect 344448 256046 344518 256102
rect 344574 256046 344642 256102
rect 344698 256046 344768 256102
rect 344448 255978 344768 256046
rect 344448 255922 344518 255978
rect 344574 255922 344642 255978
rect 344698 255922 344768 255978
rect 344448 255888 344768 255922
rect 375168 256350 375488 256384
rect 375168 256294 375238 256350
rect 375294 256294 375362 256350
rect 375418 256294 375488 256350
rect 375168 256226 375488 256294
rect 375168 256170 375238 256226
rect 375294 256170 375362 256226
rect 375418 256170 375488 256226
rect 375168 256102 375488 256170
rect 375168 256046 375238 256102
rect 375294 256046 375362 256102
rect 375418 256046 375488 256102
rect 375168 255978 375488 256046
rect 375168 255922 375238 255978
rect 375294 255922 375362 255978
rect 375418 255922 375488 255978
rect 375168 255888 375488 255922
rect 405888 256350 406208 256384
rect 405888 256294 405958 256350
rect 406014 256294 406082 256350
rect 406138 256294 406208 256350
rect 405888 256226 406208 256294
rect 405888 256170 405958 256226
rect 406014 256170 406082 256226
rect 406138 256170 406208 256226
rect 405888 256102 406208 256170
rect 405888 256046 405958 256102
rect 406014 256046 406082 256102
rect 406138 256046 406208 256102
rect 405888 255978 406208 256046
rect 405888 255922 405958 255978
rect 406014 255922 406082 255978
rect 406138 255922 406208 255978
rect 405888 255888 406208 255922
rect 436608 256350 436928 256384
rect 436608 256294 436678 256350
rect 436734 256294 436802 256350
rect 436858 256294 436928 256350
rect 436608 256226 436928 256294
rect 436608 256170 436678 256226
rect 436734 256170 436802 256226
rect 436858 256170 436928 256226
rect 436608 256102 436928 256170
rect 436608 256046 436678 256102
rect 436734 256046 436802 256102
rect 436858 256046 436928 256102
rect 436608 255978 436928 256046
rect 436608 255922 436678 255978
rect 436734 255922 436802 255978
rect 436858 255922 436928 255978
rect 436608 255888 436928 255922
rect 467328 256350 467648 256384
rect 467328 256294 467398 256350
rect 467454 256294 467522 256350
rect 467578 256294 467648 256350
rect 467328 256226 467648 256294
rect 467328 256170 467398 256226
rect 467454 256170 467522 256226
rect 467578 256170 467648 256226
rect 467328 256102 467648 256170
rect 467328 256046 467398 256102
rect 467454 256046 467522 256102
rect 467578 256046 467648 256102
rect 467328 255978 467648 256046
rect 467328 255922 467398 255978
rect 467454 255922 467522 255978
rect 467578 255922 467648 255978
rect 467328 255888 467648 255922
rect 498048 256350 498368 256384
rect 498048 256294 498118 256350
rect 498174 256294 498242 256350
rect 498298 256294 498368 256350
rect 498048 256226 498368 256294
rect 498048 256170 498118 256226
rect 498174 256170 498242 256226
rect 498298 256170 498368 256226
rect 498048 256102 498368 256170
rect 498048 256046 498118 256102
rect 498174 256046 498242 256102
rect 498298 256046 498368 256102
rect 498048 255978 498368 256046
rect 498048 255922 498118 255978
rect 498174 255922 498242 255978
rect 498298 255922 498368 255978
rect 498048 255888 498368 255922
rect 528768 256350 529088 256384
rect 528768 256294 528838 256350
rect 528894 256294 528962 256350
rect 529018 256294 529088 256350
rect 528768 256226 529088 256294
rect 528768 256170 528838 256226
rect 528894 256170 528962 256226
rect 529018 256170 529088 256226
rect 528768 256102 529088 256170
rect 528768 256046 528838 256102
rect 528894 256046 528962 256102
rect 529018 256046 529088 256102
rect 528768 255978 529088 256046
rect 528768 255922 528838 255978
rect 528894 255922 528962 255978
rect 529018 255922 529088 255978
rect 528768 255888 529088 255922
rect 559488 256350 559808 256384
rect 559488 256294 559558 256350
rect 559614 256294 559682 256350
rect 559738 256294 559808 256350
rect 559488 256226 559808 256294
rect 559488 256170 559558 256226
rect 559614 256170 559682 256226
rect 559738 256170 559808 256226
rect 559488 256102 559808 256170
rect 559488 256046 559558 256102
rect 559614 256046 559682 256102
rect 559738 256046 559808 256102
rect 559488 255978 559808 256046
rect 559488 255922 559558 255978
rect 559614 255922 559682 255978
rect 559738 255922 559808 255978
rect 559488 255888 559808 255922
rect 589098 256350 589718 273922
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 359808 244350 360128 244384
rect 359808 244294 359878 244350
rect 359934 244294 360002 244350
rect 360058 244294 360128 244350
rect 359808 244226 360128 244294
rect 359808 244170 359878 244226
rect 359934 244170 360002 244226
rect 360058 244170 360128 244226
rect 359808 244102 360128 244170
rect 359808 244046 359878 244102
rect 359934 244046 360002 244102
rect 360058 244046 360128 244102
rect 359808 243978 360128 244046
rect 359808 243922 359878 243978
rect 359934 243922 360002 243978
rect 360058 243922 360128 243978
rect 359808 243888 360128 243922
rect 390528 244350 390848 244384
rect 390528 244294 390598 244350
rect 390654 244294 390722 244350
rect 390778 244294 390848 244350
rect 390528 244226 390848 244294
rect 390528 244170 390598 244226
rect 390654 244170 390722 244226
rect 390778 244170 390848 244226
rect 390528 244102 390848 244170
rect 390528 244046 390598 244102
rect 390654 244046 390722 244102
rect 390778 244046 390848 244102
rect 390528 243978 390848 244046
rect 390528 243922 390598 243978
rect 390654 243922 390722 243978
rect 390778 243922 390848 243978
rect 390528 243888 390848 243922
rect 421248 244350 421568 244384
rect 421248 244294 421318 244350
rect 421374 244294 421442 244350
rect 421498 244294 421568 244350
rect 421248 244226 421568 244294
rect 421248 244170 421318 244226
rect 421374 244170 421442 244226
rect 421498 244170 421568 244226
rect 421248 244102 421568 244170
rect 421248 244046 421318 244102
rect 421374 244046 421442 244102
rect 421498 244046 421568 244102
rect 421248 243978 421568 244046
rect 421248 243922 421318 243978
rect 421374 243922 421442 243978
rect 421498 243922 421568 243978
rect 421248 243888 421568 243922
rect 451968 244350 452288 244384
rect 451968 244294 452038 244350
rect 452094 244294 452162 244350
rect 452218 244294 452288 244350
rect 451968 244226 452288 244294
rect 451968 244170 452038 244226
rect 452094 244170 452162 244226
rect 452218 244170 452288 244226
rect 451968 244102 452288 244170
rect 451968 244046 452038 244102
rect 452094 244046 452162 244102
rect 452218 244046 452288 244102
rect 451968 243978 452288 244046
rect 451968 243922 452038 243978
rect 452094 243922 452162 243978
rect 452218 243922 452288 243978
rect 451968 243888 452288 243922
rect 482688 244350 483008 244384
rect 482688 244294 482758 244350
rect 482814 244294 482882 244350
rect 482938 244294 483008 244350
rect 482688 244226 483008 244294
rect 482688 244170 482758 244226
rect 482814 244170 482882 244226
rect 482938 244170 483008 244226
rect 482688 244102 483008 244170
rect 482688 244046 482758 244102
rect 482814 244046 482882 244102
rect 482938 244046 483008 244102
rect 482688 243978 483008 244046
rect 482688 243922 482758 243978
rect 482814 243922 482882 243978
rect 482938 243922 483008 243978
rect 482688 243888 483008 243922
rect 513408 244350 513728 244384
rect 513408 244294 513478 244350
rect 513534 244294 513602 244350
rect 513658 244294 513728 244350
rect 513408 244226 513728 244294
rect 513408 244170 513478 244226
rect 513534 244170 513602 244226
rect 513658 244170 513728 244226
rect 513408 244102 513728 244170
rect 513408 244046 513478 244102
rect 513534 244046 513602 244102
rect 513658 244046 513728 244102
rect 513408 243978 513728 244046
rect 513408 243922 513478 243978
rect 513534 243922 513602 243978
rect 513658 243922 513728 243978
rect 513408 243888 513728 243922
rect 544128 244350 544448 244384
rect 544128 244294 544198 244350
rect 544254 244294 544322 244350
rect 544378 244294 544448 244350
rect 544128 244226 544448 244294
rect 544128 244170 544198 244226
rect 544254 244170 544322 244226
rect 544378 244170 544448 244226
rect 544128 244102 544448 244170
rect 544128 244046 544198 244102
rect 544254 244046 544322 244102
rect 544378 244046 544448 244102
rect 544128 243978 544448 244046
rect 544128 243922 544198 243978
rect 544254 243922 544322 243978
rect 544378 243922 544448 243978
rect 544128 243888 544448 243922
rect 574848 244350 575168 244384
rect 574848 244294 574918 244350
rect 574974 244294 575042 244350
rect 575098 244294 575168 244350
rect 574848 244226 575168 244294
rect 574848 244170 574918 244226
rect 574974 244170 575042 244226
rect 575098 244170 575168 244226
rect 574848 244102 575168 244170
rect 574848 244046 574918 244102
rect 574974 244046 575042 244102
rect 575098 244046 575168 244102
rect 574848 243978 575168 244046
rect 574848 243922 574918 243978
rect 574974 243922 575042 243978
rect 575098 243922 575168 243978
rect 574848 243888 575168 243922
rect 341292 239272 341348 239282
rect 344448 238350 344768 238384
rect 344448 238294 344518 238350
rect 344574 238294 344642 238350
rect 344698 238294 344768 238350
rect 344448 238226 344768 238294
rect 344448 238170 344518 238226
rect 344574 238170 344642 238226
rect 344698 238170 344768 238226
rect 344448 238102 344768 238170
rect 344448 238046 344518 238102
rect 344574 238046 344642 238102
rect 344698 238046 344768 238102
rect 344448 237978 344768 238046
rect 344448 237922 344518 237978
rect 344574 237922 344642 237978
rect 344698 237922 344768 237978
rect 344448 237888 344768 237922
rect 375168 238350 375488 238384
rect 375168 238294 375238 238350
rect 375294 238294 375362 238350
rect 375418 238294 375488 238350
rect 375168 238226 375488 238294
rect 375168 238170 375238 238226
rect 375294 238170 375362 238226
rect 375418 238170 375488 238226
rect 375168 238102 375488 238170
rect 375168 238046 375238 238102
rect 375294 238046 375362 238102
rect 375418 238046 375488 238102
rect 375168 237978 375488 238046
rect 375168 237922 375238 237978
rect 375294 237922 375362 237978
rect 375418 237922 375488 237978
rect 375168 237888 375488 237922
rect 405888 238350 406208 238384
rect 405888 238294 405958 238350
rect 406014 238294 406082 238350
rect 406138 238294 406208 238350
rect 405888 238226 406208 238294
rect 405888 238170 405958 238226
rect 406014 238170 406082 238226
rect 406138 238170 406208 238226
rect 405888 238102 406208 238170
rect 405888 238046 405958 238102
rect 406014 238046 406082 238102
rect 406138 238046 406208 238102
rect 405888 237978 406208 238046
rect 405888 237922 405958 237978
rect 406014 237922 406082 237978
rect 406138 237922 406208 237978
rect 405888 237888 406208 237922
rect 436608 238350 436928 238384
rect 436608 238294 436678 238350
rect 436734 238294 436802 238350
rect 436858 238294 436928 238350
rect 436608 238226 436928 238294
rect 436608 238170 436678 238226
rect 436734 238170 436802 238226
rect 436858 238170 436928 238226
rect 436608 238102 436928 238170
rect 436608 238046 436678 238102
rect 436734 238046 436802 238102
rect 436858 238046 436928 238102
rect 436608 237978 436928 238046
rect 436608 237922 436678 237978
rect 436734 237922 436802 237978
rect 436858 237922 436928 237978
rect 436608 237888 436928 237922
rect 467328 238350 467648 238384
rect 467328 238294 467398 238350
rect 467454 238294 467522 238350
rect 467578 238294 467648 238350
rect 467328 238226 467648 238294
rect 467328 238170 467398 238226
rect 467454 238170 467522 238226
rect 467578 238170 467648 238226
rect 467328 238102 467648 238170
rect 467328 238046 467398 238102
rect 467454 238046 467522 238102
rect 467578 238046 467648 238102
rect 467328 237978 467648 238046
rect 467328 237922 467398 237978
rect 467454 237922 467522 237978
rect 467578 237922 467648 237978
rect 467328 237888 467648 237922
rect 498048 238350 498368 238384
rect 498048 238294 498118 238350
rect 498174 238294 498242 238350
rect 498298 238294 498368 238350
rect 498048 238226 498368 238294
rect 498048 238170 498118 238226
rect 498174 238170 498242 238226
rect 498298 238170 498368 238226
rect 498048 238102 498368 238170
rect 498048 238046 498118 238102
rect 498174 238046 498242 238102
rect 498298 238046 498368 238102
rect 498048 237978 498368 238046
rect 498048 237922 498118 237978
rect 498174 237922 498242 237978
rect 498298 237922 498368 237978
rect 498048 237888 498368 237922
rect 528768 238350 529088 238384
rect 528768 238294 528838 238350
rect 528894 238294 528962 238350
rect 529018 238294 529088 238350
rect 528768 238226 529088 238294
rect 528768 238170 528838 238226
rect 528894 238170 528962 238226
rect 529018 238170 529088 238226
rect 528768 238102 529088 238170
rect 528768 238046 528838 238102
rect 528894 238046 528962 238102
rect 529018 238046 529088 238102
rect 528768 237978 529088 238046
rect 528768 237922 528838 237978
rect 528894 237922 528962 237978
rect 529018 237922 529088 237978
rect 528768 237888 529088 237922
rect 559488 238350 559808 238384
rect 559488 238294 559558 238350
rect 559614 238294 559682 238350
rect 559738 238294 559808 238350
rect 559488 238226 559808 238294
rect 559488 238170 559558 238226
rect 559614 238170 559682 238226
rect 559738 238170 559808 238226
rect 559488 238102 559808 238170
rect 559488 238046 559558 238102
rect 559614 238046 559682 238102
rect 559738 238046 559808 238102
rect 559488 237978 559808 238046
rect 559488 237922 559558 237978
rect 559614 237922 559682 237978
rect 559738 237922 559808 237978
rect 559488 237888 559808 237922
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 341068 236032 341124 236042
rect 359808 226350 360128 226384
rect 359808 226294 359878 226350
rect 359934 226294 360002 226350
rect 360058 226294 360128 226350
rect 359808 226226 360128 226294
rect 359808 226170 359878 226226
rect 359934 226170 360002 226226
rect 360058 226170 360128 226226
rect 359808 226102 360128 226170
rect 359808 226046 359878 226102
rect 359934 226046 360002 226102
rect 360058 226046 360128 226102
rect 359808 225978 360128 226046
rect 359808 225922 359878 225978
rect 359934 225922 360002 225978
rect 360058 225922 360128 225978
rect 359808 225888 360128 225922
rect 390528 226350 390848 226384
rect 390528 226294 390598 226350
rect 390654 226294 390722 226350
rect 390778 226294 390848 226350
rect 390528 226226 390848 226294
rect 390528 226170 390598 226226
rect 390654 226170 390722 226226
rect 390778 226170 390848 226226
rect 390528 226102 390848 226170
rect 390528 226046 390598 226102
rect 390654 226046 390722 226102
rect 390778 226046 390848 226102
rect 390528 225978 390848 226046
rect 390528 225922 390598 225978
rect 390654 225922 390722 225978
rect 390778 225922 390848 225978
rect 390528 225888 390848 225922
rect 421248 226350 421568 226384
rect 421248 226294 421318 226350
rect 421374 226294 421442 226350
rect 421498 226294 421568 226350
rect 421248 226226 421568 226294
rect 421248 226170 421318 226226
rect 421374 226170 421442 226226
rect 421498 226170 421568 226226
rect 421248 226102 421568 226170
rect 421248 226046 421318 226102
rect 421374 226046 421442 226102
rect 421498 226046 421568 226102
rect 421248 225978 421568 226046
rect 421248 225922 421318 225978
rect 421374 225922 421442 225978
rect 421498 225922 421568 225978
rect 421248 225888 421568 225922
rect 451968 226350 452288 226384
rect 451968 226294 452038 226350
rect 452094 226294 452162 226350
rect 452218 226294 452288 226350
rect 451968 226226 452288 226294
rect 451968 226170 452038 226226
rect 452094 226170 452162 226226
rect 452218 226170 452288 226226
rect 451968 226102 452288 226170
rect 451968 226046 452038 226102
rect 452094 226046 452162 226102
rect 452218 226046 452288 226102
rect 451968 225978 452288 226046
rect 451968 225922 452038 225978
rect 452094 225922 452162 225978
rect 452218 225922 452288 225978
rect 451968 225888 452288 225922
rect 482688 226350 483008 226384
rect 482688 226294 482758 226350
rect 482814 226294 482882 226350
rect 482938 226294 483008 226350
rect 482688 226226 483008 226294
rect 482688 226170 482758 226226
rect 482814 226170 482882 226226
rect 482938 226170 483008 226226
rect 482688 226102 483008 226170
rect 482688 226046 482758 226102
rect 482814 226046 482882 226102
rect 482938 226046 483008 226102
rect 482688 225978 483008 226046
rect 482688 225922 482758 225978
rect 482814 225922 482882 225978
rect 482938 225922 483008 225978
rect 482688 225888 483008 225922
rect 513408 226350 513728 226384
rect 513408 226294 513478 226350
rect 513534 226294 513602 226350
rect 513658 226294 513728 226350
rect 513408 226226 513728 226294
rect 513408 226170 513478 226226
rect 513534 226170 513602 226226
rect 513658 226170 513728 226226
rect 513408 226102 513728 226170
rect 513408 226046 513478 226102
rect 513534 226046 513602 226102
rect 513658 226046 513728 226102
rect 513408 225978 513728 226046
rect 513408 225922 513478 225978
rect 513534 225922 513602 225978
rect 513658 225922 513728 225978
rect 513408 225888 513728 225922
rect 544128 226350 544448 226384
rect 544128 226294 544198 226350
rect 544254 226294 544322 226350
rect 544378 226294 544448 226350
rect 544128 226226 544448 226294
rect 544128 226170 544198 226226
rect 544254 226170 544322 226226
rect 544378 226170 544448 226226
rect 544128 226102 544448 226170
rect 544128 226046 544198 226102
rect 544254 226046 544322 226102
rect 544378 226046 544448 226102
rect 544128 225978 544448 226046
rect 544128 225922 544198 225978
rect 544254 225922 544322 225978
rect 544378 225922 544448 225978
rect 544128 225888 544448 225922
rect 574848 226350 575168 226384
rect 574848 226294 574918 226350
rect 574974 226294 575042 226350
rect 575098 226294 575168 226350
rect 574848 226226 575168 226294
rect 574848 226170 574918 226226
rect 574974 226170 575042 226226
rect 575098 226170 575168 226226
rect 574848 226102 575168 226170
rect 574848 226046 574918 226102
rect 574974 226046 575042 226102
rect 575098 226046 575168 226102
rect 574848 225978 575168 226046
rect 574848 225922 574918 225978
rect 574974 225922 575042 225978
rect 575098 225922 575168 225978
rect 574848 225888 575168 225922
rect 344448 220350 344768 220384
rect 344448 220294 344518 220350
rect 344574 220294 344642 220350
rect 344698 220294 344768 220350
rect 344448 220226 344768 220294
rect 344448 220170 344518 220226
rect 344574 220170 344642 220226
rect 344698 220170 344768 220226
rect 344448 220102 344768 220170
rect 344448 220046 344518 220102
rect 344574 220046 344642 220102
rect 344698 220046 344768 220102
rect 344448 219978 344768 220046
rect 344448 219922 344518 219978
rect 344574 219922 344642 219978
rect 344698 219922 344768 219978
rect 344448 219888 344768 219922
rect 375168 220350 375488 220384
rect 375168 220294 375238 220350
rect 375294 220294 375362 220350
rect 375418 220294 375488 220350
rect 375168 220226 375488 220294
rect 375168 220170 375238 220226
rect 375294 220170 375362 220226
rect 375418 220170 375488 220226
rect 375168 220102 375488 220170
rect 375168 220046 375238 220102
rect 375294 220046 375362 220102
rect 375418 220046 375488 220102
rect 375168 219978 375488 220046
rect 375168 219922 375238 219978
rect 375294 219922 375362 219978
rect 375418 219922 375488 219978
rect 375168 219888 375488 219922
rect 405888 220350 406208 220384
rect 405888 220294 405958 220350
rect 406014 220294 406082 220350
rect 406138 220294 406208 220350
rect 405888 220226 406208 220294
rect 405888 220170 405958 220226
rect 406014 220170 406082 220226
rect 406138 220170 406208 220226
rect 405888 220102 406208 220170
rect 405888 220046 405958 220102
rect 406014 220046 406082 220102
rect 406138 220046 406208 220102
rect 405888 219978 406208 220046
rect 405888 219922 405958 219978
rect 406014 219922 406082 219978
rect 406138 219922 406208 219978
rect 405888 219888 406208 219922
rect 436608 220350 436928 220384
rect 436608 220294 436678 220350
rect 436734 220294 436802 220350
rect 436858 220294 436928 220350
rect 436608 220226 436928 220294
rect 436608 220170 436678 220226
rect 436734 220170 436802 220226
rect 436858 220170 436928 220226
rect 436608 220102 436928 220170
rect 436608 220046 436678 220102
rect 436734 220046 436802 220102
rect 436858 220046 436928 220102
rect 436608 219978 436928 220046
rect 436608 219922 436678 219978
rect 436734 219922 436802 219978
rect 436858 219922 436928 219978
rect 436608 219888 436928 219922
rect 467328 220350 467648 220384
rect 467328 220294 467398 220350
rect 467454 220294 467522 220350
rect 467578 220294 467648 220350
rect 467328 220226 467648 220294
rect 467328 220170 467398 220226
rect 467454 220170 467522 220226
rect 467578 220170 467648 220226
rect 467328 220102 467648 220170
rect 467328 220046 467398 220102
rect 467454 220046 467522 220102
rect 467578 220046 467648 220102
rect 467328 219978 467648 220046
rect 467328 219922 467398 219978
rect 467454 219922 467522 219978
rect 467578 219922 467648 219978
rect 467328 219888 467648 219922
rect 498048 220350 498368 220384
rect 498048 220294 498118 220350
rect 498174 220294 498242 220350
rect 498298 220294 498368 220350
rect 498048 220226 498368 220294
rect 498048 220170 498118 220226
rect 498174 220170 498242 220226
rect 498298 220170 498368 220226
rect 498048 220102 498368 220170
rect 498048 220046 498118 220102
rect 498174 220046 498242 220102
rect 498298 220046 498368 220102
rect 498048 219978 498368 220046
rect 498048 219922 498118 219978
rect 498174 219922 498242 219978
rect 498298 219922 498368 219978
rect 498048 219888 498368 219922
rect 528768 220350 529088 220384
rect 528768 220294 528838 220350
rect 528894 220294 528962 220350
rect 529018 220294 529088 220350
rect 528768 220226 529088 220294
rect 528768 220170 528838 220226
rect 528894 220170 528962 220226
rect 529018 220170 529088 220226
rect 528768 220102 529088 220170
rect 528768 220046 528838 220102
rect 528894 220046 528962 220102
rect 529018 220046 529088 220102
rect 528768 219978 529088 220046
rect 528768 219922 528838 219978
rect 528894 219922 528962 219978
rect 529018 219922 529088 219978
rect 528768 219888 529088 219922
rect 559488 220350 559808 220384
rect 559488 220294 559558 220350
rect 559614 220294 559682 220350
rect 559738 220294 559808 220350
rect 559488 220226 559808 220294
rect 559488 220170 559558 220226
rect 559614 220170 559682 220226
rect 559738 220170 559808 220226
rect 559488 220102 559808 220170
rect 559488 220046 559558 220102
rect 559614 220046 559682 220102
rect 559738 220046 559808 220102
rect 559488 219978 559808 220046
rect 559488 219922 559558 219978
rect 559614 219922 559682 219978
rect 559738 219922 559808 219978
rect 559488 219888 559808 219922
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 359808 208350 360128 208384
rect 359808 208294 359878 208350
rect 359934 208294 360002 208350
rect 360058 208294 360128 208350
rect 359808 208226 360128 208294
rect 359808 208170 359878 208226
rect 359934 208170 360002 208226
rect 360058 208170 360128 208226
rect 359808 208102 360128 208170
rect 359808 208046 359878 208102
rect 359934 208046 360002 208102
rect 360058 208046 360128 208102
rect 359808 207978 360128 208046
rect 359808 207922 359878 207978
rect 359934 207922 360002 207978
rect 360058 207922 360128 207978
rect 359808 207888 360128 207922
rect 390528 208350 390848 208384
rect 390528 208294 390598 208350
rect 390654 208294 390722 208350
rect 390778 208294 390848 208350
rect 390528 208226 390848 208294
rect 390528 208170 390598 208226
rect 390654 208170 390722 208226
rect 390778 208170 390848 208226
rect 390528 208102 390848 208170
rect 390528 208046 390598 208102
rect 390654 208046 390722 208102
rect 390778 208046 390848 208102
rect 390528 207978 390848 208046
rect 390528 207922 390598 207978
rect 390654 207922 390722 207978
rect 390778 207922 390848 207978
rect 390528 207888 390848 207922
rect 421248 208350 421568 208384
rect 421248 208294 421318 208350
rect 421374 208294 421442 208350
rect 421498 208294 421568 208350
rect 421248 208226 421568 208294
rect 421248 208170 421318 208226
rect 421374 208170 421442 208226
rect 421498 208170 421568 208226
rect 421248 208102 421568 208170
rect 421248 208046 421318 208102
rect 421374 208046 421442 208102
rect 421498 208046 421568 208102
rect 421248 207978 421568 208046
rect 421248 207922 421318 207978
rect 421374 207922 421442 207978
rect 421498 207922 421568 207978
rect 421248 207888 421568 207922
rect 451968 208350 452288 208384
rect 451968 208294 452038 208350
rect 452094 208294 452162 208350
rect 452218 208294 452288 208350
rect 451968 208226 452288 208294
rect 451968 208170 452038 208226
rect 452094 208170 452162 208226
rect 452218 208170 452288 208226
rect 451968 208102 452288 208170
rect 451968 208046 452038 208102
rect 452094 208046 452162 208102
rect 452218 208046 452288 208102
rect 451968 207978 452288 208046
rect 451968 207922 452038 207978
rect 452094 207922 452162 207978
rect 452218 207922 452288 207978
rect 451968 207888 452288 207922
rect 482688 208350 483008 208384
rect 482688 208294 482758 208350
rect 482814 208294 482882 208350
rect 482938 208294 483008 208350
rect 482688 208226 483008 208294
rect 482688 208170 482758 208226
rect 482814 208170 482882 208226
rect 482938 208170 483008 208226
rect 482688 208102 483008 208170
rect 482688 208046 482758 208102
rect 482814 208046 482882 208102
rect 482938 208046 483008 208102
rect 482688 207978 483008 208046
rect 482688 207922 482758 207978
rect 482814 207922 482882 207978
rect 482938 207922 483008 207978
rect 482688 207888 483008 207922
rect 513408 208350 513728 208384
rect 513408 208294 513478 208350
rect 513534 208294 513602 208350
rect 513658 208294 513728 208350
rect 513408 208226 513728 208294
rect 513408 208170 513478 208226
rect 513534 208170 513602 208226
rect 513658 208170 513728 208226
rect 513408 208102 513728 208170
rect 513408 208046 513478 208102
rect 513534 208046 513602 208102
rect 513658 208046 513728 208102
rect 513408 207978 513728 208046
rect 513408 207922 513478 207978
rect 513534 207922 513602 207978
rect 513658 207922 513728 207978
rect 513408 207888 513728 207922
rect 544128 208350 544448 208384
rect 544128 208294 544198 208350
rect 544254 208294 544322 208350
rect 544378 208294 544448 208350
rect 544128 208226 544448 208294
rect 544128 208170 544198 208226
rect 544254 208170 544322 208226
rect 544378 208170 544448 208226
rect 544128 208102 544448 208170
rect 544128 208046 544198 208102
rect 544254 208046 544322 208102
rect 544378 208046 544448 208102
rect 544128 207978 544448 208046
rect 544128 207922 544198 207978
rect 544254 207922 544322 207978
rect 544378 207922 544448 207978
rect 544128 207888 544448 207922
rect 574848 208350 575168 208384
rect 574848 208294 574918 208350
rect 574974 208294 575042 208350
rect 575098 208294 575168 208350
rect 574848 208226 575168 208294
rect 574848 208170 574918 208226
rect 574974 208170 575042 208226
rect 575098 208170 575168 208226
rect 574848 208102 575168 208170
rect 574848 208046 574918 208102
rect 574974 208046 575042 208102
rect 575098 208046 575168 208102
rect 574848 207978 575168 208046
rect 574848 207922 574918 207978
rect 574974 207922 575042 207978
rect 575098 207922 575168 207978
rect 574848 207888 575168 207922
rect 344448 202350 344768 202384
rect 344448 202294 344518 202350
rect 344574 202294 344642 202350
rect 344698 202294 344768 202350
rect 344448 202226 344768 202294
rect 344448 202170 344518 202226
rect 344574 202170 344642 202226
rect 344698 202170 344768 202226
rect 344448 202102 344768 202170
rect 344448 202046 344518 202102
rect 344574 202046 344642 202102
rect 344698 202046 344768 202102
rect 344448 201978 344768 202046
rect 344448 201922 344518 201978
rect 344574 201922 344642 201978
rect 344698 201922 344768 201978
rect 344448 201888 344768 201922
rect 375168 202350 375488 202384
rect 375168 202294 375238 202350
rect 375294 202294 375362 202350
rect 375418 202294 375488 202350
rect 375168 202226 375488 202294
rect 375168 202170 375238 202226
rect 375294 202170 375362 202226
rect 375418 202170 375488 202226
rect 375168 202102 375488 202170
rect 375168 202046 375238 202102
rect 375294 202046 375362 202102
rect 375418 202046 375488 202102
rect 375168 201978 375488 202046
rect 375168 201922 375238 201978
rect 375294 201922 375362 201978
rect 375418 201922 375488 201978
rect 375168 201888 375488 201922
rect 405888 202350 406208 202384
rect 405888 202294 405958 202350
rect 406014 202294 406082 202350
rect 406138 202294 406208 202350
rect 405888 202226 406208 202294
rect 405888 202170 405958 202226
rect 406014 202170 406082 202226
rect 406138 202170 406208 202226
rect 405888 202102 406208 202170
rect 405888 202046 405958 202102
rect 406014 202046 406082 202102
rect 406138 202046 406208 202102
rect 405888 201978 406208 202046
rect 405888 201922 405958 201978
rect 406014 201922 406082 201978
rect 406138 201922 406208 201978
rect 405888 201888 406208 201922
rect 436608 202350 436928 202384
rect 436608 202294 436678 202350
rect 436734 202294 436802 202350
rect 436858 202294 436928 202350
rect 436608 202226 436928 202294
rect 436608 202170 436678 202226
rect 436734 202170 436802 202226
rect 436858 202170 436928 202226
rect 436608 202102 436928 202170
rect 436608 202046 436678 202102
rect 436734 202046 436802 202102
rect 436858 202046 436928 202102
rect 436608 201978 436928 202046
rect 436608 201922 436678 201978
rect 436734 201922 436802 201978
rect 436858 201922 436928 201978
rect 436608 201888 436928 201922
rect 467328 202350 467648 202384
rect 467328 202294 467398 202350
rect 467454 202294 467522 202350
rect 467578 202294 467648 202350
rect 467328 202226 467648 202294
rect 467328 202170 467398 202226
rect 467454 202170 467522 202226
rect 467578 202170 467648 202226
rect 467328 202102 467648 202170
rect 467328 202046 467398 202102
rect 467454 202046 467522 202102
rect 467578 202046 467648 202102
rect 467328 201978 467648 202046
rect 467328 201922 467398 201978
rect 467454 201922 467522 201978
rect 467578 201922 467648 201978
rect 467328 201888 467648 201922
rect 498048 202350 498368 202384
rect 498048 202294 498118 202350
rect 498174 202294 498242 202350
rect 498298 202294 498368 202350
rect 498048 202226 498368 202294
rect 498048 202170 498118 202226
rect 498174 202170 498242 202226
rect 498298 202170 498368 202226
rect 498048 202102 498368 202170
rect 498048 202046 498118 202102
rect 498174 202046 498242 202102
rect 498298 202046 498368 202102
rect 498048 201978 498368 202046
rect 498048 201922 498118 201978
rect 498174 201922 498242 201978
rect 498298 201922 498368 201978
rect 498048 201888 498368 201922
rect 528768 202350 529088 202384
rect 528768 202294 528838 202350
rect 528894 202294 528962 202350
rect 529018 202294 529088 202350
rect 528768 202226 529088 202294
rect 528768 202170 528838 202226
rect 528894 202170 528962 202226
rect 529018 202170 529088 202226
rect 528768 202102 529088 202170
rect 528768 202046 528838 202102
rect 528894 202046 528962 202102
rect 529018 202046 529088 202102
rect 528768 201978 529088 202046
rect 528768 201922 528838 201978
rect 528894 201922 528962 201978
rect 529018 201922 529088 201978
rect 528768 201888 529088 201922
rect 559488 202350 559808 202384
rect 559488 202294 559558 202350
rect 559614 202294 559682 202350
rect 559738 202294 559808 202350
rect 559488 202226 559808 202294
rect 559488 202170 559558 202226
rect 559614 202170 559682 202226
rect 559738 202170 559808 202226
rect 559488 202102 559808 202170
rect 559488 202046 559558 202102
rect 559614 202046 559682 202102
rect 559738 202046 559808 202102
rect 559488 201978 559808 202046
rect 559488 201922 559558 201978
rect 559614 201922 559682 201978
rect 559738 201922 559808 201978
rect 559488 201888 559808 201922
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 359808 190350 360128 190384
rect 359808 190294 359878 190350
rect 359934 190294 360002 190350
rect 360058 190294 360128 190350
rect 359808 190226 360128 190294
rect 359808 190170 359878 190226
rect 359934 190170 360002 190226
rect 360058 190170 360128 190226
rect 359808 190102 360128 190170
rect 359808 190046 359878 190102
rect 359934 190046 360002 190102
rect 360058 190046 360128 190102
rect 359808 189978 360128 190046
rect 359808 189922 359878 189978
rect 359934 189922 360002 189978
rect 360058 189922 360128 189978
rect 359808 189888 360128 189922
rect 390528 190350 390848 190384
rect 390528 190294 390598 190350
rect 390654 190294 390722 190350
rect 390778 190294 390848 190350
rect 390528 190226 390848 190294
rect 390528 190170 390598 190226
rect 390654 190170 390722 190226
rect 390778 190170 390848 190226
rect 390528 190102 390848 190170
rect 390528 190046 390598 190102
rect 390654 190046 390722 190102
rect 390778 190046 390848 190102
rect 390528 189978 390848 190046
rect 390528 189922 390598 189978
rect 390654 189922 390722 189978
rect 390778 189922 390848 189978
rect 390528 189888 390848 189922
rect 421248 190350 421568 190384
rect 421248 190294 421318 190350
rect 421374 190294 421442 190350
rect 421498 190294 421568 190350
rect 421248 190226 421568 190294
rect 421248 190170 421318 190226
rect 421374 190170 421442 190226
rect 421498 190170 421568 190226
rect 421248 190102 421568 190170
rect 421248 190046 421318 190102
rect 421374 190046 421442 190102
rect 421498 190046 421568 190102
rect 421248 189978 421568 190046
rect 421248 189922 421318 189978
rect 421374 189922 421442 189978
rect 421498 189922 421568 189978
rect 421248 189888 421568 189922
rect 451968 190350 452288 190384
rect 451968 190294 452038 190350
rect 452094 190294 452162 190350
rect 452218 190294 452288 190350
rect 451968 190226 452288 190294
rect 451968 190170 452038 190226
rect 452094 190170 452162 190226
rect 452218 190170 452288 190226
rect 451968 190102 452288 190170
rect 451968 190046 452038 190102
rect 452094 190046 452162 190102
rect 452218 190046 452288 190102
rect 451968 189978 452288 190046
rect 451968 189922 452038 189978
rect 452094 189922 452162 189978
rect 452218 189922 452288 189978
rect 451968 189888 452288 189922
rect 482688 190350 483008 190384
rect 482688 190294 482758 190350
rect 482814 190294 482882 190350
rect 482938 190294 483008 190350
rect 482688 190226 483008 190294
rect 482688 190170 482758 190226
rect 482814 190170 482882 190226
rect 482938 190170 483008 190226
rect 482688 190102 483008 190170
rect 482688 190046 482758 190102
rect 482814 190046 482882 190102
rect 482938 190046 483008 190102
rect 482688 189978 483008 190046
rect 482688 189922 482758 189978
rect 482814 189922 482882 189978
rect 482938 189922 483008 189978
rect 482688 189888 483008 189922
rect 513408 190350 513728 190384
rect 513408 190294 513478 190350
rect 513534 190294 513602 190350
rect 513658 190294 513728 190350
rect 513408 190226 513728 190294
rect 513408 190170 513478 190226
rect 513534 190170 513602 190226
rect 513658 190170 513728 190226
rect 513408 190102 513728 190170
rect 513408 190046 513478 190102
rect 513534 190046 513602 190102
rect 513658 190046 513728 190102
rect 513408 189978 513728 190046
rect 513408 189922 513478 189978
rect 513534 189922 513602 189978
rect 513658 189922 513728 189978
rect 513408 189888 513728 189922
rect 544128 190350 544448 190384
rect 544128 190294 544198 190350
rect 544254 190294 544322 190350
rect 544378 190294 544448 190350
rect 544128 190226 544448 190294
rect 544128 190170 544198 190226
rect 544254 190170 544322 190226
rect 544378 190170 544448 190226
rect 544128 190102 544448 190170
rect 544128 190046 544198 190102
rect 544254 190046 544322 190102
rect 544378 190046 544448 190102
rect 544128 189978 544448 190046
rect 544128 189922 544198 189978
rect 544254 189922 544322 189978
rect 544378 189922 544448 189978
rect 544128 189888 544448 189922
rect 574848 190350 575168 190384
rect 574848 190294 574918 190350
rect 574974 190294 575042 190350
rect 575098 190294 575168 190350
rect 574848 190226 575168 190294
rect 574848 190170 574918 190226
rect 574974 190170 575042 190226
rect 575098 190170 575168 190226
rect 574848 190102 575168 190170
rect 574848 190046 574918 190102
rect 574974 190046 575042 190102
rect 575098 190046 575168 190102
rect 574848 189978 575168 190046
rect 574848 189922 574918 189978
rect 574974 189922 575042 189978
rect 575098 189922 575168 189978
rect 574848 189888 575168 189922
rect 344448 184350 344768 184384
rect 344448 184294 344518 184350
rect 344574 184294 344642 184350
rect 344698 184294 344768 184350
rect 344448 184226 344768 184294
rect 344448 184170 344518 184226
rect 344574 184170 344642 184226
rect 344698 184170 344768 184226
rect 344448 184102 344768 184170
rect 344448 184046 344518 184102
rect 344574 184046 344642 184102
rect 344698 184046 344768 184102
rect 344448 183978 344768 184046
rect 344448 183922 344518 183978
rect 344574 183922 344642 183978
rect 344698 183922 344768 183978
rect 344448 183888 344768 183922
rect 375168 184350 375488 184384
rect 375168 184294 375238 184350
rect 375294 184294 375362 184350
rect 375418 184294 375488 184350
rect 375168 184226 375488 184294
rect 375168 184170 375238 184226
rect 375294 184170 375362 184226
rect 375418 184170 375488 184226
rect 375168 184102 375488 184170
rect 375168 184046 375238 184102
rect 375294 184046 375362 184102
rect 375418 184046 375488 184102
rect 375168 183978 375488 184046
rect 375168 183922 375238 183978
rect 375294 183922 375362 183978
rect 375418 183922 375488 183978
rect 375168 183888 375488 183922
rect 405888 184350 406208 184384
rect 405888 184294 405958 184350
rect 406014 184294 406082 184350
rect 406138 184294 406208 184350
rect 405888 184226 406208 184294
rect 405888 184170 405958 184226
rect 406014 184170 406082 184226
rect 406138 184170 406208 184226
rect 405888 184102 406208 184170
rect 405888 184046 405958 184102
rect 406014 184046 406082 184102
rect 406138 184046 406208 184102
rect 405888 183978 406208 184046
rect 405888 183922 405958 183978
rect 406014 183922 406082 183978
rect 406138 183922 406208 183978
rect 405888 183888 406208 183922
rect 436608 184350 436928 184384
rect 436608 184294 436678 184350
rect 436734 184294 436802 184350
rect 436858 184294 436928 184350
rect 436608 184226 436928 184294
rect 436608 184170 436678 184226
rect 436734 184170 436802 184226
rect 436858 184170 436928 184226
rect 436608 184102 436928 184170
rect 436608 184046 436678 184102
rect 436734 184046 436802 184102
rect 436858 184046 436928 184102
rect 436608 183978 436928 184046
rect 436608 183922 436678 183978
rect 436734 183922 436802 183978
rect 436858 183922 436928 183978
rect 436608 183888 436928 183922
rect 467328 184350 467648 184384
rect 467328 184294 467398 184350
rect 467454 184294 467522 184350
rect 467578 184294 467648 184350
rect 467328 184226 467648 184294
rect 467328 184170 467398 184226
rect 467454 184170 467522 184226
rect 467578 184170 467648 184226
rect 467328 184102 467648 184170
rect 467328 184046 467398 184102
rect 467454 184046 467522 184102
rect 467578 184046 467648 184102
rect 467328 183978 467648 184046
rect 467328 183922 467398 183978
rect 467454 183922 467522 183978
rect 467578 183922 467648 183978
rect 467328 183888 467648 183922
rect 498048 184350 498368 184384
rect 498048 184294 498118 184350
rect 498174 184294 498242 184350
rect 498298 184294 498368 184350
rect 498048 184226 498368 184294
rect 498048 184170 498118 184226
rect 498174 184170 498242 184226
rect 498298 184170 498368 184226
rect 498048 184102 498368 184170
rect 498048 184046 498118 184102
rect 498174 184046 498242 184102
rect 498298 184046 498368 184102
rect 498048 183978 498368 184046
rect 498048 183922 498118 183978
rect 498174 183922 498242 183978
rect 498298 183922 498368 183978
rect 498048 183888 498368 183922
rect 528768 184350 529088 184384
rect 528768 184294 528838 184350
rect 528894 184294 528962 184350
rect 529018 184294 529088 184350
rect 528768 184226 529088 184294
rect 528768 184170 528838 184226
rect 528894 184170 528962 184226
rect 529018 184170 529088 184226
rect 528768 184102 529088 184170
rect 528768 184046 528838 184102
rect 528894 184046 528962 184102
rect 529018 184046 529088 184102
rect 528768 183978 529088 184046
rect 528768 183922 528838 183978
rect 528894 183922 528962 183978
rect 529018 183922 529088 183978
rect 528768 183888 529088 183922
rect 559488 184350 559808 184384
rect 559488 184294 559558 184350
rect 559614 184294 559682 184350
rect 559738 184294 559808 184350
rect 559488 184226 559808 184294
rect 559488 184170 559558 184226
rect 559614 184170 559682 184226
rect 559738 184170 559808 184226
rect 559488 184102 559808 184170
rect 559488 184046 559558 184102
rect 559614 184046 559682 184102
rect 559738 184046 559808 184102
rect 559488 183978 559808 184046
rect 559488 183922 559558 183978
rect 559614 183922 559682 183978
rect 559738 183922 559808 183978
rect 559488 183888 559808 183922
rect 589098 184350 589718 201922
rect 590492 390404 590548 390414
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 341404 173098 341460 173108
rect 341292 168058 341348 168068
rect 341180 162298 341236 162308
rect 341180 155316 341236 162242
rect 341180 155250 341236 155260
rect 341292 145236 341348 168002
rect 341404 147812 341460 173042
rect 359808 172350 360128 172384
rect 359808 172294 359878 172350
rect 359934 172294 360002 172350
rect 360058 172294 360128 172350
rect 359808 172226 360128 172294
rect 359808 172170 359878 172226
rect 359934 172170 360002 172226
rect 360058 172170 360128 172226
rect 359808 172102 360128 172170
rect 359808 172046 359878 172102
rect 359934 172046 360002 172102
rect 360058 172046 360128 172102
rect 359808 171978 360128 172046
rect 359808 171922 359878 171978
rect 359934 171922 360002 171978
rect 360058 171922 360128 171978
rect 359808 171888 360128 171922
rect 390528 172350 390848 172384
rect 390528 172294 390598 172350
rect 390654 172294 390722 172350
rect 390778 172294 390848 172350
rect 390528 172226 390848 172294
rect 390528 172170 390598 172226
rect 390654 172170 390722 172226
rect 390778 172170 390848 172226
rect 390528 172102 390848 172170
rect 390528 172046 390598 172102
rect 390654 172046 390722 172102
rect 390778 172046 390848 172102
rect 390528 171978 390848 172046
rect 390528 171922 390598 171978
rect 390654 171922 390722 171978
rect 390778 171922 390848 171978
rect 390528 171888 390848 171922
rect 421248 172350 421568 172384
rect 421248 172294 421318 172350
rect 421374 172294 421442 172350
rect 421498 172294 421568 172350
rect 421248 172226 421568 172294
rect 421248 172170 421318 172226
rect 421374 172170 421442 172226
rect 421498 172170 421568 172226
rect 421248 172102 421568 172170
rect 421248 172046 421318 172102
rect 421374 172046 421442 172102
rect 421498 172046 421568 172102
rect 421248 171978 421568 172046
rect 421248 171922 421318 171978
rect 421374 171922 421442 171978
rect 421498 171922 421568 171978
rect 421248 171888 421568 171922
rect 451968 172350 452288 172384
rect 451968 172294 452038 172350
rect 452094 172294 452162 172350
rect 452218 172294 452288 172350
rect 451968 172226 452288 172294
rect 451968 172170 452038 172226
rect 452094 172170 452162 172226
rect 452218 172170 452288 172226
rect 451968 172102 452288 172170
rect 451968 172046 452038 172102
rect 452094 172046 452162 172102
rect 452218 172046 452288 172102
rect 451968 171978 452288 172046
rect 451968 171922 452038 171978
rect 452094 171922 452162 171978
rect 452218 171922 452288 171978
rect 451968 171888 452288 171922
rect 482688 172350 483008 172384
rect 482688 172294 482758 172350
rect 482814 172294 482882 172350
rect 482938 172294 483008 172350
rect 482688 172226 483008 172294
rect 482688 172170 482758 172226
rect 482814 172170 482882 172226
rect 482938 172170 483008 172226
rect 482688 172102 483008 172170
rect 482688 172046 482758 172102
rect 482814 172046 482882 172102
rect 482938 172046 483008 172102
rect 482688 171978 483008 172046
rect 482688 171922 482758 171978
rect 482814 171922 482882 171978
rect 482938 171922 483008 171978
rect 482688 171888 483008 171922
rect 513408 172350 513728 172384
rect 513408 172294 513478 172350
rect 513534 172294 513602 172350
rect 513658 172294 513728 172350
rect 513408 172226 513728 172294
rect 513408 172170 513478 172226
rect 513534 172170 513602 172226
rect 513658 172170 513728 172226
rect 513408 172102 513728 172170
rect 513408 172046 513478 172102
rect 513534 172046 513602 172102
rect 513658 172046 513728 172102
rect 513408 171978 513728 172046
rect 513408 171922 513478 171978
rect 513534 171922 513602 171978
rect 513658 171922 513728 171978
rect 513408 171888 513728 171922
rect 544128 172350 544448 172384
rect 544128 172294 544198 172350
rect 544254 172294 544322 172350
rect 544378 172294 544448 172350
rect 544128 172226 544448 172294
rect 544128 172170 544198 172226
rect 544254 172170 544322 172226
rect 544378 172170 544448 172226
rect 544128 172102 544448 172170
rect 544128 172046 544198 172102
rect 544254 172046 544322 172102
rect 544378 172046 544448 172102
rect 544128 171978 544448 172046
rect 544128 171922 544198 171978
rect 544254 171922 544322 171978
rect 544378 171922 544448 171978
rect 544128 171888 544448 171922
rect 574848 172350 575168 172384
rect 574848 172294 574918 172350
rect 574974 172294 575042 172350
rect 575098 172294 575168 172350
rect 574848 172226 575168 172294
rect 574848 172170 574918 172226
rect 574974 172170 575042 172226
rect 575098 172170 575168 172226
rect 574848 172102 575168 172170
rect 574848 172046 574918 172102
rect 574974 172046 575042 172102
rect 575098 172046 575168 172102
rect 574848 171978 575168 172046
rect 574848 171922 574918 171978
rect 574974 171922 575042 171978
rect 575098 171922 575168 171978
rect 574848 171888 575168 171922
rect 344448 166350 344768 166384
rect 344448 166294 344518 166350
rect 344574 166294 344642 166350
rect 344698 166294 344768 166350
rect 344448 166226 344768 166294
rect 344448 166170 344518 166226
rect 344574 166170 344642 166226
rect 344698 166170 344768 166226
rect 344448 166102 344768 166170
rect 344448 166046 344518 166102
rect 344574 166046 344642 166102
rect 344698 166046 344768 166102
rect 344448 165978 344768 166046
rect 344448 165922 344518 165978
rect 344574 165922 344642 165978
rect 344698 165922 344768 165978
rect 344448 165888 344768 165922
rect 375168 166350 375488 166384
rect 375168 166294 375238 166350
rect 375294 166294 375362 166350
rect 375418 166294 375488 166350
rect 375168 166226 375488 166294
rect 375168 166170 375238 166226
rect 375294 166170 375362 166226
rect 375418 166170 375488 166226
rect 375168 166102 375488 166170
rect 375168 166046 375238 166102
rect 375294 166046 375362 166102
rect 375418 166046 375488 166102
rect 375168 165978 375488 166046
rect 375168 165922 375238 165978
rect 375294 165922 375362 165978
rect 375418 165922 375488 165978
rect 375168 165888 375488 165922
rect 405888 166350 406208 166384
rect 405888 166294 405958 166350
rect 406014 166294 406082 166350
rect 406138 166294 406208 166350
rect 405888 166226 406208 166294
rect 405888 166170 405958 166226
rect 406014 166170 406082 166226
rect 406138 166170 406208 166226
rect 405888 166102 406208 166170
rect 405888 166046 405958 166102
rect 406014 166046 406082 166102
rect 406138 166046 406208 166102
rect 405888 165978 406208 166046
rect 405888 165922 405958 165978
rect 406014 165922 406082 165978
rect 406138 165922 406208 165978
rect 405888 165888 406208 165922
rect 436608 166350 436928 166384
rect 436608 166294 436678 166350
rect 436734 166294 436802 166350
rect 436858 166294 436928 166350
rect 436608 166226 436928 166294
rect 436608 166170 436678 166226
rect 436734 166170 436802 166226
rect 436858 166170 436928 166226
rect 436608 166102 436928 166170
rect 436608 166046 436678 166102
rect 436734 166046 436802 166102
rect 436858 166046 436928 166102
rect 436608 165978 436928 166046
rect 436608 165922 436678 165978
rect 436734 165922 436802 165978
rect 436858 165922 436928 165978
rect 436608 165888 436928 165922
rect 467328 166350 467648 166384
rect 467328 166294 467398 166350
rect 467454 166294 467522 166350
rect 467578 166294 467648 166350
rect 467328 166226 467648 166294
rect 467328 166170 467398 166226
rect 467454 166170 467522 166226
rect 467578 166170 467648 166226
rect 467328 166102 467648 166170
rect 467328 166046 467398 166102
rect 467454 166046 467522 166102
rect 467578 166046 467648 166102
rect 467328 165978 467648 166046
rect 467328 165922 467398 165978
rect 467454 165922 467522 165978
rect 467578 165922 467648 165978
rect 467328 165888 467648 165922
rect 498048 166350 498368 166384
rect 498048 166294 498118 166350
rect 498174 166294 498242 166350
rect 498298 166294 498368 166350
rect 498048 166226 498368 166294
rect 498048 166170 498118 166226
rect 498174 166170 498242 166226
rect 498298 166170 498368 166226
rect 498048 166102 498368 166170
rect 498048 166046 498118 166102
rect 498174 166046 498242 166102
rect 498298 166046 498368 166102
rect 498048 165978 498368 166046
rect 498048 165922 498118 165978
rect 498174 165922 498242 165978
rect 498298 165922 498368 165978
rect 498048 165888 498368 165922
rect 528768 166350 529088 166384
rect 528768 166294 528838 166350
rect 528894 166294 528962 166350
rect 529018 166294 529088 166350
rect 528768 166226 529088 166294
rect 528768 166170 528838 166226
rect 528894 166170 528962 166226
rect 529018 166170 529088 166226
rect 528768 166102 529088 166170
rect 528768 166046 528838 166102
rect 528894 166046 528962 166102
rect 529018 166046 529088 166102
rect 528768 165978 529088 166046
rect 528768 165922 528838 165978
rect 528894 165922 528962 165978
rect 529018 165922 529088 165978
rect 528768 165888 529088 165922
rect 559488 166350 559808 166384
rect 559488 166294 559558 166350
rect 559614 166294 559682 166350
rect 559738 166294 559808 166350
rect 559488 166226 559808 166294
rect 559488 166170 559558 166226
rect 559614 166170 559682 166226
rect 559738 166170 559808 166226
rect 559488 166102 559808 166170
rect 559488 166046 559558 166102
rect 559614 166046 559682 166102
rect 559738 166046 559808 166102
rect 559488 165978 559808 166046
rect 559488 165922 559558 165978
rect 559614 165922 559682 165978
rect 559738 165922 559808 165978
rect 559488 165888 559808 165922
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 341516 162118 341572 162128
rect 341516 158900 341572 162062
rect 422604 161140 422660 161150
rect 422604 160020 422660 161084
rect 422604 159954 422660 159964
rect 422828 161028 422884 161038
rect 422828 160020 422884 160972
rect 422828 159954 422884 159964
rect 467852 160916 467908 160926
rect 467852 160020 467908 160860
rect 467852 159954 467908 159964
rect 357868 159598 357924 159608
rect 341516 158834 341572 158844
rect 341404 147746 341460 147756
rect 341516 155316 341572 155326
rect 341292 145170 341348 145180
rect 340956 138472 341012 138482
rect 341516 131012 341572 155260
rect 341516 130946 341572 130956
rect 343338 148350 343958 159418
rect 343338 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 343958 148350
rect 343338 148226 343958 148294
rect 343338 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 343958 148226
rect 343338 148102 343958 148170
rect 343338 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 343958 148102
rect 343338 147978 343958 148046
rect 343338 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 343958 147978
rect 340396 21410 340452 21420
rect 343338 130350 343958 147922
rect 343338 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 343958 130350
rect 343338 130226 343958 130294
rect 343338 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 343958 130226
rect 343338 130102 343958 130170
rect 343338 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 343958 130102
rect 343338 129978 343958 130046
rect 343338 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 343958 129978
rect 343338 112350 343958 129922
rect 343338 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 343958 112350
rect 343338 112226 343958 112294
rect 343338 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 343958 112226
rect 343338 112102 343958 112170
rect 343338 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 343958 112102
rect 343338 111978 343958 112046
rect 343338 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 343958 111978
rect 343338 94350 343958 111922
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 343338 76350 343958 93922
rect 343338 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 343958 76350
rect 343338 76226 343958 76294
rect 343338 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 343958 76226
rect 343338 76102 343958 76170
rect 343338 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 343958 76102
rect 343338 75978 343958 76046
rect 343338 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 343958 75978
rect 343338 58350 343958 75922
rect 343338 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 343958 58350
rect 343338 58226 343958 58294
rect 343338 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 343958 58226
rect 343338 58102 343958 58170
rect 343338 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 343958 58102
rect 343338 57978 343958 58046
rect 343338 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 343958 57978
rect 343338 40350 343958 57922
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 343338 22350 343958 39922
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 327516 20066 327572 20076
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 316338 -1120 316958 9922
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 4350 343958 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 154350 347678 159418
rect 357868 159236 357924 159542
rect 357868 159170 357924 159180
rect 347058 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 347678 154350
rect 347058 154226 347678 154294
rect 347058 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 347678 154226
rect 347058 154102 347678 154170
rect 347058 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 347678 154102
rect 347058 153978 347678 154046
rect 347058 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 347678 153978
rect 347058 136350 347678 153922
rect 347058 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 347678 136350
rect 347058 136226 347678 136294
rect 347058 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 347678 136226
rect 347058 136102 347678 136170
rect 347058 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 347678 136102
rect 347058 135978 347678 136046
rect 347058 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 347678 135978
rect 347058 118350 347678 135922
rect 374058 148350 374678 159418
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 347058 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 347678 118350
rect 347058 118226 347678 118294
rect 347058 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 347678 118226
rect 347058 118102 347678 118170
rect 347058 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 347678 118102
rect 347058 117978 347678 118046
rect 347058 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 347678 117978
rect 347058 100350 347678 117922
rect 347058 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 347678 100350
rect 347058 100226 347678 100294
rect 347058 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 347678 100226
rect 347058 100102 347678 100170
rect 347058 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 347678 100102
rect 347058 99978 347678 100046
rect 347058 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 347678 99978
rect 347058 82350 347678 99922
rect 367052 135478 367108 135488
rect 366268 94052 366324 94062
rect 366268 91588 366324 93996
rect 367052 94052 367108 135422
rect 374058 130350 374678 147922
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 374058 112350 374678 129922
rect 374058 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 374678 112350
rect 374058 112226 374678 112294
rect 374058 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 374678 112226
rect 374058 112102 374678 112170
rect 374058 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 374678 112102
rect 374058 111978 374678 112046
rect 374058 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 374678 111978
rect 374058 98428 374678 111922
rect 377778 154350 378398 159418
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 377778 136350 378398 153922
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 377778 118350 378398 135922
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 377778 100350 378398 117922
rect 404778 148350 405398 159418
rect 404778 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 405398 148350
rect 404778 148226 405398 148294
rect 404778 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 405398 148226
rect 404778 148102 405398 148170
rect 404778 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 405398 148102
rect 404778 147978 405398 148046
rect 404778 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 405398 147978
rect 404778 130350 405398 147922
rect 404778 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 405398 130350
rect 404778 130226 405398 130294
rect 404778 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 405398 130226
rect 404778 130102 405398 130170
rect 404778 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 405398 130102
rect 404778 129978 405398 130046
rect 404778 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 405398 129978
rect 404778 112350 405398 129922
rect 404778 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 405398 112350
rect 404778 112226 405398 112294
rect 404778 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 405398 112226
rect 404778 112102 405398 112170
rect 404778 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 405398 112102
rect 404778 111978 405398 112046
rect 404778 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 405398 111978
rect 403228 103978 403284 103988
rect 403228 103908 403284 103922
rect 403228 103842 403284 103852
rect 377778 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 378398 100350
rect 377778 100226 378398 100294
rect 377778 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 378398 100226
rect 377778 100102 378398 100170
rect 377778 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 378398 100102
rect 377778 99978 378398 100046
rect 377778 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 378398 99978
rect 377778 97622 378398 99922
rect 404778 98428 405398 111922
rect 408498 154350 409118 159418
rect 408498 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 409118 154350
rect 408498 154226 409118 154294
rect 408498 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 409118 154226
rect 408498 154102 409118 154170
rect 408498 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 409118 154102
rect 408498 153978 409118 154046
rect 408498 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 409118 153978
rect 408498 136350 409118 153922
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408498 118350 409118 135922
rect 435498 148350 436118 159418
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 423276 122724 423332 122734
rect 423276 122518 423332 122668
rect 423276 122452 423332 122462
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 406700 104158 406756 104168
rect 406700 104020 406756 104102
rect 406700 103954 406756 103964
rect 408498 100350 409118 117922
rect 413308 115318 413364 115328
rect 413308 104132 413364 115262
rect 413308 104066 413364 104076
rect 414988 115138 415044 115148
rect 414988 104132 415044 115082
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 414988 104066 415044 104076
rect 421820 107044 421876 107054
rect 408498 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 409118 100350
rect 408498 100226 409118 100294
rect 408498 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 409118 100226
rect 408498 100102 409118 100170
rect 408498 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 409118 100102
rect 408498 99978 409118 100046
rect 408498 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 409118 99978
rect 408498 97622 409118 99922
rect 421708 100212 421764 100222
rect 367052 93986 367108 93996
rect 374448 94350 374768 94384
rect 374448 94294 374518 94350
rect 374574 94294 374642 94350
rect 374698 94294 374768 94350
rect 374448 94226 374768 94294
rect 374448 94170 374518 94226
rect 374574 94170 374642 94226
rect 374698 94170 374768 94226
rect 374448 94102 374768 94170
rect 374448 94046 374518 94102
rect 374574 94046 374642 94102
rect 374698 94046 374768 94102
rect 374448 93978 374768 94046
rect 374448 93922 374518 93978
rect 374574 93922 374642 93978
rect 374698 93922 374768 93978
rect 374448 93888 374768 93922
rect 405168 94350 405488 94384
rect 405168 94294 405238 94350
rect 405294 94294 405362 94350
rect 405418 94294 405488 94350
rect 405168 94226 405488 94294
rect 405168 94170 405238 94226
rect 405294 94170 405362 94226
rect 405418 94170 405488 94226
rect 405168 94102 405488 94170
rect 405168 94046 405238 94102
rect 405294 94046 405362 94102
rect 405418 94046 405488 94102
rect 405168 93978 405488 94046
rect 405168 93922 405238 93978
rect 405294 93922 405362 93978
rect 405418 93922 405488 93978
rect 405168 93888 405488 93922
rect 366268 91522 366324 91532
rect 421708 91588 421764 100156
rect 421820 97076 421876 106988
rect 421820 97010 421876 97020
rect 424172 97076 424228 97086
rect 421708 91522 421764 91532
rect 347058 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 347678 82350
rect 347058 82226 347678 82294
rect 347058 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 347678 82226
rect 347058 82102 347678 82170
rect 347058 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 347678 82102
rect 347058 81978 347678 82046
rect 347058 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 347678 81978
rect 347058 64350 347678 81922
rect 389808 82350 390128 82384
rect 389808 82294 389878 82350
rect 389934 82294 390002 82350
rect 390058 82294 390128 82350
rect 389808 82226 390128 82294
rect 389808 82170 389878 82226
rect 389934 82170 390002 82226
rect 390058 82170 390128 82226
rect 389808 82102 390128 82170
rect 389808 82046 389878 82102
rect 389934 82046 390002 82102
rect 390058 82046 390128 82102
rect 389808 81978 390128 82046
rect 389808 81922 389878 81978
rect 389934 81922 390002 81978
rect 390058 81922 390128 81978
rect 389808 81888 390128 81922
rect 374448 76350 374768 76384
rect 374448 76294 374518 76350
rect 374574 76294 374642 76350
rect 374698 76294 374768 76350
rect 374448 76226 374768 76294
rect 374448 76170 374518 76226
rect 374574 76170 374642 76226
rect 374698 76170 374768 76226
rect 374448 76102 374768 76170
rect 374448 76046 374518 76102
rect 374574 76046 374642 76102
rect 374698 76046 374768 76102
rect 374448 75978 374768 76046
rect 374448 75922 374518 75978
rect 374574 75922 374642 75978
rect 374698 75922 374768 75978
rect 374448 75888 374768 75922
rect 405168 76350 405488 76384
rect 405168 76294 405238 76350
rect 405294 76294 405362 76350
rect 405418 76294 405488 76350
rect 405168 76226 405488 76294
rect 405168 76170 405238 76226
rect 405294 76170 405362 76226
rect 405418 76170 405488 76226
rect 405168 76102 405488 76170
rect 405168 76046 405238 76102
rect 405294 76046 405362 76102
rect 405418 76046 405488 76102
rect 405168 75978 405488 76046
rect 405168 75922 405238 75978
rect 405294 75922 405362 75978
rect 405418 75922 405488 75978
rect 405168 75888 405488 75922
rect 347058 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 347678 64350
rect 347058 64226 347678 64294
rect 347058 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 347678 64226
rect 347058 64102 347678 64170
rect 347058 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 347678 64102
rect 347058 63978 347678 64046
rect 347058 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 347678 63978
rect 347058 46350 347678 63922
rect 389808 64350 390128 64384
rect 389808 64294 389878 64350
rect 389934 64294 390002 64350
rect 390058 64294 390128 64350
rect 389808 64226 390128 64294
rect 389808 64170 389878 64226
rect 389934 64170 390002 64226
rect 390058 64170 390128 64226
rect 389808 64102 390128 64170
rect 389808 64046 389878 64102
rect 389934 64046 390002 64102
rect 390058 64046 390128 64102
rect 389808 63978 390128 64046
rect 389808 63922 389878 63978
rect 389934 63922 390002 63978
rect 390058 63922 390128 63978
rect 389808 63888 390128 63922
rect 374448 58350 374768 58384
rect 374448 58294 374518 58350
rect 374574 58294 374642 58350
rect 374698 58294 374768 58350
rect 374448 58226 374768 58294
rect 374448 58170 374518 58226
rect 374574 58170 374642 58226
rect 374698 58170 374768 58226
rect 374448 58102 374768 58170
rect 374448 58046 374518 58102
rect 374574 58046 374642 58102
rect 374698 58046 374768 58102
rect 374448 57978 374768 58046
rect 374448 57922 374518 57978
rect 374574 57922 374642 57978
rect 374698 57922 374768 57978
rect 374448 57888 374768 57922
rect 405168 58350 405488 58384
rect 405168 58294 405238 58350
rect 405294 58294 405362 58350
rect 405418 58294 405488 58350
rect 405168 58226 405488 58294
rect 405168 58170 405238 58226
rect 405294 58170 405362 58226
rect 405418 58170 405488 58226
rect 405168 58102 405488 58170
rect 405168 58046 405238 58102
rect 405294 58046 405362 58102
rect 405418 58046 405488 58102
rect 405168 57978 405488 58046
rect 405168 57922 405238 57978
rect 405294 57922 405362 57978
rect 405418 57922 405488 57978
rect 405168 57888 405488 57922
rect 347058 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 347678 46350
rect 347058 46226 347678 46294
rect 347058 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 347678 46226
rect 347058 46102 347678 46170
rect 347058 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 347678 46102
rect 347058 45978 347678 46046
rect 347058 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 347678 45978
rect 347058 28350 347678 45922
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 347058 10350 347678 27922
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 347058 -1120 347678 9922
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 40350 374678 50964
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 374058 22350 374678 39922
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 374058 4350 374678 21922
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 46350 378398 51210
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 377778 -1120 378398 9922
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 40350 405398 50964
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 404778 22350 405398 39922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 408498 46350 409118 51210
rect 408498 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 409118 46350
rect 408498 46226 409118 46294
rect 408498 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 409118 46226
rect 408498 46102 409118 46170
rect 408498 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 409118 46102
rect 408498 45978 409118 46046
rect 408498 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 409118 45978
rect 408498 28350 409118 45922
rect 424172 37828 424228 97020
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 424172 37762 424228 37772
rect 427532 91588 427588 91598
rect 427532 31332 427588 91532
rect 427532 31266 427588 31276
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 408498 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 409118 28350
rect 408498 28226 409118 28294
rect 408498 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 409118 28226
rect 408498 28102 409118 28170
rect 408498 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 409118 28102
rect 408498 27978 409118 28046
rect 408498 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 409118 27978
rect 408498 10350 409118 27922
rect 408498 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 409118 10350
rect 408498 10226 409118 10294
rect 408498 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 409118 10226
rect 408498 10102 409118 10170
rect 408498 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 409118 10102
rect 408498 9978 409118 10046
rect 408498 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 409118 9978
rect 408498 -1120 409118 9922
rect 408498 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 409118 -1120
rect 408498 -1244 409118 -1176
rect 408498 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 409118 -1244
rect 408498 -1368 409118 -1300
rect 408498 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 409118 -1368
rect 408498 -1492 409118 -1424
rect 408498 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 409118 -1492
rect 408498 -1644 409118 -1548
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 154350 439838 159418
rect 576268 158698 576324 158708
rect 558460 157668 558516 157678
rect 514108 157556 514164 157566
rect 558460 157552 558516 157562
rect 514108 157438 514164 157500
rect 514108 157372 514164 157382
rect 574812 155638 574868 155648
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 574028 155428 574084 155438
rect 462924 149716 462980 149726
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 457996 149698 458052 149708
rect 457996 136052 458052 149642
rect 457996 135986 458052 135996
rect 462812 146244 462868 146254
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 462812 132418 462868 146188
rect 462924 137458 462980 149660
rect 463708 148148 463764 148158
rect 463148 144658 463204 144668
rect 462924 137392 462980 137402
rect 463036 141428 463092 141438
rect 463036 132598 463092 141372
rect 463148 135658 463204 144602
rect 463708 142660 463764 148092
rect 463708 142594 463764 142604
rect 466396 146356 466452 146366
rect 466284 141316 466340 141326
rect 463148 135592 463204 135602
rect 463260 141238 463316 141248
rect 463260 134398 463316 141182
rect 465388 139798 465444 139808
rect 465388 135298 465444 139742
rect 466172 139636 466228 139646
rect 465388 135232 465444 135242
rect 465500 139618 465556 139628
rect 463260 134332 463316 134342
rect 463036 132532 463092 132542
rect 462812 132352 462868 132362
rect 465500 132238 465556 139562
rect 465500 132172 465556 132182
rect 464448 130350 464768 130384
rect 464448 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 464768 130350
rect 464448 130226 464768 130294
rect 464448 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 464768 130226
rect 464448 130102 464768 130170
rect 464448 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 464768 130102
rect 464448 129978 464768 130046
rect 464448 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 464768 129978
rect 464448 129888 464768 129922
rect 466172 122518 466228 139580
rect 466284 127558 466340 141260
rect 466396 135478 466452 146300
rect 466732 144838 466788 144848
rect 466396 135412 466452 135422
rect 466620 141204 466676 141214
rect 466620 134038 466676 141148
rect 466732 137638 466788 144782
rect 490028 144838 490084 144848
rect 472892 143220 472948 143230
rect 468636 143108 468692 143118
rect 468636 142498 468692 143052
rect 472892 142678 472948 143164
rect 490028 142884 490084 144782
rect 490028 142818 490084 142828
rect 497868 144658 497924 144668
rect 497868 142884 497924 144602
rect 497868 142818 497924 142828
rect 505708 144478 505764 144488
rect 505708 142884 505764 144422
rect 520156 144004 520212 144014
rect 513548 143938 513604 143948
rect 505708 142818 505764 142828
rect 507276 143758 507332 143768
rect 507276 142884 507332 143702
rect 507276 142818 507332 142828
rect 508844 143578 508900 143588
rect 508844 142884 508900 143522
rect 508844 142818 508900 142828
rect 511980 142884 512036 142896
rect 513548 142884 513604 143882
rect 520156 143668 520212 143948
rect 520156 143602 520212 143612
rect 513548 142818 513604 142828
rect 511980 142792 512036 142802
rect 472892 142612 472948 142622
rect 468636 142432 468692 142442
rect 479612 141764 479668 141774
rect 479612 141316 479668 141708
rect 479612 141250 479668 141260
rect 480620 139798 480676 139808
rect 480620 139682 480676 139692
rect 482188 139636 482244 139646
rect 482188 139542 482244 139562
rect 466732 137572 466788 137582
rect 467068 139524 467124 139534
rect 467068 134218 467124 139468
rect 501676 139524 501732 139534
rect 501676 138516 501732 139468
rect 501676 138450 501732 138460
rect 574028 137788 574084 155372
rect 574476 153076 574532 153086
rect 574252 138538 574308 138548
rect 574028 137732 574196 137788
rect 479808 136350 480128 136384
rect 479808 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 480128 136350
rect 479808 136226 480128 136294
rect 479808 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 480128 136226
rect 479808 136102 480128 136170
rect 479808 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 480128 136102
rect 479808 135978 480128 136046
rect 479808 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 480128 135978
rect 479808 135888 480128 135922
rect 510528 136350 510848 136384
rect 510528 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 510848 136350
rect 510528 136226 510848 136294
rect 510528 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 510848 136226
rect 510528 136102 510848 136170
rect 510528 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 510848 136102
rect 510528 135978 510848 136046
rect 510528 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 510848 135978
rect 510528 135888 510848 135922
rect 541248 136350 541568 136384
rect 541248 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 541568 136350
rect 541248 136226 541568 136294
rect 541248 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 541568 136226
rect 541248 136102 541568 136170
rect 541248 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 541568 136102
rect 541248 135978 541568 136046
rect 541248 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 541568 135978
rect 541248 135888 541568 135922
rect 571968 136350 572288 136384
rect 571968 136294 572038 136350
rect 572094 136294 572162 136350
rect 572218 136294 572288 136350
rect 571968 136226 572288 136294
rect 571968 136170 572038 136226
rect 572094 136170 572162 136226
rect 572218 136170 572288 136226
rect 571968 136102 572288 136170
rect 571968 136046 572038 136102
rect 572094 136046 572162 136102
rect 572218 136046 572288 136102
rect 571968 135978 572288 136046
rect 571968 135922 572038 135978
rect 572094 135922 572162 135978
rect 572218 135922 572288 135978
rect 571968 135888 572288 135922
rect 467068 134152 467124 134162
rect 466620 133972 466676 133982
rect 495168 130350 495488 130384
rect 495168 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 495488 130350
rect 495168 130226 495488 130294
rect 495168 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 495488 130226
rect 495168 130102 495488 130170
rect 495168 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 495488 130102
rect 495168 129978 495488 130046
rect 495168 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 495488 129978
rect 495168 129888 495488 129922
rect 525888 130350 526208 130384
rect 525888 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 526208 130350
rect 525888 130226 526208 130294
rect 525888 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 526208 130226
rect 525888 130102 526208 130170
rect 525888 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 526208 130102
rect 525888 129978 526208 130046
rect 525888 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 526208 129978
rect 525888 129888 526208 129922
rect 556608 130350 556928 130384
rect 556608 130294 556678 130350
rect 556734 130294 556802 130350
rect 556858 130294 556928 130350
rect 556608 130226 556928 130294
rect 556608 130170 556678 130226
rect 556734 130170 556802 130226
rect 556858 130170 556928 130226
rect 556608 130102 556928 130170
rect 556608 130046 556678 130102
rect 556734 130046 556802 130102
rect 556858 130046 556928 130102
rect 556608 129978 556928 130046
rect 556608 129922 556678 129978
rect 556734 129922 556802 129978
rect 556858 129922 556928 129978
rect 556608 129888 556928 129922
rect 466284 127492 466340 127502
rect 466172 122452 466228 122462
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 479808 118350 480128 118384
rect 479808 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 480128 118350
rect 479808 118226 480128 118294
rect 479808 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 480128 118226
rect 479808 118102 480128 118170
rect 479808 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 480128 118102
rect 479808 117978 480128 118046
rect 479808 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 480128 117978
rect 479808 117888 480128 117922
rect 510528 118350 510848 118384
rect 510528 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 510848 118350
rect 510528 118226 510848 118294
rect 510528 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 510848 118226
rect 510528 118102 510848 118170
rect 510528 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 510848 118102
rect 510528 117978 510848 118046
rect 510528 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 510848 117978
rect 510528 117888 510848 117922
rect 541248 118350 541568 118384
rect 541248 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 541568 118350
rect 541248 118226 541568 118294
rect 541248 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 541568 118226
rect 541248 118102 541568 118170
rect 541248 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 541568 118102
rect 541248 117978 541568 118046
rect 541248 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 541568 117978
rect 541248 117888 541568 117922
rect 571968 118350 572288 118384
rect 571968 118294 572038 118350
rect 572094 118294 572162 118350
rect 572218 118294 572288 118350
rect 571968 118226 572288 118294
rect 571968 118170 572038 118226
rect 572094 118170 572162 118226
rect 572218 118170 572288 118226
rect 571968 118102 572288 118170
rect 571968 118046 572038 118102
rect 572094 118046 572162 118102
rect 572218 118046 572288 118102
rect 571968 117978 572288 118046
rect 571968 117922 572038 117978
rect 572094 117922 572162 117978
rect 572218 117922 572288 117978
rect 571968 117888 572288 117922
rect 574140 113878 574196 137732
rect 574140 113812 574196 113822
rect 464448 112350 464768 112384
rect 464448 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 464768 112350
rect 464448 112226 464768 112294
rect 464448 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 464768 112226
rect 464448 112102 464768 112170
rect 464448 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 464768 112102
rect 464448 111978 464768 112046
rect 464448 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 464768 111978
rect 464448 111888 464768 111922
rect 495168 112350 495488 112384
rect 495168 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 495488 112350
rect 495168 112226 495488 112294
rect 495168 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 495488 112226
rect 495168 112102 495488 112170
rect 495168 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 495488 112102
rect 495168 111978 495488 112046
rect 495168 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 495488 111978
rect 495168 111888 495488 111922
rect 525888 112350 526208 112384
rect 525888 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 526208 112350
rect 525888 112226 526208 112294
rect 525888 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 526208 112226
rect 525888 112102 526208 112170
rect 525888 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 526208 112102
rect 525888 111978 526208 112046
rect 525888 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 526208 111978
rect 525888 111888 526208 111922
rect 556608 112350 556928 112384
rect 556608 112294 556678 112350
rect 556734 112294 556802 112350
rect 556858 112294 556928 112350
rect 556608 112226 556928 112294
rect 556608 112170 556678 112226
rect 556734 112170 556802 112226
rect 556858 112170 556928 112226
rect 556608 112102 556928 112170
rect 556608 112046 556678 112102
rect 556734 112046 556802 112102
rect 556858 112046 556928 112102
rect 556608 111978 556928 112046
rect 556608 111922 556678 111978
rect 556734 111922 556802 111978
rect 556858 111922 556928 111978
rect 556608 111888 556928 111922
rect 458108 110404 458164 110414
rect 457884 110180 457940 110190
rect 457772 106708 457828 106718
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 456988 101668 457044 101678
rect 456988 97636 457044 101612
rect 456988 97570 457044 97580
rect 457548 98644 457604 98654
rect 457548 85092 457604 98588
rect 457548 85026 457604 85036
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 457772 54852 457828 106652
rect 457884 58212 457940 110124
rect 457884 58146 457940 58156
rect 457996 98308 458052 98318
rect 457772 54786 457828 54796
rect 457996 48132 458052 98252
rect 458108 61572 458164 110348
rect 458556 101780 458612 101790
rect 458220 100100 458276 100110
rect 458220 64932 458276 100044
rect 458444 99988 458500 99998
rect 458332 98980 458388 98990
rect 458332 75012 458388 98924
rect 458332 74946 458388 74956
rect 458444 68292 458500 99932
rect 458556 88452 458612 101724
rect 479808 100350 480128 100384
rect 479808 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 480128 100350
rect 479808 100226 480128 100294
rect 479808 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 480128 100226
rect 479808 100102 480128 100170
rect 479808 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 480128 100102
rect 479808 99978 480128 100046
rect 479808 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 480128 99978
rect 479808 99888 480128 99922
rect 510528 100350 510848 100384
rect 510528 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 510848 100350
rect 510528 100226 510848 100294
rect 510528 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 510848 100226
rect 510528 100102 510848 100170
rect 510528 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 510848 100102
rect 510528 99978 510848 100046
rect 510528 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 510848 99978
rect 510528 99888 510848 99922
rect 541248 100350 541568 100384
rect 541248 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 541568 100350
rect 541248 100226 541568 100294
rect 541248 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 541568 100226
rect 541248 100102 541568 100170
rect 541248 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 541568 100102
rect 541248 99978 541568 100046
rect 541248 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 541568 99978
rect 541248 99888 541568 99922
rect 571968 100350 572288 100384
rect 571968 100294 572038 100350
rect 572094 100294 572162 100350
rect 572218 100294 572288 100350
rect 571968 100226 572288 100294
rect 571968 100170 572038 100226
rect 572094 100170 572162 100226
rect 572218 100170 572288 100226
rect 571968 100102 572288 100170
rect 571968 100046 572038 100102
rect 572094 100046 572162 100102
rect 572218 100046 572288 100102
rect 571968 99978 572288 100046
rect 571968 99922 572038 99978
rect 572094 99922 572162 99978
rect 572218 99922 572288 99978
rect 571968 99888 572288 99922
rect 464448 94350 464768 94384
rect 464448 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 464768 94350
rect 464448 94226 464768 94294
rect 464448 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 464768 94226
rect 464448 94102 464768 94170
rect 464448 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 464768 94102
rect 464448 93978 464768 94046
rect 464448 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 464768 93978
rect 464448 93888 464768 93922
rect 495168 94350 495488 94384
rect 495168 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 495488 94350
rect 495168 94226 495488 94294
rect 495168 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 495488 94226
rect 495168 94102 495488 94170
rect 495168 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 495488 94102
rect 495168 93978 495488 94046
rect 495168 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 495488 93978
rect 495168 93888 495488 93922
rect 525888 94350 526208 94384
rect 525888 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 526208 94350
rect 525888 94226 526208 94294
rect 525888 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 526208 94226
rect 525888 94102 526208 94170
rect 525888 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 526208 94102
rect 525888 93978 526208 94046
rect 525888 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 526208 93978
rect 525888 93888 526208 93922
rect 556608 94350 556928 94384
rect 556608 94294 556678 94350
rect 556734 94294 556802 94350
rect 556858 94294 556928 94350
rect 556608 94226 556928 94294
rect 556608 94170 556678 94226
rect 556734 94170 556802 94226
rect 556858 94170 556928 94226
rect 556608 94102 556928 94170
rect 556608 94046 556678 94102
rect 556734 94046 556802 94102
rect 556858 94046 556928 94102
rect 556608 93978 556928 94046
rect 556608 93922 556678 93978
rect 556734 93922 556802 93978
rect 556858 93922 556928 93978
rect 556608 93888 556928 93922
rect 458556 88386 458612 88396
rect 479808 82350 480128 82384
rect 479808 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 480128 82350
rect 479808 82226 480128 82294
rect 479808 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 480128 82226
rect 479808 82102 480128 82170
rect 479808 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 480128 82102
rect 479808 81978 480128 82046
rect 479808 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 480128 81978
rect 479808 81888 480128 81922
rect 510528 82350 510848 82384
rect 510528 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 510848 82350
rect 510528 82226 510848 82294
rect 510528 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 510848 82226
rect 510528 82102 510848 82170
rect 510528 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 510848 82102
rect 510528 81978 510848 82046
rect 510528 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 510848 81978
rect 510528 81888 510848 81922
rect 541248 82350 541568 82384
rect 541248 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 541568 82350
rect 541248 82226 541568 82294
rect 541248 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 541568 82226
rect 541248 82102 541568 82170
rect 541248 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 541568 82102
rect 541248 81978 541568 82046
rect 541248 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 541568 81978
rect 541248 81888 541568 81922
rect 571968 82350 572288 82384
rect 571968 82294 572038 82350
rect 572094 82294 572162 82350
rect 572218 82294 572288 82350
rect 571968 82226 572288 82294
rect 571968 82170 572038 82226
rect 572094 82170 572162 82226
rect 572218 82170 572288 82226
rect 571968 82102 572288 82170
rect 571968 82046 572038 82102
rect 572094 82046 572162 82102
rect 572218 82046 572288 82102
rect 571968 81978 572288 82046
rect 571968 81922 572038 81978
rect 572094 81922 572162 81978
rect 572218 81922 572288 81978
rect 571968 81888 572288 81922
rect 464448 76350 464768 76384
rect 464448 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 464768 76350
rect 464448 76226 464768 76294
rect 464448 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 464768 76226
rect 464448 76102 464768 76170
rect 464448 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 464768 76102
rect 464448 75978 464768 76046
rect 464448 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 464768 75978
rect 464448 75888 464768 75922
rect 495168 76350 495488 76384
rect 495168 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 495488 76350
rect 495168 76226 495488 76294
rect 495168 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 495488 76226
rect 495168 76102 495488 76170
rect 495168 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 495488 76102
rect 495168 75978 495488 76046
rect 495168 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 495488 75978
rect 495168 75888 495488 75922
rect 525888 76350 526208 76384
rect 525888 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 526208 76350
rect 525888 76226 526208 76294
rect 525888 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 526208 76226
rect 525888 76102 526208 76170
rect 525888 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 526208 76102
rect 525888 75978 526208 76046
rect 525888 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 526208 75978
rect 525888 75888 526208 75922
rect 556608 76350 556928 76384
rect 556608 76294 556678 76350
rect 556734 76294 556802 76350
rect 556858 76294 556928 76350
rect 556608 76226 556928 76294
rect 556608 76170 556678 76226
rect 556734 76170 556802 76226
rect 556858 76170 556928 76226
rect 556608 76102 556928 76170
rect 556608 76046 556678 76102
rect 556734 76046 556802 76102
rect 556858 76046 556928 76102
rect 556608 75978 556928 76046
rect 556608 75922 556678 75978
rect 556734 75922 556802 75978
rect 556858 75922 556928 75978
rect 556608 75888 556928 75922
rect 458444 68226 458500 68236
rect 458220 64866 458276 64876
rect 479808 64350 480128 64384
rect 479808 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 480128 64350
rect 479808 64226 480128 64294
rect 479808 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 480128 64226
rect 479808 64102 480128 64170
rect 479808 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 480128 64102
rect 479808 63978 480128 64046
rect 479808 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 480128 63978
rect 479808 63888 480128 63922
rect 510528 64350 510848 64384
rect 510528 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 510848 64350
rect 510528 64226 510848 64294
rect 510528 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 510848 64226
rect 510528 64102 510848 64170
rect 510528 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 510848 64102
rect 510528 63978 510848 64046
rect 510528 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 510848 63978
rect 510528 63888 510848 63922
rect 541248 64350 541568 64384
rect 541248 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 541568 64350
rect 541248 64226 541568 64294
rect 541248 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 541568 64226
rect 541248 64102 541568 64170
rect 541248 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 541568 64102
rect 541248 63978 541568 64046
rect 541248 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 541568 63978
rect 541248 63888 541568 63922
rect 571968 64350 572288 64384
rect 571968 64294 572038 64350
rect 572094 64294 572162 64350
rect 572218 64294 572288 64350
rect 571968 64226 572288 64294
rect 571968 64170 572038 64226
rect 572094 64170 572162 64226
rect 572218 64170 572288 64226
rect 571968 64102 572288 64170
rect 571968 64046 572038 64102
rect 572094 64046 572162 64102
rect 572218 64046 572288 64102
rect 571968 63978 572288 64046
rect 571968 63922 572038 63978
rect 572094 63922 572162 63978
rect 572218 63922 572288 63978
rect 571968 63888 572288 63922
rect 458108 61506 458164 61516
rect 574252 61138 574308 138482
rect 574476 61318 574532 153020
rect 574700 152180 574756 152190
rect 574588 145378 574644 145388
rect 574588 64932 574644 145322
rect 574700 75012 574756 152124
rect 574812 81060 574868 155582
rect 575036 148148 575092 148158
rect 574924 146998 574980 147008
rect 574924 83076 574980 146942
rect 575036 89684 575092 148092
rect 575148 113878 575204 113914
rect 575148 113810 575204 113820
rect 575036 89618 575092 89628
rect 574924 83010 574980 83020
rect 574812 80994 574868 81004
rect 574700 74946 574756 74956
rect 574588 64866 574644 64876
rect 574476 61262 574756 61318
rect 574252 61124 574644 61138
rect 574252 61082 574588 61124
rect 574588 61058 574644 61068
rect 574700 60958 574756 61262
rect 574476 60902 574756 60958
rect 464448 58350 464768 58384
rect 464448 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 464768 58350
rect 464448 58226 464768 58294
rect 464448 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 464768 58226
rect 464448 58102 464768 58170
rect 464448 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 464768 58102
rect 464448 57978 464768 58046
rect 464448 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 464768 57978
rect 464448 57888 464768 57922
rect 495168 58350 495488 58384
rect 495168 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 495488 58350
rect 495168 58226 495488 58294
rect 495168 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 495488 58226
rect 495168 58102 495488 58170
rect 495168 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 495488 58102
rect 495168 57978 495488 58046
rect 495168 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 495488 57978
rect 495168 57888 495488 57922
rect 525888 58350 526208 58384
rect 525888 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 526208 58350
rect 525888 58226 526208 58294
rect 525888 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 526208 58226
rect 525888 58102 526208 58170
rect 525888 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 526208 58102
rect 525888 57978 526208 58046
rect 525888 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 526208 57978
rect 525888 57888 526208 57922
rect 556608 58350 556928 58384
rect 556608 58294 556678 58350
rect 556734 58294 556802 58350
rect 556858 58294 556928 58350
rect 556608 58226 556928 58294
rect 556608 58170 556678 58226
rect 556734 58170 556802 58226
rect 556858 58170 556928 58226
rect 556608 58102 556928 58170
rect 556608 58046 556678 58102
rect 556734 58046 556802 58102
rect 556858 58046 556928 58102
rect 556608 57978 556928 58046
rect 556608 57922 556678 57978
rect 556734 57922 556802 57978
rect 556858 57922 556928 57978
rect 556608 57888 556928 57922
rect 574476 52836 574532 60902
rect 574476 52770 574532 52780
rect 457996 48066 458052 48076
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 457660 47908 457716 47918
rect 457660 44772 457716 47852
rect 479808 46350 480128 46384
rect 479808 46294 479878 46350
rect 479934 46294 480002 46350
rect 480058 46294 480128 46350
rect 479808 46226 480128 46294
rect 479808 46170 479878 46226
rect 479934 46170 480002 46226
rect 480058 46170 480128 46226
rect 479808 46102 480128 46170
rect 479808 46046 479878 46102
rect 479934 46046 480002 46102
rect 480058 46046 480128 46102
rect 479808 45978 480128 46046
rect 479808 45922 479878 45978
rect 479934 45922 480002 45978
rect 480058 45922 480128 45978
rect 479808 45888 480128 45922
rect 510528 46350 510848 46384
rect 510528 46294 510598 46350
rect 510654 46294 510722 46350
rect 510778 46294 510848 46350
rect 510528 46226 510848 46294
rect 510528 46170 510598 46226
rect 510654 46170 510722 46226
rect 510778 46170 510848 46226
rect 510528 46102 510848 46170
rect 510528 46046 510598 46102
rect 510654 46046 510722 46102
rect 510778 46046 510848 46102
rect 510528 45978 510848 46046
rect 510528 45922 510598 45978
rect 510654 45922 510722 45978
rect 510778 45922 510848 45978
rect 510528 45888 510848 45922
rect 541248 46350 541568 46384
rect 541248 46294 541318 46350
rect 541374 46294 541442 46350
rect 541498 46294 541568 46350
rect 541248 46226 541568 46294
rect 541248 46170 541318 46226
rect 541374 46170 541442 46226
rect 541498 46170 541568 46226
rect 541248 46102 541568 46170
rect 541248 46046 541318 46102
rect 541374 46046 541442 46102
rect 541498 46046 541568 46102
rect 541248 45978 541568 46046
rect 541248 45922 541318 45978
rect 541374 45922 541442 45978
rect 541498 45922 541568 45978
rect 541248 45888 541568 45922
rect 571968 46350 572288 46384
rect 571968 46294 572038 46350
rect 572094 46294 572162 46350
rect 572218 46294 572288 46350
rect 571968 46226 572288 46294
rect 571968 46170 572038 46226
rect 572094 46170 572162 46226
rect 572218 46170 572288 46226
rect 571968 46102 572288 46170
rect 571968 46046 572038 46102
rect 572094 46046 572162 46102
rect 572218 46046 572288 46102
rect 571968 45978 572288 46046
rect 571968 45922 572038 45978
rect 572094 45922 572162 45978
rect 572218 45922 572288 45978
rect 571968 45888 572288 45922
rect 457660 44706 457716 44716
rect 456988 44548 457044 44558
rect 456988 41412 457044 44492
rect 456988 41346 457044 41356
rect 457100 42868 457156 42878
rect 457100 38052 457156 42812
rect 576268 40740 576324 158642
rect 578508 155652 578564 155662
rect 578060 155458 578116 155468
rect 576380 149698 576436 149708
rect 576380 56868 576436 149642
rect 576380 56802 576436 56812
rect 576492 143220 576548 143230
rect 576492 54852 576548 143164
rect 577948 141958 578004 141968
rect 577948 58884 578004 141902
rect 578060 77028 578116 155402
rect 578396 150836 578452 150846
rect 578284 143108 578340 143118
rect 578060 76962 578116 76972
rect 578172 139076 578228 139086
rect 578172 66948 578228 139020
rect 578284 70980 578340 143052
rect 578396 79044 578452 150780
rect 578508 87108 578564 155596
rect 589098 148350 589718 165922
rect 590380 192164 590436 192174
rect 590380 160692 590436 192108
rect 590492 161038 590548 390348
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 590492 160972 590548 160982
rect 590604 350756 590660 350766
rect 590380 160626 590436 160636
rect 590604 158676 590660 350700
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 590716 311108 590772 311118
rect 590716 160580 590772 311052
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 590828 297892 590884 297902
rect 590828 160858 590884 297836
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 590828 160792 590884 160802
rect 590940 271460 590996 271470
rect 590716 160514 590772 160524
rect 590940 159348 590996 271404
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 590940 159282 590996 159292
rect 591052 258244 591108 258254
rect 590604 158610 590660 158620
rect 591052 157798 591108 258188
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 591164 231924 591220 231934
rect 591164 159460 591220 231868
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 591276 218596 591332 218606
rect 591276 161218 591332 218540
rect 591276 161152 591332 161162
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 591164 159394 591220 159404
rect 591276 159684 591332 159694
rect 591052 157732 591108 157742
rect 591276 154532 591332 159628
rect 591276 154466 591332 154476
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 590828 153748 590884 153758
rect 590044 152758 590100 152778
rect 590044 152674 590100 152684
rect 590604 152038 590660 152048
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 578732 142324 578788 142334
rect 578508 87042 578564 87052
rect 578620 138628 578676 138638
rect 578396 78978 578452 78988
rect 578620 72996 578676 138572
rect 578732 85092 578788 142268
rect 578844 140338 578900 140348
rect 578844 91140 578900 140282
rect 578844 91074 578900 91084
rect 589098 130350 589718 147922
rect 590492 150418 590548 150428
rect 590156 139438 590212 139450
rect 590156 139346 590212 139356
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 578732 85026 578788 85036
rect 578620 72930 578676 72940
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 578284 70914 578340 70924
rect 578172 66882 578228 66892
rect 577948 58818 578004 58828
rect 576492 54786 576548 54796
rect 589098 58350 589718 75922
rect 590492 60228 590548 150362
rect 590604 73444 590660 151982
rect 590716 141238 590772 141248
rect 590716 99876 590772 141182
rect 590828 113092 590884 153692
rect 590828 113026 590884 113036
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 590716 99810 590772 99820
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 590604 73378 590660 73388
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 590492 60162 590548 60172
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 576268 40674 576324 40684
rect 577948 50820 578004 50830
rect 464448 40350 464768 40384
rect 464448 40294 464518 40350
rect 464574 40294 464642 40350
rect 464698 40294 464768 40350
rect 464448 40226 464768 40294
rect 464448 40170 464518 40226
rect 464574 40170 464642 40226
rect 464698 40170 464768 40226
rect 464448 40102 464768 40170
rect 464448 40046 464518 40102
rect 464574 40046 464642 40102
rect 464698 40046 464768 40102
rect 464448 39978 464768 40046
rect 464448 39922 464518 39978
rect 464574 39922 464642 39978
rect 464698 39922 464768 39978
rect 464448 39888 464768 39922
rect 495168 40350 495488 40384
rect 495168 40294 495238 40350
rect 495294 40294 495362 40350
rect 495418 40294 495488 40350
rect 495168 40226 495488 40294
rect 495168 40170 495238 40226
rect 495294 40170 495362 40226
rect 495418 40170 495488 40226
rect 495168 40102 495488 40170
rect 495168 40046 495238 40102
rect 495294 40046 495362 40102
rect 495418 40046 495488 40102
rect 495168 39978 495488 40046
rect 495168 39922 495238 39978
rect 495294 39922 495362 39978
rect 495418 39922 495488 39978
rect 495168 39888 495488 39922
rect 525888 40350 526208 40384
rect 525888 40294 525958 40350
rect 526014 40294 526082 40350
rect 526138 40294 526208 40350
rect 525888 40226 526208 40294
rect 525888 40170 525958 40226
rect 526014 40170 526082 40226
rect 526138 40170 526208 40226
rect 525888 40102 526208 40170
rect 525888 40046 525958 40102
rect 526014 40046 526082 40102
rect 526138 40046 526208 40102
rect 525888 39978 526208 40046
rect 525888 39922 525958 39978
rect 526014 39922 526082 39978
rect 526138 39922 526208 39978
rect 525888 39888 526208 39922
rect 556608 40350 556928 40384
rect 556608 40294 556678 40350
rect 556734 40294 556802 40350
rect 556858 40294 556928 40350
rect 556608 40226 556928 40294
rect 556608 40170 556678 40226
rect 556734 40170 556802 40226
rect 556858 40170 556928 40226
rect 556608 40102 556928 40170
rect 556608 40046 556678 40102
rect 556734 40046 556802 40102
rect 556858 40046 556928 40102
rect 556608 39978 556928 40046
rect 556608 39922 556678 39978
rect 556734 39922 556802 39978
rect 556858 39922 556928 39978
rect 556608 39888 556928 39922
rect 457100 37986 457156 37996
rect 457660 37828 457716 37838
rect 457660 34692 457716 37772
rect 457660 34626 457716 34636
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 439218 -1120 439838 9922
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 22350 466838 34090
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 466218 4350 466838 21922
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 28350 470558 34090
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 479808 28350 480128 28384
rect 479808 28294 479878 28350
rect 479934 28294 480002 28350
rect 480058 28294 480128 28350
rect 479808 28226 480128 28294
rect 479808 28170 479878 28226
rect 479934 28170 480002 28226
rect 480058 28170 480128 28226
rect 479808 28102 480128 28170
rect 479808 28046 479878 28102
rect 479934 28046 480002 28102
rect 480058 28046 480128 28102
rect 479808 27978 480128 28046
rect 479808 27922 479878 27978
rect 479934 27922 480002 27978
rect 480058 27922 480128 27978
rect 479808 27888 480128 27922
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 22350 497558 34090
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 496938 4350 497558 21922
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 28350 501278 34090
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 510528 28350 510848 28384
rect 510528 28294 510598 28350
rect 510654 28294 510722 28350
rect 510778 28294 510848 28350
rect 510528 28226 510848 28294
rect 510528 28170 510598 28226
rect 510654 28170 510722 28226
rect 510778 28170 510848 28226
rect 510528 28102 510848 28170
rect 510528 28046 510598 28102
rect 510654 28046 510722 28102
rect 510778 28046 510848 28102
rect 510528 27978 510848 28046
rect 510528 27922 510598 27978
rect 510654 27922 510722 27978
rect 510778 27922 510848 27978
rect 510528 27888 510848 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 500658 -1120 501278 9922
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 22350 528278 34090
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 28350 531998 34090
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 531378 10350 531998 27922
rect 541248 28350 541568 28384
rect 541248 28294 541318 28350
rect 541374 28294 541442 28350
rect 541498 28294 541568 28350
rect 541248 28226 541568 28294
rect 541248 28170 541318 28226
rect 541374 28170 541442 28226
rect 541498 28170 541568 28226
rect 541248 28102 541568 28170
rect 541248 28046 541318 28102
rect 541374 28046 541442 28102
rect 541498 28046 541568 28102
rect 541248 27978 541568 28046
rect 541248 27922 541318 27978
rect 541374 27922 541442 27978
rect 541498 27922 541568 27978
rect 541248 27888 541568 27922
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 531378 -1120 531998 9922
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 22350 558998 34090
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 28350 562718 34090
rect 577948 31798 578004 50764
rect 578172 44772 578228 44782
rect 577948 31732 578004 31742
rect 578060 36708 578116 36718
rect 574588 30178 574644 30188
rect 574588 29316 574644 30122
rect 574588 29250 574644 29260
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 562098 10350 562718 27922
rect 571968 28350 572288 28384
rect 571968 28294 572038 28350
rect 572094 28294 572162 28350
rect 572218 28294 572288 28350
rect 571968 28226 572288 28294
rect 571968 28170 572038 28226
rect 572094 28170 572162 28226
rect 572218 28170 572288 28226
rect 571968 28102 572288 28170
rect 571968 28046 572038 28102
rect 572094 28046 572162 28102
rect 572218 28046 572288 28102
rect 571968 27978 572288 28046
rect 571968 27922 572038 27978
rect 572094 27922 572162 27978
rect 572218 27922 572288 27978
rect 571968 27888 572288 27922
rect 574588 26068 574644 26078
rect 574588 22932 574644 26012
rect 574588 22866 574644 22876
rect 578060 21588 578116 36652
rect 578172 33598 578228 44716
rect 578172 33532 578228 33542
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 578172 32676 578228 32686
rect 578172 22820 578228 32620
rect 578172 22754 578228 22764
rect 578060 21522 578116 21532
rect 589098 22350 589718 39922
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 589932 35218 589988 35228
rect 589932 33796 589988 35162
rect 589932 33730 589988 33740
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 4350 589718 21922
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect 4172 416762 4228 416818
rect 4284 410642 4340 410698
rect 4396 409382 4452 409438
rect 4508 409202 4564 409258
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect 4060 380222 4116 380278
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 4172 376262 4228 376318
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect 4060 206522 4116 206578
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 12572 402362 12628 402418
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 4620 247022 4676 247078
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 7532 378782 7588 378838
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 20076 384722 20132 384778
rect 18396 383642 18452 383698
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 9234 316294 9290 316350
rect 9358 316294 9414 316350
rect 9482 316294 9538 316350
rect 9606 316294 9662 316350
rect 9234 316170 9290 316226
rect 9358 316170 9414 316226
rect 9482 316170 9538 316226
rect 9606 316170 9662 316226
rect 9234 316046 9290 316102
rect 9358 316046 9414 316102
rect 9482 316046 9538 316102
rect 9606 316046 9662 316102
rect 9234 315922 9290 315978
rect 9358 315922 9414 315978
rect 9482 315922 9538 315978
rect 9606 315922 9662 315978
rect 9234 298294 9290 298350
rect 9358 298294 9414 298350
rect 9482 298294 9538 298350
rect 9606 298294 9662 298350
rect 9234 298170 9290 298226
rect 9358 298170 9414 298226
rect 9482 298170 9538 298226
rect 9606 298170 9662 298226
rect 9234 298046 9290 298102
rect 9358 298046 9414 298102
rect 9482 298046 9538 298102
rect 9606 298046 9662 298102
rect 9234 297922 9290 297978
rect 9358 297922 9414 297978
rect 9482 297922 9538 297978
rect 9606 297922 9662 297978
rect 14252 383282 14308 383338
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 4284 55322 4340 55378
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 16716 372122 16772 372178
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 31052 379142 31108 379198
rect 32732 378962 32788 379018
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 36234 310294 36290 310350
rect 36358 310294 36414 310350
rect 36482 310294 36538 310350
rect 36606 310294 36662 310350
rect 36234 310170 36290 310226
rect 36358 310170 36414 310226
rect 36482 310170 36538 310226
rect 36606 310170 36662 310226
rect 36234 310046 36290 310102
rect 36358 310046 36414 310102
rect 36482 310046 36538 310102
rect 36606 310046 36662 310102
rect 36234 309922 36290 309978
rect 36358 309922 36414 309978
rect 36482 309922 36538 309978
rect 36606 309922 36662 309978
rect 36234 292294 36290 292350
rect 36358 292294 36414 292350
rect 36482 292294 36538 292350
rect 36606 292294 36662 292350
rect 36234 292170 36290 292226
rect 36358 292170 36414 292226
rect 36482 292170 36538 292226
rect 36606 292170 36662 292226
rect 36234 292046 36290 292102
rect 36358 292046 36414 292102
rect 36482 292046 36538 292102
rect 36606 292046 36662 292102
rect 36234 291922 36290 291978
rect 36358 291922 36414 291978
rect 36482 291922 36538 291978
rect 36606 291922 36662 291978
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 35196 229202 35252 229258
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568294 40010 568350
rect 40078 568294 40134 568350
rect 40202 568294 40258 568350
rect 40326 568294 40382 568350
rect 39954 568170 40010 568226
rect 40078 568170 40134 568226
rect 40202 568170 40258 568226
rect 40326 568170 40382 568226
rect 39954 568046 40010 568102
rect 40078 568046 40134 568102
rect 40202 568046 40258 568102
rect 40326 568046 40382 568102
rect 39954 567922 40010 567978
rect 40078 567922 40134 567978
rect 40202 567922 40258 567978
rect 40326 567922 40382 567978
rect 39954 550294 40010 550350
rect 40078 550294 40134 550350
rect 40202 550294 40258 550350
rect 40326 550294 40382 550350
rect 39954 550170 40010 550226
rect 40078 550170 40134 550226
rect 40202 550170 40258 550226
rect 40326 550170 40382 550226
rect 39954 550046 40010 550102
rect 40078 550046 40134 550102
rect 40202 550046 40258 550102
rect 40326 550046 40382 550102
rect 39954 549922 40010 549978
rect 40078 549922 40134 549978
rect 40202 549922 40258 549978
rect 40326 549922 40382 549978
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 130346 580007 130402 580063
rect 130470 580007 130526 580063
rect 130594 580007 130650 580063
rect 130718 580007 130774 580063
rect 130346 579883 130402 579939
rect 130470 579883 130526 579939
rect 130594 579883 130650 579939
rect 130718 579883 130774 579939
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 101394 568294 101450 568350
rect 101518 568294 101574 568350
rect 101642 568294 101698 568350
rect 101766 568294 101822 568350
rect 101394 568170 101450 568226
rect 101518 568170 101574 568226
rect 101642 568170 101698 568226
rect 101766 568170 101822 568226
rect 101394 568046 101450 568102
rect 101518 568046 101574 568102
rect 101642 568046 101698 568102
rect 101766 568046 101822 568102
rect 101394 567922 101450 567978
rect 101518 567922 101574 567978
rect 101642 567922 101698 567978
rect 101766 567922 101822 567978
rect 116228 562216 116284 562272
rect 116352 562216 116408 562272
rect 116476 562216 116532 562272
rect 116600 562216 116656 562272
rect 116724 562216 116780 562272
rect 116848 562216 116904 562272
rect 116972 562216 117028 562272
rect 117096 562216 117152 562272
rect 117220 562216 117276 562272
rect 117344 562216 117400 562272
rect 117468 562216 117524 562272
rect 117592 562216 117648 562272
rect 117716 562216 117772 562272
rect 117840 562216 117896 562272
rect 117964 562216 118020 562272
rect 118088 562216 118144 562272
rect 118212 562216 118268 562272
rect 118336 562216 118392 562272
rect 118460 562216 118516 562272
rect 118584 562216 118640 562272
rect 118708 562216 118764 562272
rect 118832 562216 118888 562272
rect 118956 562216 119012 562272
rect 119080 562216 119136 562272
rect 119204 562216 119260 562272
rect 119328 562216 119384 562272
rect 119452 562216 119508 562272
rect 119576 562216 119632 562272
rect 119700 562216 119756 562272
rect 119824 562216 119880 562272
rect 119948 562216 120004 562272
rect 120072 562216 120128 562272
rect 120196 562216 120252 562272
rect 120320 562216 120376 562272
rect 120444 562216 120500 562272
rect 120568 562216 120624 562272
rect 120692 562216 120748 562272
rect 120816 562216 120872 562272
rect 120940 562216 120996 562272
rect 121064 562216 121120 562272
rect 121188 562216 121244 562272
rect 121312 562216 121368 562272
rect 121436 562216 121492 562272
rect 121560 562216 121616 562272
rect 121684 562216 121740 562272
rect 121808 562216 121864 562272
rect 121932 562216 121988 562272
rect 122056 562216 122112 562272
rect 122180 562216 122236 562272
rect 122304 562216 122360 562272
rect 122428 562216 122484 562272
rect 122552 562216 122608 562272
rect 122676 562216 122732 562272
rect 122800 562216 122856 562272
rect 122924 562216 122980 562272
rect 123048 562216 123104 562272
rect 123172 562216 123228 562272
rect 123296 562216 123352 562272
rect 123420 562216 123476 562272
rect 123544 562216 123600 562272
rect 123668 562216 123724 562272
rect 123792 562216 123848 562272
rect 123916 562216 123972 562272
rect 124040 562216 124096 562272
rect 124164 562216 124220 562272
rect 124288 562216 124344 562272
rect 124412 562216 124468 562272
rect 124536 562216 124592 562272
rect 124660 562216 124716 562272
rect 124784 562216 124840 562272
rect 124908 562216 124964 562272
rect 125032 562216 125088 562272
rect 125156 562216 125212 562272
rect 125280 562216 125336 562272
rect 125404 562216 125460 562272
rect 125528 562216 125584 562272
rect 125652 562216 125708 562272
rect 125776 562216 125832 562272
rect 125900 562216 125956 562272
rect 126024 562216 126080 562272
rect 126148 562216 126204 562272
rect 126272 562216 126328 562272
rect 126396 562216 126452 562272
rect 126520 562216 126576 562272
rect 126644 562216 126700 562272
rect 126768 562216 126824 562272
rect 126892 562216 126948 562272
rect 127016 562216 127072 562272
rect 127140 562216 127196 562272
rect 127264 562216 127320 562272
rect 127388 562216 127444 562272
rect 127512 562216 127568 562272
rect 127636 562216 127692 562272
rect 127760 562216 127816 562272
rect 127884 562216 127940 562272
rect 128008 562216 128064 562272
rect 128132 562216 128188 562272
rect 128256 562216 128312 562272
rect 128380 562216 128436 562272
rect 128504 562216 128560 562272
rect 128628 562216 128684 562272
rect 128752 562216 128808 562272
rect 128876 562216 128932 562272
rect 129000 562216 129056 562272
rect 129124 562216 129180 562272
rect 129248 562216 129304 562272
rect 129372 562216 129428 562272
rect 129496 562216 129552 562272
rect 129620 562216 129676 562272
rect 129744 562216 129800 562272
rect 129868 562216 129924 562272
rect 129992 562216 130048 562272
rect 130116 562216 130172 562272
rect 130240 562216 130296 562272
rect 130364 562216 130420 562272
rect 130488 562216 130544 562272
rect 130612 562216 130668 562272
rect 130736 562216 130792 562272
rect 130860 562216 130916 562272
rect 130984 562216 131040 562272
rect 131108 562216 131164 562272
rect 131232 562216 131288 562272
rect 131356 562216 131412 562272
rect 131480 562216 131536 562272
rect 131604 562216 131660 562272
rect 131728 562216 131784 562272
rect 131852 562216 131908 562272
rect 131976 562216 132032 562272
rect 132100 562216 132156 562272
rect 132224 562216 132280 562272
rect 132348 562216 132404 562272
rect 132472 562216 132528 562272
rect 132596 562216 132652 562272
rect 116228 562092 116284 562148
rect 116352 562092 116408 562148
rect 116476 562092 116532 562148
rect 116600 562092 116656 562148
rect 116724 562092 116780 562148
rect 116848 562092 116904 562148
rect 116972 562092 117028 562148
rect 117096 562092 117152 562148
rect 117220 562092 117276 562148
rect 117344 562092 117400 562148
rect 117468 562092 117524 562148
rect 117592 562092 117648 562148
rect 117716 562092 117772 562148
rect 117840 562092 117896 562148
rect 117964 562092 118020 562148
rect 118088 562092 118144 562148
rect 118212 562092 118268 562148
rect 118336 562092 118392 562148
rect 118460 562092 118516 562148
rect 118584 562092 118640 562148
rect 118708 562092 118764 562148
rect 118832 562092 118888 562148
rect 118956 562092 119012 562148
rect 119080 562092 119136 562148
rect 119204 562092 119260 562148
rect 119328 562092 119384 562148
rect 119452 562092 119508 562148
rect 119576 562092 119632 562148
rect 119700 562092 119756 562148
rect 119824 562092 119880 562148
rect 119948 562092 120004 562148
rect 120072 562092 120128 562148
rect 120196 562092 120252 562148
rect 120320 562092 120376 562148
rect 120444 562092 120500 562148
rect 120568 562092 120624 562148
rect 120692 562092 120748 562148
rect 120816 562092 120872 562148
rect 120940 562092 120996 562148
rect 121064 562092 121120 562148
rect 121188 562092 121244 562148
rect 121312 562092 121368 562148
rect 121436 562092 121492 562148
rect 121560 562092 121616 562148
rect 121684 562092 121740 562148
rect 121808 562092 121864 562148
rect 121932 562092 121988 562148
rect 122056 562092 122112 562148
rect 122180 562092 122236 562148
rect 122304 562092 122360 562148
rect 122428 562092 122484 562148
rect 122552 562092 122608 562148
rect 122676 562092 122732 562148
rect 122800 562092 122856 562148
rect 122924 562092 122980 562148
rect 123048 562092 123104 562148
rect 123172 562092 123228 562148
rect 123296 562092 123352 562148
rect 123420 562092 123476 562148
rect 123544 562092 123600 562148
rect 123668 562092 123724 562148
rect 123792 562092 123848 562148
rect 123916 562092 123972 562148
rect 124040 562092 124096 562148
rect 124164 562092 124220 562148
rect 124288 562092 124344 562148
rect 124412 562092 124468 562148
rect 124536 562092 124592 562148
rect 124660 562092 124716 562148
rect 124784 562092 124840 562148
rect 124908 562092 124964 562148
rect 125032 562092 125088 562148
rect 125156 562092 125212 562148
rect 125280 562092 125336 562148
rect 125404 562092 125460 562148
rect 125528 562092 125584 562148
rect 125652 562092 125708 562148
rect 125776 562092 125832 562148
rect 125900 562092 125956 562148
rect 126024 562092 126080 562148
rect 126148 562092 126204 562148
rect 126272 562092 126328 562148
rect 126396 562092 126452 562148
rect 126520 562092 126576 562148
rect 126644 562092 126700 562148
rect 126768 562092 126824 562148
rect 126892 562092 126948 562148
rect 127016 562092 127072 562148
rect 127140 562092 127196 562148
rect 127264 562092 127320 562148
rect 127388 562092 127444 562148
rect 127512 562092 127568 562148
rect 127636 562092 127692 562148
rect 127760 562092 127816 562148
rect 127884 562092 127940 562148
rect 128008 562092 128064 562148
rect 128132 562092 128188 562148
rect 128256 562092 128312 562148
rect 128380 562092 128436 562148
rect 128504 562092 128560 562148
rect 128628 562092 128684 562148
rect 128752 562092 128808 562148
rect 128876 562092 128932 562148
rect 129000 562092 129056 562148
rect 129124 562092 129180 562148
rect 129248 562092 129304 562148
rect 129372 562092 129428 562148
rect 129496 562092 129552 562148
rect 129620 562092 129676 562148
rect 129744 562092 129800 562148
rect 129868 562092 129924 562148
rect 129992 562092 130048 562148
rect 130116 562092 130172 562148
rect 130240 562092 130296 562148
rect 130364 562092 130420 562148
rect 130488 562092 130544 562148
rect 130612 562092 130668 562148
rect 130736 562092 130792 562148
rect 130860 562092 130916 562148
rect 130984 562092 131040 562148
rect 131108 562092 131164 562148
rect 131232 562092 131288 562148
rect 131356 562092 131412 562148
rect 131480 562092 131536 562148
rect 131604 562092 131660 562148
rect 131728 562092 131784 562148
rect 131852 562092 131908 562148
rect 131976 562092 132032 562148
rect 132100 562092 132156 562148
rect 132224 562092 132280 562148
rect 132348 562092 132404 562148
rect 132472 562092 132528 562148
rect 132596 562092 132652 562148
rect 116228 561968 116284 562024
rect 116352 561968 116408 562024
rect 116476 561968 116532 562024
rect 116600 561968 116656 562024
rect 116724 561968 116780 562024
rect 116848 561968 116904 562024
rect 116972 561968 117028 562024
rect 117096 561968 117152 562024
rect 117220 561968 117276 562024
rect 117344 561968 117400 562024
rect 117468 561968 117524 562024
rect 117592 561968 117648 562024
rect 117716 561968 117772 562024
rect 117840 561968 117896 562024
rect 117964 561968 118020 562024
rect 118088 561968 118144 562024
rect 118212 561968 118268 562024
rect 118336 561968 118392 562024
rect 118460 561968 118516 562024
rect 118584 561968 118640 562024
rect 118708 561968 118764 562024
rect 118832 561968 118888 562024
rect 118956 561968 119012 562024
rect 119080 561968 119136 562024
rect 119204 561968 119260 562024
rect 119328 561968 119384 562024
rect 119452 561968 119508 562024
rect 119576 561968 119632 562024
rect 119700 561968 119756 562024
rect 119824 561968 119880 562024
rect 119948 561968 120004 562024
rect 120072 561968 120128 562024
rect 120196 561968 120252 562024
rect 120320 561968 120376 562024
rect 120444 561968 120500 562024
rect 120568 561968 120624 562024
rect 120692 561968 120748 562024
rect 120816 561968 120872 562024
rect 120940 561968 120996 562024
rect 121064 561968 121120 562024
rect 121188 561968 121244 562024
rect 121312 561968 121368 562024
rect 121436 561968 121492 562024
rect 121560 561968 121616 562024
rect 121684 561968 121740 562024
rect 121808 561968 121864 562024
rect 121932 561968 121988 562024
rect 122056 561968 122112 562024
rect 122180 561968 122236 562024
rect 122304 561968 122360 562024
rect 122428 561968 122484 562024
rect 122552 561968 122608 562024
rect 122676 561968 122732 562024
rect 122800 561968 122856 562024
rect 122924 561968 122980 562024
rect 123048 561968 123104 562024
rect 123172 561968 123228 562024
rect 123296 561968 123352 562024
rect 123420 561968 123476 562024
rect 123544 561968 123600 562024
rect 123668 561968 123724 562024
rect 123792 561968 123848 562024
rect 123916 561968 123972 562024
rect 124040 561968 124096 562024
rect 124164 561968 124220 562024
rect 124288 561968 124344 562024
rect 124412 561968 124468 562024
rect 124536 561968 124592 562024
rect 124660 561968 124716 562024
rect 124784 561968 124840 562024
rect 124908 561968 124964 562024
rect 125032 561968 125088 562024
rect 125156 561968 125212 562024
rect 125280 561968 125336 562024
rect 125404 561968 125460 562024
rect 125528 561968 125584 562024
rect 125652 561968 125708 562024
rect 125776 561968 125832 562024
rect 125900 561968 125956 562024
rect 126024 561968 126080 562024
rect 126148 561968 126204 562024
rect 126272 561968 126328 562024
rect 126396 561968 126452 562024
rect 126520 561968 126576 562024
rect 126644 561968 126700 562024
rect 126768 561968 126824 562024
rect 126892 561968 126948 562024
rect 127016 561968 127072 562024
rect 127140 561968 127196 562024
rect 127264 561968 127320 562024
rect 127388 561968 127444 562024
rect 127512 561968 127568 562024
rect 127636 561968 127692 562024
rect 127760 561968 127816 562024
rect 127884 561968 127940 562024
rect 128008 561968 128064 562024
rect 128132 561968 128188 562024
rect 128256 561968 128312 562024
rect 128380 561968 128436 562024
rect 128504 561968 128560 562024
rect 128628 561968 128684 562024
rect 128752 561968 128808 562024
rect 128876 561968 128932 562024
rect 129000 561968 129056 562024
rect 129124 561968 129180 562024
rect 129248 561968 129304 562024
rect 129372 561968 129428 562024
rect 129496 561968 129552 562024
rect 129620 561968 129676 562024
rect 129744 561968 129800 562024
rect 129868 561968 129924 562024
rect 129992 561968 130048 562024
rect 130116 561968 130172 562024
rect 130240 561968 130296 562024
rect 130364 561968 130420 562024
rect 130488 561968 130544 562024
rect 130612 561968 130668 562024
rect 130736 561968 130792 562024
rect 130860 561968 130916 562024
rect 130984 561968 131040 562024
rect 131108 561968 131164 562024
rect 131232 561968 131288 562024
rect 131356 561968 131412 562024
rect 131480 561968 131536 562024
rect 131604 561968 131660 562024
rect 131728 561968 131784 562024
rect 131852 561968 131908 562024
rect 131976 561968 132032 562024
rect 132100 561968 132156 562024
rect 132224 561968 132280 562024
rect 132348 561968 132404 562024
rect 132472 561968 132528 562024
rect 132596 561968 132652 562024
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 101394 550294 101450 550350
rect 101518 550294 101574 550350
rect 101642 550294 101698 550350
rect 101766 550294 101822 550350
rect 101394 550170 101450 550226
rect 101518 550170 101574 550226
rect 101642 550170 101698 550226
rect 101766 550170 101822 550226
rect 101394 550046 101450 550102
rect 101518 550046 101574 550102
rect 101642 550046 101698 550102
rect 101766 550046 101822 550102
rect 101394 549922 101450 549978
rect 101518 549922 101574 549978
rect 101642 549922 101698 549978
rect 101766 549922 101822 549978
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 104348 544002 104404 544058
rect 104472 544002 104528 544058
rect 104596 544002 104652 544058
rect 104720 544002 104776 544058
rect 104844 544002 104900 544058
rect 104968 544002 105024 544058
rect 105092 544002 105148 544058
rect 105216 544002 105272 544058
rect 105340 544002 105396 544058
rect 105464 544002 105520 544058
rect 105588 544002 105644 544058
rect 105712 544002 105768 544058
rect 105836 544002 105892 544058
rect 105960 544002 106016 544058
rect 106084 544002 106140 544058
rect 106208 544002 106264 544058
rect 106332 544002 106388 544058
rect 106456 544002 106512 544058
rect 106580 544002 106636 544058
rect 106704 544002 106760 544058
rect 106828 544002 106884 544058
rect 106952 544002 107008 544058
rect 107076 544002 107132 544058
rect 107200 544002 107256 544058
rect 107324 544002 107380 544058
rect 107448 544002 107504 544058
rect 107572 544002 107628 544058
rect 107696 544002 107752 544058
rect 107820 544002 107876 544058
rect 107944 544002 108000 544058
rect 108068 544002 108124 544058
rect 108192 544002 108248 544058
rect 108316 544002 108372 544058
rect 108440 544002 108496 544058
rect 108564 544002 108620 544058
rect 108688 544002 108744 544058
rect 108812 544002 108868 544058
rect 108936 544002 108992 544058
rect 109060 544002 109116 544058
rect 109184 544002 109240 544058
rect 109308 544002 109364 544058
rect 109432 544002 109488 544058
rect 109556 544002 109612 544058
rect 109680 544002 109736 544058
rect 109804 544002 109860 544058
rect 109928 544002 109984 544058
rect 110052 544002 110108 544058
rect 110176 544002 110232 544058
rect 110300 544002 110356 544058
rect 110424 544002 110480 544058
rect 110548 544002 110604 544058
rect 110672 544002 110728 544058
rect 110796 544002 110852 544058
rect 110920 544002 110976 544058
rect 111044 544002 111100 544058
rect 111168 544002 111224 544058
rect 111292 544002 111348 544058
rect 111416 544002 111472 544058
rect 111540 544002 111596 544058
rect 111664 544002 111720 544058
rect 111788 544002 111844 544058
rect 111912 544002 111968 544058
rect 112036 544002 112092 544058
rect 112160 544002 112216 544058
rect 112284 544002 112340 544058
rect 112408 544002 112464 544058
rect 112532 544002 112588 544058
rect 112656 544002 112712 544058
rect 112780 544002 112836 544058
rect 112904 544002 112960 544058
rect 113028 544002 113084 544058
rect 113152 544002 113208 544058
rect 113276 544002 113332 544058
rect 113400 544002 113456 544058
rect 113524 544002 113580 544058
rect 113648 544002 113704 544058
rect 113772 544002 113828 544058
rect 113896 544002 113952 544058
rect 114020 544002 114076 544058
rect 114144 544002 114200 544058
rect 114268 544002 114324 544058
rect 114392 544002 114448 544058
rect 114516 544002 114572 544058
rect 114640 544002 114696 544058
rect 114764 544002 114820 544058
rect 114888 544002 114944 544058
rect 115012 544002 115068 544058
rect 115136 544002 115192 544058
rect 115260 544002 115316 544058
rect 115384 544002 115440 544058
rect 115508 544002 115564 544058
rect 115632 544002 115688 544058
rect 115756 544002 115812 544058
rect 115880 544002 115936 544058
rect 116004 544002 116060 544058
rect 116128 544002 116184 544058
rect 116252 544002 116308 544058
rect 116376 544002 116432 544058
rect 116500 544002 116556 544058
rect 116624 544002 116680 544058
rect 116748 544002 116804 544058
rect 116872 544002 116928 544058
rect 116996 544002 117052 544058
rect 117120 544002 117176 544058
rect 117244 544002 117300 544058
rect 117368 544002 117424 544058
rect 117492 544002 117548 544058
rect 117616 544002 117672 544058
rect 117740 544002 117796 544058
rect 117864 544002 117920 544058
rect 117988 544002 118044 544058
rect 118112 544002 118168 544058
rect 118236 544002 118292 544058
rect 118360 544002 118416 544058
rect 118484 544002 118540 544058
rect 118608 544002 118664 544058
rect 118732 544002 118788 544058
rect 118856 544002 118912 544058
rect 118980 544002 119036 544058
rect 119104 544002 119160 544058
rect 119228 544002 119284 544058
rect 119352 544002 119408 544058
rect 119476 544002 119532 544058
rect 119600 544002 119656 544058
rect 119724 544002 119780 544058
rect 119848 544002 119904 544058
rect 119972 544002 120028 544058
rect 120096 544002 120152 544058
rect 120220 544002 120276 544058
rect 120344 544002 120400 544058
rect 120468 544002 120524 544058
rect 120592 544002 120648 544058
rect 120716 544002 120772 544058
rect 120840 544002 120896 544058
rect 120964 544002 121020 544058
rect 121088 544002 121144 544058
rect 121212 544002 121268 544058
rect 121336 544002 121392 544058
rect 121460 544002 121516 544058
rect 121584 544002 121640 544058
rect 121708 544002 121764 544058
rect 121832 544002 121888 544058
rect 121956 544002 122012 544058
rect 122080 544002 122136 544058
rect 122204 544002 122260 544058
rect 122328 544002 122384 544058
rect 122452 544002 122508 544058
rect 122576 544002 122632 544058
rect 122700 544002 122756 544058
rect 122824 544002 122880 544058
rect 122948 544002 123004 544058
rect 123072 544002 123128 544058
rect 123196 544002 123252 544058
rect 123320 544002 123376 544058
rect 123444 544002 123500 544058
rect 123568 544002 123624 544058
rect 123692 544002 123748 544058
rect 123816 544002 123872 544058
rect 123940 544002 123996 544058
rect 124064 544002 124120 544058
rect 124188 544002 124244 544058
rect 124312 544002 124368 544058
rect 124436 544002 124492 544058
rect 124560 544002 124616 544058
rect 124684 544002 124740 544058
rect 124808 544002 124864 544058
rect 124932 544002 124988 544058
rect 125056 544002 125112 544058
rect 125180 544002 125236 544058
rect 125304 544002 125360 544058
rect 125428 544002 125484 544058
rect 125552 544002 125608 544058
rect 125676 544002 125732 544058
rect 125800 544002 125856 544058
rect 125924 544002 125980 544058
rect 126048 544002 126104 544058
rect 126172 544002 126228 544058
rect 126296 544002 126352 544058
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 39954 532294 40010 532350
rect 40078 532294 40134 532350
rect 40202 532294 40258 532350
rect 40326 532294 40382 532350
rect 66714 532302 66770 532358
rect 66838 532302 66894 532358
rect 66962 532302 67018 532358
rect 67086 532302 67142 532358
rect 67210 532302 67266 532358
rect 67334 532302 67390 532358
rect 67458 532302 67514 532358
rect 67582 532302 67638 532358
rect 67706 532302 67762 532358
rect 67830 532302 67886 532358
rect 67954 532302 68010 532358
rect 68078 532302 68134 532358
rect 68202 532302 68258 532358
rect 68326 532302 68382 532358
rect 68450 532302 68506 532358
rect 68574 532302 68630 532358
rect 68698 532302 68754 532358
rect 68822 532302 68878 532358
rect 68946 532302 69002 532358
rect 69070 532302 69126 532358
rect 69194 532302 69250 532358
rect 69318 532302 69374 532358
rect 69442 532302 69498 532358
rect 69566 532302 69622 532358
rect 69690 532302 69746 532358
rect 69814 532302 69870 532358
rect 69938 532302 69994 532358
rect 70062 532302 70118 532358
rect 70186 532302 70242 532358
rect 70310 532302 70366 532358
rect 70434 532302 70490 532358
rect 70558 532302 70614 532358
rect 70682 532302 70738 532358
rect 70806 532302 70862 532358
rect 70930 532302 70986 532358
rect 71054 532302 71110 532358
rect 71178 532302 71234 532358
rect 71302 532302 71358 532358
rect 71426 532302 71482 532358
rect 71550 532302 71606 532358
rect 71674 532302 71730 532358
rect 71798 532302 71854 532358
rect 71922 532302 71978 532358
rect 72046 532302 72102 532358
rect 72170 532302 72226 532358
rect 72294 532302 72350 532358
rect 72418 532302 72474 532358
rect 72542 532302 72598 532358
rect 72666 532302 72722 532358
rect 72790 532302 72846 532358
rect 72914 532302 72970 532358
rect 73038 532302 73094 532358
rect 73162 532302 73218 532358
rect 73286 532302 73342 532358
rect 73410 532302 73466 532358
rect 73534 532302 73590 532358
rect 73658 532302 73714 532358
rect 73782 532302 73838 532358
rect 73906 532302 73962 532358
rect 74030 532302 74086 532358
rect 74154 532302 74210 532358
rect 74278 532302 74334 532358
rect 74402 532302 74458 532358
rect 74526 532302 74582 532358
rect 74650 532302 74706 532358
rect 39954 532170 40010 532226
rect 40078 532170 40134 532226
rect 40202 532170 40258 532226
rect 40326 532170 40382 532226
rect 39954 532046 40010 532102
rect 40078 532046 40134 532102
rect 40202 532046 40258 532102
rect 40326 532046 40382 532102
rect 39954 531922 40010 531978
rect 40078 531922 40134 531978
rect 40202 531922 40258 531978
rect 40326 531922 40382 531978
rect 66506 531942 66562 531998
rect 66630 531942 66686 531998
rect 66754 531942 66810 531998
rect 66878 531942 66934 531998
rect 67002 531942 67058 531998
rect 67126 531942 67182 531998
rect 67250 531942 67306 531998
rect 67374 531942 67430 531998
rect 67498 531942 67554 531998
rect 67622 531942 67678 531998
rect 67746 531942 67802 531998
rect 67870 531942 67926 531998
rect 67994 531942 68050 531998
rect 68118 531942 68174 531998
rect 68242 531942 68298 531998
rect 68366 531942 68422 531998
rect 68490 531942 68546 531998
rect 68614 531942 68670 531998
rect 68738 531942 68794 531998
rect 68862 531942 68918 531998
rect 68986 531942 69042 531998
rect 69110 531942 69166 531998
rect 69234 531942 69290 531998
rect 69358 531942 69414 531998
rect 69482 531942 69538 531998
rect 69606 531942 69662 531998
rect 69730 531942 69786 531998
rect 69854 531942 69910 531998
rect 69978 531942 70034 531998
rect 70102 531942 70158 531998
rect 70226 531942 70282 531998
rect 70350 531942 70406 531998
rect 70474 531942 70530 531998
rect 70598 531942 70654 531998
rect 70722 531942 70778 531998
rect 70846 531942 70902 531998
rect 70970 531942 71026 531998
rect 71094 531942 71150 531998
rect 71218 531942 71274 531998
rect 71342 531942 71398 531998
rect 71466 531942 71522 531998
rect 71590 531942 71646 531998
rect 71714 531942 71770 531998
rect 71838 531942 71894 531998
rect 71962 531942 72018 531998
rect 72086 531942 72142 531998
rect 72210 531942 72266 531998
rect 72334 531942 72390 531998
rect 72458 531942 72514 531998
rect 72582 531942 72638 531998
rect 72706 531942 72762 531998
rect 72830 531942 72886 531998
rect 72954 531942 73010 531998
rect 73078 531942 73134 531998
rect 73202 531942 73258 531998
rect 73326 531942 73382 531998
rect 73450 531942 73506 531998
rect 73574 531942 73630 531998
rect 73698 531942 73754 531998
rect 73822 531942 73878 531998
rect 73946 531942 74002 531998
rect 74070 531942 74126 531998
rect 74194 531942 74250 531998
rect 74318 531942 74374 531998
rect 39954 514294 40010 514350
rect 40078 514294 40134 514350
rect 40202 514294 40258 514350
rect 40326 514294 40382 514350
rect 39954 514170 40010 514226
rect 40078 514170 40134 514226
rect 40202 514170 40258 514226
rect 40326 514170 40382 514226
rect 39954 514046 40010 514102
rect 40078 514046 40134 514102
rect 40202 514046 40258 514102
rect 40326 514046 40382 514102
rect 39954 513922 40010 513978
rect 40078 513922 40134 513978
rect 40202 513922 40258 513978
rect 40326 513922 40382 513978
rect 39954 496294 40010 496350
rect 40078 496294 40134 496350
rect 40202 496294 40258 496350
rect 40326 496294 40382 496350
rect 39954 496170 40010 496226
rect 40078 496170 40134 496226
rect 40202 496170 40258 496226
rect 40326 496170 40382 496226
rect 39954 496046 40010 496102
rect 40078 496046 40134 496102
rect 40202 496046 40258 496102
rect 40326 496046 40382 496102
rect 39954 495922 40010 495978
rect 40078 495922 40134 495978
rect 40202 495922 40258 495978
rect 40326 495922 40382 495978
rect 39954 478294 40010 478350
rect 40078 478294 40134 478350
rect 40202 478294 40258 478350
rect 40326 478294 40382 478350
rect 39954 478170 40010 478226
rect 40078 478170 40134 478226
rect 40202 478170 40258 478226
rect 40326 478170 40382 478226
rect 39954 478046 40010 478102
rect 40078 478046 40134 478102
rect 40202 478046 40258 478102
rect 40326 478046 40382 478102
rect 39954 477922 40010 477978
rect 40078 477922 40134 477978
rect 40202 477922 40258 477978
rect 40326 477922 40382 477978
rect 39954 460294 40010 460350
rect 40078 460294 40134 460350
rect 40202 460294 40258 460350
rect 40326 460294 40382 460350
rect 39954 460170 40010 460226
rect 40078 460170 40134 460226
rect 40202 460170 40258 460226
rect 40326 460170 40382 460226
rect 39954 460046 40010 460102
rect 40078 460046 40134 460102
rect 40202 460046 40258 460102
rect 40326 460046 40382 460102
rect 39954 459922 40010 459978
rect 40078 459922 40134 459978
rect 40202 459922 40258 459978
rect 40326 459922 40382 459978
rect 39954 442294 40010 442350
rect 40078 442294 40134 442350
rect 40202 442294 40258 442350
rect 40326 442294 40382 442350
rect 39954 442170 40010 442226
rect 40078 442170 40134 442226
rect 40202 442170 40258 442226
rect 40326 442170 40382 442226
rect 39954 442046 40010 442102
rect 40078 442046 40134 442102
rect 40202 442046 40258 442102
rect 40326 442046 40382 442102
rect 39954 441922 40010 441978
rect 40078 441922 40134 441978
rect 40202 441922 40258 441978
rect 40326 441922 40382 441978
rect 39954 424294 40010 424350
rect 40078 424294 40134 424350
rect 40202 424294 40258 424350
rect 40326 424294 40382 424350
rect 39954 424170 40010 424226
rect 40078 424170 40134 424226
rect 40202 424170 40258 424226
rect 40326 424170 40382 424226
rect 39954 424046 40010 424102
rect 40078 424046 40134 424102
rect 40202 424046 40258 424102
rect 40326 424046 40382 424102
rect 39954 423922 40010 423978
rect 40078 423922 40134 423978
rect 40202 423922 40258 423978
rect 40326 423922 40382 423978
rect 39954 406294 40010 406350
rect 40078 406294 40134 406350
rect 40202 406294 40258 406350
rect 40326 406294 40382 406350
rect 39954 406170 40010 406226
rect 40078 406170 40134 406226
rect 40202 406170 40258 406226
rect 40326 406170 40382 406226
rect 39954 406046 40010 406102
rect 40078 406046 40134 406102
rect 40202 406046 40258 406102
rect 40326 406046 40382 406102
rect 39954 405922 40010 405978
rect 40078 405922 40134 405978
rect 40202 405922 40258 405978
rect 40326 405922 40382 405978
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 95846 526002 95902 526058
rect 95970 526002 96026 526058
rect 96094 526002 96150 526058
rect 96218 526002 96274 526058
rect 96342 526002 96398 526058
rect 96466 526002 96522 526058
rect 96590 526002 96646 526058
rect 96714 526002 96770 526058
rect 96838 526002 96894 526058
rect 96962 526002 97018 526058
rect 97086 526002 97142 526058
rect 97210 526002 97266 526058
rect 97334 526002 97390 526058
rect 97458 526002 97514 526058
rect 97582 526002 97638 526058
rect 97706 526002 97762 526058
rect 97830 526002 97886 526058
rect 97954 526002 98010 526058
rect 98078 526002 98134 526058
rect 98202 526002 98258 526058
rect 98326 526002 98382 526058
rect 98450 526002 98506 526058
rect 98574 526002 98630 526058
rect 98698 526002 98754 526058
rect 98822 526002 98878 526058
rect 98946 526002 99002 526058
rect 99070 526002 99126 526058
rect 99194 526002 99250 526058
rect 99318 526002 99374 526058
rect 99442 526002 99498 526058
rect 99566 526002 99622 526058
rect 99690 526002 99746 526058
rect 99814 526002 99870 526058
rect 99938 526002 99994 526058
rect 100062 526002 100118 526058
rect 100186 526002 100242 526058
rect 100310 526002 100366 526058
rect 100434 526002 100490 526058
rect 100558 526002 100614 526058
rect 100682 526002 100738 526058
rect 100806 526002 100862 526058
rect 100930 526002 100986 526058
rect 101054 526002 101110 526058
rect 101178 526002 101234 526058
rect 101302 526002 101358 526058
rect 101426 526002 101482 526058
rect 101550 526002 101606 526058
rect 101674 526002 101730 526058
rect 101798 526002 101854 526058
rect 101922 526002 101978 526058
rect 102046 526002 102102 526058
rect 102170 526002 102226 526058
rect 102294 526002 102350 526058
rect 102418 526002 102474 526058
rect 102542 526002 102598 526058
rect 102666 526002 102722 526058
rect 102790 526002 102846 526058
rect 102914 526002 102970 526058
rect 103038 526002 103094 526058
rect 103162 526002 103218 526058
rect 103286 526002 103342 526058
rect 103410 526002 103466 526058
rect 103534 526002 103590 526058
rect 103658 526002 103714 526058
rect 103782 526002 103838 526058
rect 103906 526002 103962 526058
rect 104030 526002 104086 526058
rect 104154 526002 104210 526058
rect 104278 526002 104334 526058
rect 104402 526002 104458 526058
rect 104526 526002 104582 526058
rect 104650 526002 104706 526058
rect 104774 526002 104830 526058
rect 104898 526002 104954 526058
rect 105022 526002 105078 526058
rect 105146 526002 105202 526058
rect 105270 526002 105326 526058
rect 105394 526002 105450 526058
rect 105518 526002 105574 526058
rect 105642 526002 105698 526058
rect 105766 526002 105822 526058
rect 105890 526002 105946 526058
rect 106014 526002 106070 526058
rect 106138 526002 106194 526058
rect 106262 526002 106318 526058
rect 106386 526002 106442 526058
rect 106510 526002 106566 526058
rect 106634 526002 106690 526058
rect 106758 526002 106814 526058
rect 106882 526002 106938 526058
rect 107006 526002 107062 526058
rect 107130 526002 107186 526058
rect 107254 526002 107310 526058
rect 107378 526002 107434 526058
rect 107502 526002 107558 526058
rect 107626 526002 107682 526058
rect 107750 526002 107806 526058
rect 107874 526002 107930 526058
rect 107998 526002 108054 526058
rect 108122 526002 108178 526058
rect 108246 526002 108302 526058
rect 108370 526002 108426 526058
rect 108494 526002 108550 526058
rect 108618 526002 108674 526058
rect 108742 526002 108798 526058
rect 108866 526002 108922 526058
rect 108990 526002 109046 526058
rect 109114 526002 109170 526058
rect 109238 526002 109294 526058
rect 109362 526002 109418 526058
rect 109486 526002 109542 526058
rect 109610 526002 109666 526058
rect 109734 526002 109790 526058
rect 109858 526002 109914 526058
rect 109982 526002 110038 526058
rect 110106 526002 110162 526058
rect 110230 526002 110286 526058
rect 110354 526002 110410 526058
rect 110478 526002 110534 526058
rect 110602 526002 110658 526058
rect 110726 526002 110782 526058
rect 110850 526002 110906 526058
rect 110974 526002 111030 526058
rect 111098 526002 111154 526058
rect 111222 526002 111278 526058
rect 111346 526002 111402 526058
rect 111470 526002 111526 526058
rect 111594 526002 111650 526058
rect 111718 526002 111774 526058
rect 111842 526002 111898 526058
rect 111966 526002 112022 526058
rect 112090 526002 112146 526058
rect 112214 526002 112270 526058
rect 112338 526002 112394 526058
rect 112462 526002 112518 526058
rect 112586 526002 112642 526058
rect 112710 526002 112766 526058
rect 112834 526002 112890 526058
rect 112958 526002 113014 526058
rect 113082 526002 113138 526058
rect 113206 526002 113262 526058
rect 113330 526002 113386 526058
rect 113454 526002 113510 526058
rect 113578 526002 113634 526058
rect 113702 526002 113758 526058
rect 113826 526002 113882 526058
rect 113950 526002 114006 526058
rect 114074 526002 114130 526058
rect 114198 526002 114254 526058
rect 114322 526002 114378 526058
rect 114446 526002 114502 526058
rect 114570 526002 114626 526058
rect 114694 526002 114750 526058
rect 114818 526002 114874 526058
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 60202 514356 60258 514412
rect 60326 514356 60382 514412
rect 60450 514356 60506 514412
rect 60202 514232 60258 514288
rect 60326 514232 60382 514288
rect 60450 514232 60506 514288
rect 60202 514108 60258 514164
rect 60326 514108 60382 514164
rect 60450 514108 60506 514164
rect 60202 513984 60258 514040
rect 60326 513984 60382 514040
rect 60450 513984 60506 514040
rect 60202 513860 60258 513916
rect 60326 513860 60382 513916
rect 60450 513860 60506 513916
rect 60574 514356 60630 514412
rect 60698 514356 60754 514412
rect 60822 514356 60878 514412
rect 60946 514356 61002 514412
rect 60574 514232 60630 514288
rect 60698 514232 60754 514288
rect 60822 514232 60878 514288
rect 60946 514232 61002 514288
rect 60574 514108 60630 514164
rect 60698 514108 60754 514164
rect 60822 514108 60878 514164
rect 60946 514108 61002 514164
rect 60574 513984 60630 514040
rect 60698 513984 60754 514040
rect 60822 513984 60878 514040
rect 60946 513984 61002 514040
rect 60574 513860 60630 513916
rect 60698 513860 60754 513916
rect 60822 513860 60878 513916
rect 60946 513860 61002 513916
rect 61070 514356 61126 514412
rect 61194 514356 61250 514412
rect 61318 514356 61374 514412
rect 61442 514356 61498 514412
rect 61070 514232 61126 514288
rect 61194 514232 61250 514288
rect 61318 514232 61374 514288
rect 61442 514232 61498 514288
rect 61070 514108 61126 514164
rect 61194 514108 61250 514164
rect 61318 514108 61374 514164
rect 61442 514108 61498 514164
rect 61070 513984 61126 514040
rect 61194 513984 61250 514040
rect 61318 513984 61374 514040
rect 61442 513984 61498 514040
rect 61070 513860 61126 513916
rect 61194 513860 61250 513916
rect 61318 513860 61374 513916
rect 61442 513860 61498 513916
rect 61566 514356 61622 514412
rect 61690 514356 61746 514412
rect 61814 514356 61870 514412
rect 61938 514356 61994 514412
rect 61566 514232 61622 514288
rect 61690 514232 61746 514288
rect 61814 514232 61870 514288
rect 61938 514232 61994 514288
rect 61566 514108 61622 514164
rect 61690 514108 61746 514164
rect 61814 514108 61870 514164
rect 61938 514108 61994 514164
rect 61566 513984 61622 514040
rect 61690 513984 61746 514040
rect 61814 513984 61870 514040
rect 61938 513984 61994 514040
rect 61566 513860 61622 513916
rect 61690 513860 61746 513916
rect 61814 513860 61870 513916
rect 61938 513860 61994 513916
rect 62062 514356 62118 514412
rect 62186 514356 62242 514412
rect 62310 514356 62366 514412
rect 62434 514356 62490 514412
rect 62062 514232 62118 514288
rect 62186 514232 62242 514288
rect 62310 514232 62366 514288
rect 62434 514232 62490 514288
rect 62062 514108 62118 514164
rect 62186 514108 62242 514164
rect 62310 514108 62366 514164
rect 62434 514108 62490 514164
rect 62062 513984 62118 514040
rect 62186 513984 62242 514040
rect 62310 513984 62366 514040
rect 62434 513984 62490 514040
rect 62062 513860 62118 513916
rect 62186 513860 62242 513916
rect 62310 513860 62366 513916
rect 62434 513860 62490 513916
rect 62558 514356 62614 514412
rect 62682 514356 62738 514412
rect 62806 514356 62862 514412
rect 62930 514356 62986 514412
rect 62558 514232 62614 514288
rect 62682 514232 62738 514288
rect 62806 514232 62862 514288
rect 62930 514232 62986 514288
rect 62558 514108 62614 514164
rect 62682 514108 62738 514164
rect 62806 514108 62862 514164
rect 62930 514108 62986 514164
rect 62558 513984 62614 514040
rect 62682 513984 62738 514040
rect 62806 513984 62862 514040
rect 62930 513984 62986 514040
rect 62558 513860 62614 513916
rect 62682 513860 62738 513916
rect 62806 513860 62862 513916
rect 62930 513860 62986 513916
rect 63054 514356 63110 514412
rect 63178 514356 63234 514412
rect 63302 514356 63358 514412
rect 63426 514356 63482 514412
rect 63054 514232 63110 514288
rect 63178 514232 63234 514288
rect 63302 514232 63358 514288
rect 63426 514232 63482 514288
rect 63054 514108 63110 514164
rect 63178 514108 63234 514164
rect 63302 514108 63358 514164
rect 63426 514108 63482 514164
rect 63054 513984 63110 514040
rect 63178 513984 63234 514040
rect 63302 513984 63358 514040
rect 63426 513984 63482 514040
rect 63054 513860 63110 513916
rect 63178 513860 63234 513916
rect 63302 513860 63358 513916
rect 63426 513860 63482 513916
rect 63550 514356 63606 514412
rect 63674 514356 63730 514412
rect 63798 514356 63854 514412
rect 63922 514356 63978 514412
rect 63550 514232 63606 514288
rect 63674 514232 63730 514288
rect 63798 514232 63854 514288
rect 63922 514232 63978 514288
rect 63550 514108 63606 514164
rect 63674 514108 63730 514164
rect 63798 514108 63854 514164
rect 63922 514108 63978 514164
rect 63550 513984 63606 514040
rect 63674 513984 63730 514040
rect 63798 513984 63854 514040
rect 63922 513984 63978 514040
rect 63550 513860 63606 513916
rect 63674 513860 63730 513916
rect 63798 513860 63854 513916
rect 63922 513860 63978 513916
rect 64046 514356 64102 514412
rect 64170 514356 64226 514412
rect 64294 514356 64350 514412
rect 64418 514356 64474 514412
rect 64046 514232 64102 514288
rect 64170 514232 64226 514288
rect 64294 514232 64350 514288
rect 64418 514232 64474 514288
rect 64046 514108 64102 514164
rect 64170 514108 64226 514164
rect 64294 514108 64350 514164
rect 64418 514108 64474 514164
rect 64046 513984 64102 514040
rect 64170 513984 64226 514040
rect 64294 513984 64350 514040
rect 64418 513984 64474 514040
rect 64046 513860 64102 513916
rect 64170 513860 64226 513916
rect 64294 513860 64350 513916
rect 64418 513860 64474 513916
rect 64542 514356 64598 514412
rect 64666 514356 64722 514412
rect 64790 514356 64846 514412
rect 64914 514356 64970 514412
rect 64542 514232 64598 514288
rect 64666 514232 64722 514288
rect 64790 514232 64846 514288
rect 64914 514232 64970 514288
rect 64542 514108 64598 514164
rect 64666 514108 64722 514164
rect 64790 514108 64846 514164
rect 64914 514108 64970 514164
rect 64542 513984 64598 514040
rect 64666 513984 64722 514040
rect 64790 513984 64846 514040
rect 64914 513984 64970 514040
rect 64542 513860 64598 513916
rect 64666 513860 64722 513916
rect 64790 513860 64846 513916
rect 64914 513860 64970 513916
rect 65038 514356 65094 514412
rect 65162 514356 65218 514412
rect 65286 514356 65342 514412
rect 65410 514356 65466 514412
rect 65038 514232 65094 514288
rect 65162 514232 65218 514288
rect 65286 514232 65342 514288
rect 65410 514232 65466 514288
rect 65038 514108 65094 514164
rect 65162 514108 65218 514164
rect 65286 514108 65342 514164
rect 65410 514108 65466 514164
rect 65038 513984 65094 514040
rect 65162 513984 65218 514040
rect 65286 513984 65342 514040
rect 65410 513984 65466 514040
rect 65038 513860 65094 513916
rect 65162 513860 65218 513916
rect 65286 513860 65342 513916
rect 65410 513860 65466 513916
rect 65534 514356 65590 514412
rect 65658 514356 65714 514412
rect 65782 514356 65838 514412
rect 65906 514356 65962 514412
rect 65534 514232 65590 514288
rect 65658 514232 65714 514288
rect 65782 514232 65838 514288
rect 65906 514232 65962 514288
rect 65534 514108 65590 514164
rect 65658 514108 65714 514164
rect 65782 514108 65838 514164
rect 65906 514108 65962 514164
rect 65534 513984 65590 514040
rect 65658 513984 65714 514040
rect 65782 513984 65838 514040
rect 65906 513984 65962 514040
rect 65534 513860 65590 513916
rect 65658 513860 65714 513916
rect 65782 513860 65838 513916
rect 65906 513860 65962 513916
rect 66030 514356 66086 514412
rect 66154 514356 66210 514412
rect 66278 514356 66334 514412
rect 66402 514356 66458 514412
rect 66030 514232 66086 514288
rect 66154 514232 66210 514288
rect 66278 514232 66334 514288
rect 66402 514232 66458 514288
rect 66030 514108 66086 514164
rect 66154 514108 66210 514164
rect 66278 514108 66334 514164
rect 66402 514108 66458 514164
rect 66030 513984 66086 514040
rect 66154 513984 66210 514040
rect 66278 513984 66334 514040
rect 66402 513984 66458 514040
rect 66030 513860 66086 513916
rect 66154 513860 66210 513916
rect 66278 513860 66334 513916
rect 66402 513860 66458 513916
rect 90112 508379 90168 508435
rect 90236 508379 90292 508435
rect 90360 508379 90416 508435
rect 90484 508379 90540 508435
rect 90608 508379 90664 508435
rect 90732 508379 90788 508435
rect 90856 508379 90912 508435
rect 90980 508379 91036 508435
rect 91104 508379 91160 508435
rect 91228 508379 91284 508435
rect 91352 508379 91408 508435
rect 91476 508379 91532 508435
rect 91600 508379 91656 508435
rect 91724 508379 91780 508435
rect 91848 508379 91904 508435
rect 91972 508379 92028 508435
rect 92096 508379 92152 508435
rect 92220 508379 92276 508435
rect 92344 508379 92400 508435
rect 92468 508379 92524 508435
rect 92592 508379 92648 508435
rect 92716 508379 92772 508435
rect 92840 508379 92896 508435
rect 92964 508379 93020 508435
rect 93088 508379 93144 508435
rect 93212 508379 93268 508435
rect 93336 508379 93392 508435
rect 93460 508379 93516 508435
rect 93584 508379 93640 508435
rect 93708 508379 93764 508435
rect 93832 508379 93888 508435
rect 93956 508379 94012 508435
rect 94080 508379 94136 508435
rect 94204 508379 94260 508435
rect 94328 508379 94384 508435
rect 94452 508379 94508 508435
rect 94576 508379 94632 508435
rect 94700 508379 94756 508435
rect 94824 508379 94880 508435
rect 94948 508379 95004 508435
rect 95072 508379 95128 508435
rect 95196 508379 95252 508435
rect 95320 508379 95376 508435
rect 95444 508379 95500 508435
rect 95568 508379 95624 508435
rect 95692 508379 95748 508435
rect 95816 508379 95872 508435
rect 95940 508379 95996 508435
rect 96064 508379 96120 508435
rect 96188 508379 96244 508435
rect 96312 508379 96368 508435
rect 96436 508379 96492 508435
rect 96560 508379 96616 508435
rect 96684 508379 96740 508435
rect 96808 508379 96864 508435
rect 96932 508379 96988 508435
rect 97056 508379 97112 508435
rect 97180 508379 97236 508435
rect 97304 508379 97360 508435
rect 97428 508379 97484 508435
rect 97552 508379 97608 508435
rect 97676 508379 97732 508435
rect 97800 508379 97856 508435
rect 97924 508379 97980 508435
rect 98048 508379 98104 508435
rect 98172 508379 98228 508435
rect 98296 508379 98352 508435
rect 98420 508379 98476 508435
rect 98544 508379 98600 508435
rect 98668 508379 98724 508435
rect 98792 508379 98848 508435
rect 98916 508379 98972 508435
rect 99040 508379 99096 508435
rect 99164 508379 99220 508435
rect 99288 508379 99344 508435
rect 99412 508379 99468 508435
rect 99536 508379 99592 508435
rect 99660 508379 99716 508435
rect 99784 508379 99840 508435
rect 99908 508379 99964 508435
rect 100032 508379 100088 508435
rect 90112 508255 90168 508311
rect 90236 508255 90292 508311
rect 90360 508255 90416 508311
rect 90484 508255 90540 508311
rect 90608 508255 90664 508311
rect 90732 508255 90788 508311
rect 90856 508255 90912 508311
rect 90980 508255 91036 508311
rect 91104 508255 91160 508311
rect 91228 508255 91284 508311
rect 91352 508255 91408 508311
rect 91476 508255 91532 508311
rect 91600 508255 91656 508311
rect 91724 508255 91780 508311
rect 91848 508255 91904 508311
rect 91972 508255 92028 508311
rect 92096 508255 92152 508311
rect 92220 508255 92276 508311
rect 92344 508255 92400 508311
rect 92468 508255 92524 508311
rect 92592 508255 92648 508311
rect 92716 508255 92772 508311
rect 92840 508255 92896 508311
rect 92964 508255 93020 508311
rect 93088 508255 93144 508311
rect 93212 508255 93268 508311
rect 93336 508255 93392 508311
rect 93460 508255 93516 508311
rect 93584 508255 93640 508311
rect 93708 508255 93764 508311
rect 93832 508255 93888 508311
rect 93956 508255 94012 508311
rect 94080 508255 94136 508311
rect 94204 508255 94260 508311
rect 94328 508255 94384 508311
rect 94452 508255 94508 508311
rect 94576 508255 94632 508311
rect 94700 508255 94756 508311
rect 94824 508255 94880 508311
rect 94948 508255 95004 508311
rect 95072 508255 95128 508311
rect 95196 508255 95252 508311
rect 95320 508255 95376 508311
rect 95444 508255 95500 508311
rect 95568 508255 95624 508311
rect 95692 508255 95748 508311
rect 95816 508255 95872 508311
rect 95940 508255 95996 508311
rect 96064 508255 96120 508311
rect 96188 508255 96244 508311
rect 96312 508255 96368 508311
rect 96436 508255 96492 508311
rect 96560 508255 96616 508311
rect 96684 508255 96740 508311
rect 96808 508255 96864 508311
rect 96932 508255 96988 508311
rect 97056 508255 97112 508311
rect 97180 508255 97236 508311
rect 97304 508255 97360 508311
rect 97428 508255 97484 508311
rect 97552 508255 97608 508311
rect 97676 508255 97732 508311
rect 97800 508255 97856 508311
rect 97924 508255 97980 508311
rect 98048 508255 98104 508311
rect 98172 508255 98228 508311
rect 98296 508255 98352 508311
rect 98420 508255 98476 508311
rect 98544 508255 98600 508311
rect 98668 508255 98724 508311
rect 98792 508255 98848 508311
rect 98916 508255 98972 508311
rect 99040 508255 99096 508311
rect 99164 508255 99220 508311
rect 99288 508255 99344 508311
rect 99412 508255 99468 508311
rect 99536 508255 99592 508311
rect 99660 508255 99716 508311
rect 99784 508255 99840 508311
rect 99908 508255 99964 508311
rect 100032 508255 100088 508311
rect 90112 508131 90168 508187
rect 90236 508131 90292 508187
rect 90360 508131 90416 508187
rect 90484 508131 90540 508187
rect 90608 508131 90664 508187
rect 90732 508131 90788 508187
rect 90856 508131 90912 508187
rect 90980 508131 91036 508187
rect 91104 508131 91160 508187
rect 91228 508131 91284 508187
rect 91352 508131 91408 508187
rect 91476 508131 91532 508187
rect 91600 508131 91656 508187
rect 91724 508131 91780 508187
rect 91848 508131 91904 508187
rect 91972 508131 92028 508187
rect 92096 508131 92152 508187
rect 92220 508131 92276 508187
rect 92344 508131 92400 508187
rect 92468 508131 92524 508187
rect 92592 508131 92648 508187
rect 92716 508131 92772 508187
rect 92840 508131 92896 508187
rect 92964 508131 93020 508187
rect 93088 508131 93144 508187
rect 93212 508131 93268 508187
rect 93336 508131 93392 508187
rect 93460 508131 93516 508187
rect 93584 508131 93640 508187
rect 93708 508131 93764 508187
rect 93832 508131 93888 508187
rect 93956 508131 94012 508187
rect 94080 508131 94136 508187
rect 94204 508131 94260 508187
rect 94328 508131 94384 508187
rect 94452 508131 94508 508187
rect 94576 508131 94632 508187
rect 94700 508131 94756 508187
rect 94824 508131 94880 508187
rect 94948 508131 95004 508187
rect 95072 508131 95128 508187
rect 95196 508131 95252 508187
rect 95320 508131 95376 508187
rect 95444 508131 95500 508187
rect 95568 508131 95624 508187
rect 95692 508131 95748 508187
rect 95816 508131 95872 508187
rect 95940 508131 95996 508187
rect 96064 508131 96120 508187
rect 96188 508131 96244 508187
rect 96312 508131 96368 508187
rect 96436 508131 96492 508187
rect 96560 508131 96616 508187
rect 96684 508131 96740 508187
rect 96808 508131 96864 508187
rect 96932 508131 96988 508187
rect 97056 508131 97112 508187
rect 97180 508131 97236 508187
rect 97304 508131 97360 508187
rect 97428 508131 97484 508187
rect 97552 508131 97608 508187
rect 97676 508131 97732 508187
rect 97800 508131 97856 508187
rect 97924 508131 97980 508187
rect 98048 508131 98104 508187
rect 98172 508131 98228 508187
rect 98296 508131 98352 508187
rect 98420 508131 98476 508187
rect 98544 508131 98600 508187
rect 98668 508131 98724 508187
rect 98792 508131 98848 508187
rect 98916 508131 98972 508187
rect 99040 508131 99096 508187
rect 99164 508131 99220 508187
rect 99288 508131 99344 508187
rect 99412 508131 99468 508187
rect 99536 508131 99592 508187
rect 99660 508131 99716 508187
rect 99784 508131 99840 508187
rect 99908 508131 99964 508187
rect 100032 508131 100088 508187
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 89904 507855 89960 507911
rect 90028 507855 90084 507911
rect 90152 507855 90208 507911
rect 90276 507855 90332 507911
rect 90400 507855 90456 507911
rect 90524 507855 90580 507911
rect 90648 507855 90704 507911
rect 90772 507855 90828 507911
rect 90896 507855 90952 507911
rect 91020 507855 91076 507911
rect 91144 507855 91200 507911
rect 91268 507855 91324 507911
rect 91392 507855 91448 507911
rect 91516 507855 91572 507911
rect 91640 507855 91696 507911
rect 91764 507855 91820 507911
rect 91888 507855 91944 507911
rect 92012 507855 92068 507911
rect 92136 507855 92192 507911
rect 92260 507855 92316 507911
rect 92384 507855 92440 507911
rect 92508 507855 92564 507911
rect 92632 507855 92688 507911
rect 92756 507855 92812 507911
rect 92880 507855 92936 507911
rect 93004 507855 93060 507911
rect 93128 507855 93184 507911
rect 93252 507855 93308 507911
rect 93376 507855 93432 507911
rect 93500 507855 93556 507911
rect 93624 507855 93680 507911
rect 93748 507855 93804 507911
rect 93872 507855 93928 507911
rect 93996 507855 94052 507911
rect 94120 507855 94176 507911
rect 94244 507855 94300 507911
rect 94368 507855 94424 507911
rect 94492 507855 94548 507911
rect 94616 507855 94672 507911
rect 94740 507855 94796 507911
rect 94864 507855 94920 507911
rect 94988 507855 95044 507911
rect 95112 507855 95168 507911
rect 95236 507855 95292 507911
rect 95360 507855 95416 507911
rect 95484 507855 95540 507911
rect 95608 507855 95664 507911
rect 95732 507855 95788 507911
rect 95856 507855 95912 507911
rect 95980 507855 96036 507911
rect 96104 507855 96160 507911
rect 96228 507855 96284 507911
rect 96352 507855 96408 507911
rect 96476 507855 96532 507911
rect 96600 507855 96656 507911
rect 96724 507855 96780 507911
rect 96848 507855 96904 507911
rect 96972 507855 97028 507911
rect 97096 507855 97152 507911
rect 97220 507855 97276 507911
rect 97344 507855 97400 507911
rect 97468 507855 97524 507911
rect 97592 507855 97648 507911
rect 97716 507855 97772 507911
rect 97840 507855 97896 507911
rect 97964 507855 98020 507911
rect 98088 507855 98144 507911
rect 98212 507855 98268 507911
rect 98336 507855 98392 507911
rect 98460 507855 98516 507911
rect 98584 507855 98640 507911
rect 98708 507855 98764 507911
rect 98832 507855 98888 507911
rect 98956 507855 99012 507911
rect 99080 507855 99136 507911
rect 99204 507855 99260 507911
rect 99328 507855 99384 507911
rect 99452 507855 99508 507911
rect 99576 507855 99632 507911
rect 99700 507855 99756 507911
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 63430 496156 63486 496212
rect 63430 496032 63486 496088
rect 63430 495908 63486 495964
rect 63554 496156 63610 496212
rect 63678 496156 63734 496212
rect 63802 496156 63858 496212
rect 63926 496156 63982 496212
rect 63554 496032 63610 496088
rect 63678 496032 63734 496088
rect 63802 496032 63858 496088
rect 63926 496032 63982 496088
rect 63554 495908 63610 495964
rect 63678 495908 63734 495964
rect 63802 495908 63858 495964
rect 63926 495908 63982 495964
rect 64050 496156 64106 496212
rect 64174 496156 64230 496212
rect 64298 496156 64354 496212
rect 64422 496156 64478 496212
rect 64050 496032 64106 496088
rect 64174 496032 64230 496088
rect 64298 496032 64354 496088
rect 64422 496032 64478 496088
rect 64050 495908 64106 495964
rect 64174 495908 64230 495964
rect 64298 495908 64354 495964
rect 64422 495908 64478 495964
rect 64546 496156 64602 496212
rect 64670 496156 64726 496212
rect 64794 496156 64850 496212
rect 64918 496156 64974 496212
rect 64546 496032 64602 496088
rect 64670 496032 64726 496088
rect 64794 496032 64850 496088
rect 64918 496032 64974 496088
rect 64546 495908 64602 495964
rect 64670 495908 64726 495964
rect 64794 495908 64850 495964
rect 64918 495908 64974 495964
rect 65042 496156 65098 496212
rect 65166 496156 65222 496212
rect 65290 496156 65346 496212
rect 65414 496156 65470 496212
rect 65042 496032 65098 496088
rect 65166 496032 65222 496088
rect 65290 496032 65346 496088
rect 65414 496032 65470 496088
rect 65042 495908 65098 495964
rect 65166 495908 65222 495964
rect 65290 495908 65346 495964
rect 65414 495908 65470 495964
rect 65538 496156 65594 496212
rect 65662 496156 65718 496212
rect 65786 496156 65842 496212
rect 65910 496156 65966 496212
rect 65538 496032 65594 496088
rect 65662 496032 65718 496088
rect 65786 496032 65842 496088
rect 65910 496032 65966 496088
rect 65538 495908 65594 495964
rect 65662 495908 65718 495964
rect 65786 495908 65842 495964
rect 65910 495908 65966 495964
rect 66034 496156 66090 496212
rect 66158 496156 66214 496212
rect 66282 496156 66338 496212
rect 66406 496156 66462 496212
rect 66034 496032 66090 496088
rect 66158 496032 66214 496088
rect 66282 496032 66338 496088
rect 66406 496032 66462 496088
rect 66034 495908 66090 495964
rect 66158 495908 66214 495964
rect 66282 495908 66338 495964
rect 66406 495908 66462 495964
rect 66530 496156 66586 496212
rect 66654 496156 66710 496212
rect 66778 496156 66834 496212
rect 66902 496156 66958 496212
rect 66530 496032 66586 496088
rect 66654 496032 66710 496088
rect 66778 496032 66834 496088
rect 66902 496032 66958 496088
rect 66530 495908 66586 495964
rect 66654 495908 66710 495964
rect 66778 495908 66834 495964
rect 66902 495908 66958 495964
rect 67026 496156 67082 496212
rect 67150 496156 67206 496212
rect 67274 496156 67330 496212
rect 67398 496156 67454 496212
rect 67026 496032 67082 496088
rect 67150 496032 67206 496088
rect 67274 496032 67330 496088
rect 67398 496032 67454 496088
rect 67026 495908 67082 495964
rect 67150 495908 67206 495964
rect 67274 495908 67330 495964
rect 67398 495908 67454 495964
rect 67522 496156 67578 496212
rect 67646 496156 67702 496212
rect 67770 496156 67826 496212
rect 67894 496156 67950 496212
rect 67522 496032 67578 496088
rect 67646 496032 67702 496088
rect 67770 496032 67826 496088
rect 67894 496032 67950 496088
rect 67522 495908 67578 495964
rect 67646 495908 67702 495964
rect 67770 495908 67826 495964
rect 67894 495908 67950 495964
rect 68018 496156 68074 496212
rect 68142 496156 68198 496212
rect 68266 496156 68322 496212
rect 68390 496156 68446 496212
rect 68018 496032 68074 496088
rect 68142 496032 68198 496088
rect 68266 496032 68322 496088
rect 68390 496032 68446 496088
rect 68018 495908 68074 495964
rect 68142 495908 68198 495964
rect 68266 495908 68322 495964
rect 68390 495908 68446 495964
rect 68514 496156 68570 496212
rect 68638 496156 68694 496212
rect 68762 496156 68818 496212
rect 68886 496156 68942 496212
rect 68514 496032 68570 496088
rect 68638 496032 68694 496088
rect 68762 496032 68818 496088
rect 68886 496032 68942 496088
rect 68514 495908 68570 495964
rect 68638 495908 68694 495964
rect 68762 495908 68818 495964
rect 68886 495908 68942 495964
rect 69010 496156 69066 496212
rect 69134 496156 69190 496212
rect 69258 496156 69314 496212
rect 69382 496156 69438 496212
rect 69010 496032 69066 496088
rect 69134 496032 69190 496088
rect 69258 496032 69314 496088
rect 69382 496032 69438 496088
rect 69010 495908 69066 495964
rect 69134 495908 69190 495964
rect 69258 495908 69314 495964
rect 69382 495908 69438 495964
rect 69506 496156 69562 496212
rect 69630 496156 69686 496212
rect 69754 496156 69810 496212
rect 69878 496156 69934 496212
rect 69506 496032 69562 496088
rect 69630 496032 69686 496088
rect 69754 496032 69810 496088
rect 69878 496032 69934 496088
rect 69506 495908 69562 495964
rect 69630 495908 69686 495964
rect 69754 495908 69810 495964
rect 69878 495908 69934 495964
rect 70002 496156 70058 496212
rect 70126 496156 70182 496212
rect 70250 496156 70306 496212
rect 70374 496156 70430 496212
rect 70002 496032 70058 496088
rect 70126 496032 70182 496088
rect 70250 496032 70306 496088
rect 70374 496032 70430 496088
rect 70002 495908 70058 495964
rect 70126 495908 70182 495964
rect 70250 495908 70306 495964
rect 70374 495908 70430 495964
rect 85236 490216 85292 490272
rect 85360 490216 85416 490272
rect 85484 490216 85540 490272
rect 85608 490216 85664 490272
rect 85732 490216 85788 490272
rect 85856 490216 85912 490272
rect 85980 490216 86036 490272
rect 86104 490216 86160 490272
rect 86228 490216 86284 490272
rect 86352 490216 86408 490272
rect 86476 490216 86532 490272
rect 86600 490216 86656 490272
rect 86724 490216 86780 490272
rect 86848 490216 86904 490272
rect 86972 490216 87028 490272
rect 87096 490216 87152 490272
rect 87220 490216 87276 490272
rect 87344 490216 87400 490272
rect 87468 490216 87524 490272
rect 87592 490216 87648 490272
rect 87716 490216 87772 490272
rect 87840 490216 87896 490272
rect 87964 490216 88020 490272
rect 88088 490216 88144 490272
rect 88212 490216 88268 490272
rect 88336 490216 88392 490272
rect 88460 490216 88516 490272
rect 88584 490216 88640 490272
rect 88708 490216 88764 490272
rect 85236 490092 85292 490148
rect 85360 490092 85416 490148
rect 85484 490092 85540 490148
rect 85608 490092 85664 490148
rect 85732 490092 85788 490148
rect 85856 490092 85912 490148
rect 85980 490092 86036 490148
rect 86104 490092 86160 490148
rect 86228 490092 86284 490148
rect 86352 490092 86408 490148
rect 86476 490092 86532 490148
rect 86600 490092 86656 490148
rect 86724 490092 86780 490148
rect 86848 490092 86904 490148
rect 86972 490092 87028 490148
rect 87096 490092 87152 490148
rect 87220 490092 87276 490148
rect 87344 490092 87400 490148
rect 87468 490092 87524 490148
rect 87592 490092 87648 490148
rect 87716 490092 87772 490148
rect 87840 490092 87896 490148
rect 87964 490092 88020 490148
rect 88088 490092 88144 490148
rect 88212 490092 88268 490148
rect 88336 490092 88392 490148
rect 88460 490092 88516 490148
rect 88584 490092 88640 490148
rect 88708 490092 88764 490148
rect 85236 489968 85292 490024
rect 85360 489968 85416 490024
rect 85484 489968 85540 490024
rect 85608 489968 85664 490024
rect 85732 489968 85788 490024
rect 85856 489968 85912 490024
rect 85980 489968 86036 490024
rect 86104 489968 86160 490024
rect 86228 489968 86284 490024
rect 86352 489968 86408 490024
rect 86476 489968 86532 490024
rect 86600 489968 86656 490024
rect 86724 489968 86780 490024
rect 86848 489968 86904 490024
rect 86972 489968 87028 490024
rect 87096 489968 87152 490024
rect 87220 489968 87276 490024
rect 87344 489968 87400 490024
rect 87468 489968 87524 490024
rect 87592 489968 87648 490024
rect 87716 489968 87772 490024
rect 87840 489968 87896 490024
rect 87964 489968 88020 490024
rect 88088 489968 88144 490024
rect 88212 489968 88268 490024
rect 88336 489968 88392 490024
rect 88460 489968 88516 490024
rect 88584 489968 88640 490024
rect 88708 489968 88764 490024
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 57932 403982 57988 404038
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 80936 478302 80992 478358
rect 81060 478302 81116 478358
rect 81184 478302 81240 478358
rect 81308 478302 81364 478358
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 66574 406294 66630 406350
rect 66698 406294 66754 406350
rect 66574 406170 66630 406226
rect 66698 406170 66754 406226
rect 66574 406046 66630 406102
rect 66698 406046 66754 406102
rect 66574 405922 66630 405978
rect 66698 405922 66754 405978
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 97674 418294 97730 418350
rect 97798 418294 97854 418350
rect 97922 418294 97978 418350
rect 98046 418294 98102 418350
rect 97674 418170 97730 418226
rect 97798 418170 97854 418226
rect 97922 418170 97978 418226
rect 98046 418170 98102 418226
rect 97674 418046 97730 418102
rect 97798 418046 97854 418102
rect 97922 418046 97978 418102
rect 98046 418046 98102 418102
rect 97674 417922 97730 417978
rect 97798 417922 97854 417978
rect 97922 417922 97978 417978
rect 98046 417922 98102 417978
rect 83916 416762 83972 416818
rect 70674 406294 70730 406350
rect 70798 406294 70854 406350
rect 70922 406294 70978 406350
rect 71046 406294 71102 406350
rect 70674 406170 70730 406226
rect 70798 406170 70854 406226
rect 70922 406170 70978 406226
rect 71046 406170 71102 406226
rect 70674 406046 70730 406102
rect 70798 406046 70854 406102
rect 70922 406046 70978 406102
rect 71046 406046 71102 406102
rect 70674 405922 70730 405978
rect 70798 405922 70854 405978
rect 70922 405922 70978 405978
rect 71046 405922 71102 405978
rect 71894 406294 71950 406350
rect 72018 406294 72074 406350
rect 71894 406170 71950 406226
rect 72018 406170 72074 406226
rect 71894 406046 71950 406102
rect 72018 406046 72074 406102
rect 71894 405922 71950 405978
rect 72018 405922 72074 405978
rect 77214 406294 77270 406350
rect 77338 406294 77394 406350
rect 77214 406170 77270 406226
rect 77338 406170 77394 406226
rect 77214 406046 77270 406102
rect 77338 406046 77394 406102
rect 77214 405922 77270 405978
rect 77338 405922 77394 405978
rect 82534 406294 82590 406350
rect 82658 406294 82714 406350
rect 82534 406170 82590 406226
rect 82658 406170 82714 406226
rect 82534 406046 82590 406102
rect 82658 406046 82714 406102
rect 82534 405922 82590 405978
rect 82658 405922 82714 405978
rect 63914 400294 63970 400350
rect 64038 400294 64094 400350
rect 63914 400170 63970 400226
rect 64038 400170 64094 400226
rect 63914 400046 63970 400102
rect 64038 400046 64094 400102
rect 63914 399922 63970 399978
rect 64038 399922 64094 399978
rect 69234 400294 69290 400350
rect 69358 400294 69414 400350
rect 69234 400170 69290 400226
rect 69358 400170 69414 400226
rect 74554 400294 74610 400350
rect 74678 400294 74734 400350
rect 74554 400170 74610 400226
rect 74678 400170 74734 400226
rect 69234 400046 69290 400102
rect 69358 400046 69414 400102
rect 69234 399922 69290 399978
rect 69358 399922 69414 399978
rect 62076 395522 62132 395578
rect 39954 388294 40010 388350
rect 40078 388294 40134 388350
rect 40202 388294 40258 388350
rect 40326 388294 40382 388350
rect 39954 388170 40010 388226
rect 40078 388170 40134 388226
rect 40202 388170 40258 388226
rect 40326 388170 40382 388226
rect 39954 388046 40010 388102
rect 40078 388046 40134 388102
rect 40202 388046 40258 388102
rect 40326 388046 40382 388102
rect 39954 387922 40010 387978
rect 40078 387922 40134 387978
rect 40202 387922 40258 387978
rect 40326 387922 40382 387978
rect 39954 370294 40010 370350
rect 40078 370294 40134 370350
rect 40202 370294 40258 370350
rect 40326 370294 40382 370350
rect 39954 370170 40010 370226
rect 40078 370170 40134 370226
rect 40202 370170 40258 370226
rect 40326 370170 40382 370226
rect 39954 370046 40010 370102
rect 40078 370046 40134 370102
rect 40202 370046 40258 370102
rect 40326 370046 40382 370102
rect 39954 369922 40010 369978
rect 40078 369922 40134 369978
rect 40202 369922 40258 369978
rect 40326 369922 40382 369978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 39954 352294 40010 352350
rect 40078 352294 40134 352350
rect 40202 352294 40258 352350
rect 40326 352294 40382 352350
rect 39954 352170 40010 352226
rect 40078 352170 40134 352226
rect 40202 352170 40258 352226
rect 40326 352170 40382 352226
rect 39954 352046 40010 352102
rect 40078 352046 40134 352102
rect 40202 352046 40258 352102
rect 40326 352046 40382 352102
rect 39954 351922 40010 351978
rect 40078 351922 40134 351978
rect 40202 351922 40258 351978
rect 40326 351922 40382 351978
rect 64878 352294 64934 352350
rect 65002 352294 65058 352350
rect 64878 352170 64934 352226
rect 65002 352170 65058 352226
rect 64878 352046 64934 352102
rect 65002 352046 65058 352102
rect 64878 351922 64934 351978
rect 65002 351922 65058 351978
rect 74554 400046 74610 400102
rect 74678 400046 74734 400102
rect 74554 399922 74610 399978
rect 74678 399922 74734 399978
rect 79874 400294 79930 400350
rect 79998 400294 80054 400350
rect 79874 400170 79930 400226
rect 79998 400170 80054 400226
rect 79874 400046 79930 400102
rect 79998 400046 80054 400102
rect 79874 399922 79930 399978
rect 79998 399922 80054 399978
rect 97674 400294 97730 400350
rect 97798 400294 97854 400350
rect 97922 400294 97978 400350
rect 98046 400294 98102 400350
rect 97674 400170 97730 400226
rect 97798 400170 97854 400226
rect 97922 400170 97978 400226
rect 98046 400170 98102 400226
rect 97674 400046 97730 400102
rect 97798 400046 97854 400102
rect 97922 400046 97978 400102
rect 98046 400046 98102 400102
rect 97674 399922 97730 399978
rect 97798 399922 97854 399978
rect 97922 399922 97978 399978
rect 98046 399922 98102 399978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 70674 352294 70730 352350
rect 70798 352294 70854 352350
rect 70922 352294 70978 352350
rect 71046 352294 71102 352350
rect 70674 352170 70730 352226
rect 70798 352170 70854 352226
rect 70922 352170 70978 352226
rect 71046 352170 71102 352226
rect 70674 352046 70730 352102
rect 70798 352046 70854 352102
rect 70922 352046 70978 352102
rect 71046 352046 71102 352102
rect 70674 351922 70730 351978
rect 70798 351922 70854 351978
rect 70922 351922 70978 351978
rect 71046 351922 71102 351978
rect 49518 346294 49574 346350
rect 49642 346294 49698 346350
rect 49518 346170 49574 346226
rect 49642 346170 49698 346226
rect 49518 346046 49574 346102
rect 49642 346046 49698 346102
rect 49518 345922 49574 345978
rect 49642 345922 49698 345978
rect 80238 346294 80294 346350
rect 80362 346294 80418 346350
rect 80238 346170 80294 346226
rect 80362 346170 80418 346226
rect 80238 346046 80294 346102
rect 80362 346046 80418 346102
rect 80238 345922 80294 345978
rect 80362 345922 80418 345978
rect 39954 334294 40010 334350
rect 40078 334294 40134 334350
rect 40202 334294 40258 334350
rect 40326 334294 40382 334350
rect 39954 334170 40010 334226
rect 40078 334170 40134 334226
rect 40202 334170 40258 334226
rect 40326 334170 40382 334226
rect 39954 334046 40010 334102
rect 40078 334046 40134 334102
rect 40202 334046 40258 334102
rect 40326 334046 40382 334102
rect 39954 333922 40010 333978
rect 40078 333922 40134 333978
rect 40202 333922 40258 333978
rect 40326 333922 40382 333978
rect 64878 334294 64934 334350
rect 65002 334294 65058 334350
rect 64878 334170 64934 334226
rect 65002 334170 65058 334226
rect 64878 334046 64934 334102
rect 65002 334046 65058 334102
rect 64878 333922 64934 333978
rect 65002 333922 65058 333978
rect 49518 328294 49574 328350
rect 49642 328294 49698 328350
rect 49518 328170 49574 328226
rect 49642 328170 49698 328226
rect 49518 328046 49574 328102
rect 49642 328046 49698 328102
rect 49518 327922 49574 327978
rect 49642 327922 49698 327978
rect 66954 328294 67010 328350
rect 67078 328294 67134 328350
rect 67202 328294 67258 328350
rect 67326 328294 67382 328350
rect 66954 328170 67010 328226
rect 67078 328170 67134 328226
rect 67202 328170 67258 328226
rect 67326 328170 67382 328226
rect 66954 328046 67010 328102
rect 67078 328046 67134 328102
rect 67202 328046 67258 328102
rect 67326 328046 67382 328102
rect 66954 327922 67010 327978
rect 67078 327922 67134 327978
rect 67202 327922 67258 327978
rect 67326 327922 67382 327978
rect 39954 316294 40010 316350
rect 40078 316294 40134 316350
rect 40202 316294 40258 316350
rect 40326 316294 40382 316350
rect 39954 316170 40010 316226
rect 40078 316170 40134 316226
rect 40202 316170 40258 316226
rect 40326 316170 40382 316226
rect 39954 316046 40010 316102
rect 40078 316046 40134 316102
rect 40202 316046 40258 316102
rect 40326 316046 40382 316102
rect 39954 315922 40010 315978
rect 40078 315922 40134 315978
rect 40202 315922 40258 315978
rect 40326 315922 40382 315978
rect 39954 298294 40010 298350
rect 40078 298294 40134 298350
rect 40202 298294 40258 298350
rect 40326 298294 40382 298350
rect 39954 298170 40010 298226
rect 40078 298170 40134 298226
rect 40202 298170 40258 298226
rect 40326 298170 40382 298226
rect 39954 298046 40010 298102
rect 40078 298046 40134 298102
rect 40202 298046 40258 298102
rect 40326 298046 40382 298102
rect 39954 297922 40010 297978
rect 40078 297922 40134 297978
rect 40202 297922 40258 297978
rect 40326 297922 40382 297978
rect 66954 310294 67010 310350
rect 67078 310294 67134 310350
rect 67202 310294 67258 310350
rect 67326 310294 67382 310350
rect 66954 310170 67010 310226
rect 67078 310170 67134 310226
rect 67202 310170 67258 310226
rect 67326 310170 67382 310226
rect 66954 310046 67010 310102
rect 67078 310046 67134 310102
rect 67202 310046 67258 310102
rect 67326 310046 67382 310102
rect 66954 309922 67010 309978
rect 67078 309922 67134 309978
rect 67202 309922 67258 309978
rect 67326 309922 67382 309978
rect 66954 292294 67010 292350
rect 67078 292294 67134 292350
rect 67202 292294 67258 292350
rect 67326 292294 67382 292350
rect 66954 292170 67010 292226
rect 67078 292170 67134 292226
rect 67202 292170 67258 292226
rect 67326 292170 67382 292226
rect 66954 292046 67010 292102
rect 67078 292046 67134 292102
rect 67202 292046 67258 292102
rect 67326 292046 67382 292102
rect 66954 291922 67010 291978
rect 67078 291922 67134 291978
rect 67202 291922 67258 291978
rect 67326 291922 67382 291978
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 80238 328294 80294 328350
rect 80362 328294 80418 328350
rect 80238 328170 80294 328226
rect 80362 328170 80418 328226
rect 80238 328046 80294 328102
rect 80362 328046 80418 328102
rect 80238 327922 80294 327978
rect 80362 327922 80418 327978
rect 70674 316294 70730 316350
rect 70798 316294 70854 316350
rect 70922 316294 70978 316350
rect 71046 316294 71102 316350
rect 70674 316170 70730 316226
rect 70798 316170 70854 316226
rect 70922 316170 70978 316226
rect 71046 316170 71102 316226
rect 70674 316046 70730 316102
rect 70798 316046 70854 316102
rect 70922 316046 70978 316102
rect 71046 316046 71102 316102
rect 70674 315922 70730 315978
rect 70798 315922 70854 315978
rect 70922 315922 70978 315978
rect 71046 315922 71102 315978
rect 85596 305882 85652 305938
rect 70674 298294 70730 298350
rect 70798 298294 70854 298350
rect 70922 298294 70978 298350
rect 71046 298294 71102 298350
rect 70674 298170 70730 298226
rect 70798 298170 70854 298226
rect 70922 298170 70978 298226
rect 71046 298170 71102 298226
rect 70674 298046 70730 298102
rect 70798 298046 70854 298102
rect 70922 298046 70978 298102
rect 71046 298046 71102 298102
rect 70674 297922 70730 297978
rect 70798 297922 70854 297978
rect 70922 297922 70978 297978
rect 71046 297922 71102 297978
rect 72156 302462 72212 302518
rect 39954 280294 40010 280350
rect 40078 280294 40134 280350
rect 40202 280294 40258 280350
rect 40326 280294 40382 280350
rect 39954 280170 40010 280226
rect 40078 280170 40134 280226
rect 40202 280170 40258 280226
rect 40326 280170 40382 280226
rect 39954 280046 40010 280102
rect 40078 280046 40134 280102
rect 40202 280046 40258 280102
rect 40326 280046 40382 280102
rect 39954 279922 40010 279978
rect 40078 279922 40134 279978
rect 40202 279922 40258 279978
rect 40326 279922 40382 279978
rect 59878 280294 59934 280350
rect 60002 280294 60058 280350
rect 59878 280170 59934 280226
rect 60002 280170 60058 280226
rect 59878 280046 59934 280102
rect 60002 280046 60058 280102
rect 59878 279922 59934 279978
rect 60002 279922 60058 279978
rect 44518 274294 44574 274350
rect 44642 274294 44698 274350
rect 44518 274170 44574 274226
rect 44642 274170 44698 274226
rect 44518 274046 44574 274102
rect 44642 274046 44698 274102
rect 44518 273922 44574 273978
rect 44642 273922 44698 273978
rect 75238 274294 75294 274350
rect 75362 274294 75418 274350
rect 75238 274170 75294 274226
rect 75362 274170 75418 274226
rect 75238 274046 75294 274102
rect 75362 274046 75418 274102
rect 75238 273922 75294 273978
rect 75362 273922 75418 273978
rect 39954 262294 40010 262350
rect 40078 262294 40134 262350
rect 40202 262294 40258 262350
rect 40326 262294 40382 262350
rect 39954 262170 40010 262226
rect 40078 262170 40134 262226
rect 40202 262170 40258 262226
rect 40326 262170 40382 262226
rect 39954 262046 40010 262102
rect 40078 262046 40134 262102
rect 40202 262046 40258 262102
rect 40326 262046 40382 262102
rect 39954 261922 40010 261978
rect 40078 261922 40134 261978
rect 40202 261922 40258 261978
rect 40326 261922 40382 261978
rect 59878 262294 59934 262350
rect 60002 262294 60058 262350
rect 59878 262170 59934 262226
rect 60002 262170 60058 262226
rect 59878 262046 59934 262102
rect 60002 262046 60058 262102
rect 59878 261922 59934 261978
rect 60002 261922 60058 261978
rect 44518 256294 44574 256350
rect 44642 256294 44698 256350
rect 44518 256170 44574 256226
rect 44642 256170 44698 256226
rect 44518 256046 44574 256102
rect 44642 256046 44698 256102
rect 44518 255922 44574 255978
rect 44642 255922 44698 255978
rect 75238 256294 75294 256350
rect 75362 256294 75418 256350
rect 75238 256170 75294 256226
rect 75362 256170 75418 256226
rect 75238 256046 75294 256102
rect 75362 256046 75418 256102
rect 75238 255922 75294 255978
rect 75362 255922 75418 255978
rect 39954 244294 40010 244350
rect 40078 244294 40134 244350
rect 40202 244294 40258 244350
rect 40326 244294 40382 244350
rect 39954 244170 40010 244226
rect 40078 244170 40134 244226
rect 40202 244170 40258 244226
rect 40326 244170 40382 244226
rect 39954 244046 40010 244102
rect 40078 244046 40134 244102
rect 40202 244046 40258 244102
rect 40326 244046 40382 244102
rect 39954 243922 40010 243978
rect 40078 243922 40134 243978
rect 40202 243922 40258 243978
rect 40326 243922 40382 243978
rect 42812 247022 42868 247078
rect 59878 244294 59934 244350
rect 60002 244294 60058 244350
rect 59878 244170 59934 244226
rect 60002 244170 60058 244226
rect 59878 244046 59934 244102
rect 60002 244046 60058 244102
rect 59878 243922 59934 243978
rect 60002 243922 60058 243978
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 39954 226294 40010 226350
rect 40078 226294 40134 226350
rect 40202 226294 40258 226350
rect 40326 226294 40382 226350
rect 39954 226170 40010 226226
rect 40078 226170 40134 226226
rect 40202 226170 40258 226226
rect 40326 226170 40382 226226
rect 39954 226046 40010 226102
rect 40078 226046 40134 226102
rect 40202 226046 40258 226102
rect 40326 226046 40382 226102
rect 39954 225922 40010 225978
rect 40078 225922 40134 225978
rect 40202 225922 40258 225978
rect 40326 225922 40382 225978
rect 39954 208294 40010 208350
rect 40078 208294 40134 208350
rect 40202 208294 40258 208350
rect 40326 208294 40382 208350
rect 39954 208170 40010 208226
rect 40078 208170 40134 208226
rect 40202 208170 40258 208226
rect 40326 208170 40382 208226
rect 39954 208046 40010 208102
rect 40078 208046 40134 208102
rect 40202 208046 40258 208102
rect 40326 208046 40382 208102
rect 39954 207922 40010 207978
rect 40078 207922 40134 207978
rect 40202 207922 40258 207978
rect 40326 207922 40382 207978
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 39452 205802 39508 205858
rect 39954 190294 40010 190350
rect 40078 190294 40134 190350
rect 40202 190294 40258 190350
rect 40326 190294 40382 190350
rect 39954 190170 40010 190226
rect 40078 190170 40134 190226
rect 40202 190170 40258 190226
rect 40326 190170 40382 190226
rect 39954 190046 40010 190102
rect 40078 190046 40134 190102
rect 40202 190046 40258 190102
rect 40326 190046 40382 190102
rect 39954 189922 40010 189978
rect 40078 189922 40134 189978
rect 40202 189922 40258 189978
rect 40326 189922 40382 189978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 39954 136294 40010 136350
rect 40078 136294 40134 136350
rect 40202 136294 40258 136350
rect 40326 136294 40382 136350
rect 39954 136170 40010 136226
rect 40078 136170 40134 136226
rect 40202 136170 40258 136226
rect 40326 136170 40382 136226
rect 39954 136046 40010 136102
rect 40078 136046 40134 136102
rect 40202 136046 40258 136102
rect 40326 136046 40382 136102
rect 39954 135922 40010 135978
rect 40078 135922 40134 135978
rect 40202 135922 40258 135978
rect 40326 135922 40382 135978
rect 39954 118294 40010 118350
rect 40078 118294 40134 118350
rect 40202 118294 40258 118350
rect 40326 118294 40382 118350
rect 39954 118170 40010 118226
rect 40078 118170 40134 118226
rect 40202 118170 40258 118226
rect 40326 118170 40382 118226
rect 39954 118046 40010 118102
rect 40078 118046 40134 118102
rect 40202 118046 40258 118102
rect 40326 118046 40382 118102
rect 39954 117922 40010 117978
rect 40078 117922 40134 117978
rect 40202 117922 40258 117978
rect 40326 117922 40382 117978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 39954 64294 40010 64350
rect 40078 64294 40134 64350
rect 40202 64294 40258 64350
rect 40326 64294 40382 64350
rect 39954 64170 40010 64226
rect 40078 64170 40134 64226
rect 40202 64170 40258 64226
rect 40326 64170 40382 64226
rect 39954 64046 40010 64102
rect 40078 64046 40134 64102
rect 40202 64046 40258 64102
rect 40326 64046 40382 64102
rect 39954 63922 40010 63978
rect 40078 63922 40134 63978
rect 40202 63922 40258 63978
rect 40326 63922 40382 63978
rect 39954 46294 40010 46350
rect 40078 46294 40134 46350
rect 40202 46294 40258 46350
rect 40326 46294 40382 46350
rect 39954 46170 40010 46226
rect 40078 46170 40134 46226
rect 40202 46170 40258 46226
rect 40326 46170 40382 46226
rect 39954 46046 40010 46102
rect 40078 46046 40134 46102
rect 40202 46046 40258 46102
rect 40326 46046 40382 46102
rect 39954 45922 40010 45978
rect 40078 45922 40134 45978
rect 40202 45922 40258 45978
rect 40326 45922 40382 45978
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 41804 210842 41860 210898
rect 68012 237692 68068 237718
rect 68012 237662 68068 237692
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 71596 237482 71652 237538
rect 97674 382294 97730 382350
rect 97798 382294 97854 382350
rect 97922 382294 97978 382350
rect 98046 382294 98102 382350
rect 97674 382170 97730 382226
rect 97798 382170 97854 382226
rect 97922 382170 97978 382226
rect 98046 382170 98102 382226
rect 97674 382046 97730 382102
rect 97798 382046 97854 382102
rect 97922 382046 97978 382102
rect 98046 382046 98102 382102
rect 97674 381922 97730 381978
rect 97798 381922 97854 381978
rect 97922 381922 97978 381978
rect 98046 381922 98102 381978
rect 97674 364294 97730 364350
rect 97798 364294 97854 364350
rect 97922 364294 97978 364350
rect 98046 364294 98102 364350
rect 97674 364170 97730 364226
rect 97798 364170 97854 364226
rect 97922 364170 97978 364226
rect 98046 364170 98102 364226
rect 97674 364046 97730 364102
rect 97798 364046 97854 364102
rect 97922 364046 97978 364102
rect 98046 364046 98102 364102
rect 97674 363922 97730 363978
rect 97798 363922 97854 363978
rect 97922 363922 97978 363978
rect 98046 363922 98102 363978
rect 97674 346294 97730 346350
rect 97798 346294 97854 346350
rect 97922 346294 97978 346350
rect 98046 346294 98102 346350
rect 97674 346170 97730 346226
rect 97798 346170 97854 346226
rect 97922 346170 97978 346226
rect 98046 346170 98102 346226
rect 97674 346046 97730 346102
rect 97798 346046 97854 346102
rect 97922 346046 97978 346102
rect 98046 346046 98102 346102
rect 97674 345922 97730 345978
rect 97798 345922 97854 345978
rect 97922 345922 97978 345978
rect 98046 345922 98102 345978
rect 97674 328294 97730 328350
rect 97798 328294 97854 328350
rect 97922 328294 97978 328350
rect 98046 328294 98102 328350
rect 97674 328170 97730 328226
rect 97798 328170 97854 328226
rect 97922 328170 97978 328226
rect 98046 328170 98102 328226
rect 97674 328046 97730 328102
rect 97798 328046 97854 328102
rect 97922 328046 97978 328102
rect 98046 328046 98102 328102
rect 97674 327922 97730 327978
rect 97798 327922 97854 327978
rect 97922 327922 97978 327978
rect 98046 327922 98102 327978
rect 97674 310294 97730 310350
rect 97798 310294 97854 310350
rect 97922 310294 97978 310350
rect 98046 310294 98102 310350
rect 97674 310170 97730 310226
rect 97798 310170 97854 310226
rect 97922 310170 97978 310226
rect 98046 310170 98102 310226
rect 97674 310046 97730 310102
rect 97798 310046 97854 310102
rect 97922 310046 97978 310102
rect 98046 310046 98102 310102
rect 97674 309922 97730 309978
rect 97798 309922 97854 309978
rect 97922 309922 97978 309978
rect 98046 309922 98102 309978
rect 97674 292294 97730 292350
rect 97798 292294 97854 292350
rect 97922 292294 97978 292350
rect 98046 292294 98102 292350
rect 97674 292170 97730 292226
rect 97798 292170 97854 292226
rect 97922 292170 97978 292226
rect 98046 292170 98102 292226
rect 97674 292046 97730 292102
rect 97798 292046 97854 292102
rect 97922 292046 97978 292102
rect 98046 292046 98102 292102
rect 97674 291922 97730 291978
rect 97798 291922 97854 291978
rect 97922 291922 97978 291978
rect 98046 291922 98102 291978
rect 93996 275642 94052 275698
rect 97674 274294 97730 274350
rect 97798 274294 97854 274350
rect 97922 274294 97978 274350
rect 98046 274294 98102 274350
rect 97674 274170 97730 274226
rect 97798 274170 97854 274226
rect 97922 274170 97978 274226
rect 98046 274170 98102 274226
rect 97674 274046 97730 274102
rect 97798 274046 97854 274102
rect 97922 274046 97978 274102
rect 98046 274046 98102 274102
rect 97674 273922 97730 273978
rect 97798 273922 97854 273978
rect 97922 273922 97978 273978
rect 98046 273922 98102 273978
rect 93436 270602 93492 270658
rect 91756 237662 91812 237718
rect 97674 256294 97730 256350
rect 97798 256294 97854 256350
rect 97922 256294 97978 256350
rect 98046 256294 98102 256350
rect 97674 256170 97730 256226
rect 97798 256170 97854 256226
rect 97922 256170 97978 256226
rect 98046 256170 98102 256226
rect 97674 256046 97730 256102
rect 97798 256046 97854 256102
rect 97922 256046 97978 256102
rect 98046 256046 98102 256102
rect 97674 255922 97730 255978
rect 97798 255922 97854 255978
rect 97922 255922 97978 255978
rect 98046 255922 98102 255978
rect 97674 238294 97730 238350
rect 97798 238294 97854 238350
rect 97922 238294 97978 238350
rect 98046 238294 98102 238350
rect 97674 238170 97730 238226
rect 97798 238170 97854 238226
rect 97922 238170 97978 238226
rect 98046 238170 98102 238226
rect 97674 238046 97730 238102
rect 97798 238046 97854 238102
rect 97922 238046 97978 238102
rect 98046 238046 98102 238102
rect 97674 237922 97730 237978
rect 97798 237922 97854 237978
rect 97922 237922 97978 237978
rect 98046 237922 98102 237978
rect 91532 237482 91588 237538
rect 70674 226294 70730 226350
rect 70798 226294 70854 226350
rect 70922 226294 70978 226350
rect 71046 226294 71102 226350
rect 70674 226170 70730 226226
rect 70798 226170 70854 226226
rect 70922 226170 70978 226226
rect 71046 226170 71102 226226
rect 70674 226046 70730 226102
rect 70798 226046 70854 226102
rect 70922 226046 70978 226102
rect 71046 226046 71102 226102
rect 70674 225922 70730 225978
rect 70798 225922 70854 225978
rect 70922 225922 70978 225978
rect 71046 225922 71102 225978
rect 70674 208294 70730 208350
rect 70798 208294 70854 208350
rect 70922 208294 70978 208350
rect 71046 208294 71102 208350
rect 70674 208170 70730 208226
rect 70798 208170 70854 208226
rect 70922 208170 70978 208226
rect 71046 208170 71102 208226
rect 70674 208046 70730 208102
rect 70798 208046 70854 208102
rect 70922 208046 70978 208102
rect 71046 208046 71102 208102
rect 70674 207922 70730 207978
rect 70798 207922 70854 207978
rect 70922 207922 70978 207978
rect 71046 207922 71102 207978
rect 97674 220294 97730 220350
rect 97798 220294 97854 220350
rect 97922 220294 97978 220350
rect 98046 220294 98102 220350
rect 97674 220170 97730 220226
rect 97798 220170 97854 220226
rect 97922 220170 97978 220226
rect 98046 220170 98102 220226
rect 97674 220046 97730 220102
rect 97798 220046 97854 220102
rect 97922 220046 97978 220102
rect 98046 220046 98102 220102
rect 97674 219922 97730 219978
rect 97798 219922 97854 219978
rect 97922 219922 97978 219978
rect 98046 219922 98102 219978
rect 101394 460294 101450 460350
rect 101518 460294 101574 460350
rect 101642 460294 101698 460350
rect 101766 460294 101822 460350
rect 101394 460170 101450 460226
rect 101518 460170 101574 460226
rect 101642 460170 101698 460226
rect 101766 460170 101822 460226
rect 101394 460046 101450 460102
rect 101518 460046 101574 460102
rect 101642 460046 101698 460102
rect 101766 460046 101822 460102
rect 101394 459922 101450 459978
rect 101518 459922 101574 459978
rect 101642 459922 101698 459978
rect 101766 459922 101822 459978
rect 101394 442294 101450 442350
rect 101518 442294 101574 442350
rect 101642 442294 101698 442350
rect 101766 442294 101822 442350
rect 101394 442170 101450 442226
rect 101518 442170 101574 442226
rect 101642 442170 101698 442226
rect 101766 442170 101822 442226
rect 101394 442046 101450 442102
rect 101518 442046 101574 442102
rect 101642 442046 101698 442102
rect 101766 442046 101822 442102
rect 101394 441922 101450 441978
rect 101518 441922 101574 441978
rect 101642 441922 101698 441978
rect 101766 441922 101822 441978
rect 101394 424294 101450 424350
rect 101518 424294 101574 424350
rect 101642 424294 101698 424350
rect 101766 424294 101822 424350
rect 101394 424170 101450 424226
rect 101518 424170 101574 424226
rect 101642 424170 101698 424226
rect 101766 424170 101822 424226
rect 101394 424046 101450 424102
rect 101518 424046 101574 424102
rect 101642 424046 101698 424102
rect 101766 424046 101822 424102
rect 101394 423922 101450 423978
rect 101518 423922 101574 423978
rect 101642 423922 101698 423978
rect 101766 423922 101822 423978
rect 101394 406294 101450 406350
rect 101518 406294 101574 406350
rect 101642 406294 101698 406350
rect 101766 406294 101822 406350
rect 101394 406170 101450 406226
rect 101518 406170 101574 406226
rect 101642 406170 101698 406226
rect 101766 406170 101822 406226
rect 101394 406046 101450 406102
rect 101518 406046 101574 406102
rect 101642 406046 101698 406102
rect 101766 406046 101822 406102
rect 101394 405922 101450 405978
rect 101518 405922 101574 405978
rect 101642 405922 101698 405978
rect 101766 405922 101822 405978
rect 101394 388294 101450 388350
rect 101518 388294 101574 388350
rect 101642 388294 101698 388350
rect 101766 388294 101822 388350
rect 101394 388170 101450 388226
rect 101518 388170 101574 388226
rect 101642 388170 101698 388226
rect 101766 388170 101822 388226
rect 101394 388046 101450 388102
rect 101518 388046 101574 388102
rect 101642 388046 101698 388102
rect 101766 388046 101822 388102
rect 101394 387922 101450 387978
rect 101518 387922 101574 387978
rect 101642 387922 101698 387978
rect 101766 387922 101822 387978
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 128394 418294 128450 418350
rect 128518 418294 128574 418350
rect 128642 418294 128698 418350
rect 128766 418294 128822 418350
rect 128394 418170 128450 418226
rect 128518 418170 128574 418226
rect 128642 418170 128698 418226
rect 128766 418170 128822 418226
rect 128394 418046 128450 418102
rect 128518 418046 128574 418102
rect 128642 418046 128698 418102
rect 128766 418046 128822 418102
rect 128394 417922 128450 417978
rect 128518 417922 128574 417978
rect 128642 417922 128698 417978
rect 128766 417922 128822 417978
rect 128394 400294 128450 400350
rect 128518 400294 128574 400350
rect 128642 400294 128698 400350
rect 128766 400294 128822 400350
rect 128394 400170 128450 400226
rect 128518 400170 128574 400226
rect 128642 400170 128698 400226
rect 128766 400170 128822 400226
rect 128394 400046 128450 400102
rect 128518 400046 128574 400102
rect 128642 400046 128698 400102
rect 128766 400046 128822 400102
rect 128394 399922 128450 399978
rect 128518 399922 128574 399978
rect 128642 399922 128698 399978
rect 128766 399922 128822 399978
rect 128394 382294 128450 382350
rect 128518 382294 128574 382350
rect 128642 382294 128698 382350
rect 128766 382294 128822 382350
rect 128394 382170 128450 382226
rect 128518 382170 128574 382226
rect 128642 382170 128698 382226
rect 128766 382170 128822 382226
rect 128394 382046 128450 382102
rect 128518 382046 128574 382102
rect 128642 382046 128698 382102
rect 128766 382046 128822 382102
rect 128394 381922 128450 381978
rect 128518 381922 128574 381978
rect 128642 381922 128698 381978
rect 128766 381922 128822 381978
rect 101394 370294 101450 370350
rect 101518 370294 101574 370350
rect 101642 370294 101698 370350
rect 101766 370294 101822 370350
rect 101394 370170 101450 370226
rect 101518 370170 101574 370226
rect 101642 370170 101698 370226
rect 101766 370170 101822 370226
rect 101394 370046 101450 370102
rect 101518 370046 101574 370102
rect 101642 370046 101698 370102
rect 101766 370046 101822 370102
rect 101394 369922 101450 369978
rect 101518 369922 101574 369978
rect 101642 369922 101698 369978
rect 101766 369922 101822 369978
rect 101394 352294 101450 352350
rect 101518 352294 101574 352350
rect 101642 352294 101698 352350
rect 101766 352294 101822 352350
rect 101394 352170 101450 352226
rect 101518 352170 101574 352226
rect 101642 352170 101698 352226
rect 101766 352170 101822 352226
rect 101394 352046 101450 352102
rect 101518 352046 101574 352102
rect 101642 352046 101698 352102
rect 101766 352046 101822 352102
rect 101394 351922 101450 351978
rect 101518 351922 101574 351978
rect 101642 351922 101698 351978
rect 101766 351922 101822 351978
rect 101394 334294 101450 334350
rect 101518 334294 101574 334350
rect 101642 334294 101698 334350
rect 101766 334294 101822 334350
rect 101394 334170 101450 334226
rect 101518 334170 101574 334226
rect 101642 334170 101698 334226
rect 101766 334170 101822 334226
rect 101394 334046 101450 334102
rect 101518 334046 101574 334102
rect 101642 334046 101698 334102
rect 101766 334046 101822 334102
rect 101394 333922 101450 333978
rect 101518 333922 101574 333978
rect 101642 333922 101698 333978
rect 101766 333922 101822 333978
rect 101394 316294 101450 316350
rect 101518 316294 101574 316350
rect 101642 316294 101698 316350
rect 101766 316294 101822 316350
rect 101394 316170 101450 316226
rect 101518 316170 101574 316226
rect 101642 316170 101698 316226
rect 101766 316170 101822 316226
rect 101394 316046 101450 316102
rect 101518 316046 101574 316102
rect 101642 316046 101698 316102
rect 101766 316046 101822 316102
rect 101394 315922 101450 315978
rect 101518 315922 101574 315978
rect 101642 315922 101698 315978
rect 101766 315922 101822 315978
rect 101394 298294 101450 298350
rect 101518 298294 101574 298350
rect 101642 298294 101698 298350
rect 101766 298294 101822 298350
rect 101394 298170 101450 298226
rect 101518 298170 101574 298226
rect 101642 298170 101698 298226
rect 101766 298170 101822 298226
rect 101394 298046 101450 298102
rect 101518 298046 101574 298102
rect 101642 298046 101698 298102
rect 101766 298046 101822 298102
rect 101394 297922 101450 297978
rect 101518 297922 101574 297978
rect 101642 297922 101698 297978
rect 101766 297922 101822 297978
rect 108332 376442 108388 376498
rect 128394 364294 128450 364350
rect 128518 364294 128574 364350
rect 128642 364294 128698 364350
rect 128766 364294 128822 364350
rect 128394 364170 128450 364226
rect 128518 364170 128574 364226
rect 128642 364170 128698 364226
rect 128766 364170 128822 364226
rect 128394 364046 128450 364102
rect 128518 364046 128574 364102
rect 128642 364046 128698 364102
rect 128766 364046 128822 364102
rect 128394 363922 128450 363978
rect 128518 363922 128574 363978
rect 128642 363922 128698 363978
rect 128766 363922 128822 363978
rect 119518 346294 119574 346350
rect 119642 346294 119698 346350
rect 119518 346170 119574 346226
rect 119642 346170 119698 346226
rect 119518 346046 119574 346102
rect 119642 346046 119698 346102
rect 119518 345922 119574 345978
rect 119642 345922 119698 345978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 132114 424294 132170 424350
rect 132238 424294 132294 424350
rect 132362 424294 132418 424350
rect 132486 424294 132542 424350
rect 132114 424170 132170 424226
rect 132238 424170 132294 424226
rect 132362 424170 132418 424226
rect 132486 424170 132542 424226
rect 132114 424046 132170 424102
rect 132238 424046 132294 424102
rect 132362 424046 132418 424102
rect 132486 424046 132542 424102
rect 132114 423922 132170 423978
rect 132238 423922 132294 423978
rect 132362 423922 132418 423978
rect 132486 423922 132542 423978
rect 132114 406294 132170 406350
rect 132238 406294 132294 406350
rect 132362 406294 132418 406350
rect 132486 406294 132542 406350
rect 132114 406170 132170 406226
rect 132238 406170 132294 406226
rect 132362 406170 132418 406226
rect 132486 406170 132542 406226
rect 132114 406046 132170 406102
rect 132238 406046 132294 406102
rect 132362 406046 132418 406102
rect 132486 406046 132542 406102
rect 132114 405922 132170 405978
rect 132238 405922 132294 405978
rect 132362 405922 132418 405978
rect 132486 405922 132542 405978
rect 132114 388294 132170 388350
rect 132238 388294 132294 388350
rect 132362 388294 132418 388350
rect 132486 388294 132542 388350
rect 132114 388170 132170 388226
rect 132238 388170 132294 388226
rect 132362 388170 132418 388226
rect 132486 388170 132542 388226
rect 132114 388046 132170 388102
rect 132238 388046 132294 388102
rect 132362 388046 132418 388102
rect 132486 388046 132542 388102
rect 132114 387922 132170 387978
rect 132238 387922 132294 387978
rect 132362 387922 132418 387978
rect 132486 387922 132542 387978
rect 132114 370294 132170 370350
rect 132238 370294 132294 370350
rect 132362 370294 132418 370350
rect 132486 370294 132542 370350
rect 132114 370170 132170 370226
rect 132238 370170 132294 370226
rect 132362 370170 132418 370226
rect 132486 370170 132542 370226
rect 132114 370046 132170 370102
rect 132238 370046 132294 370102
rect 132362 370046 132418 370102
rect 132486 370046 132542 370102
rect 132114 369922 132170 369978
rect 132238 369922 132294 369978
rect 132362 369922 132418 369978
rect 132486 369922 132542 369978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 162834 550294 162890 550350
rect 162958 550294 163014 550350
rect 163082 550294 163138 550350
rect 163206 550294 163262 550350
rect 162834 550170 162890 550226
rect 162958 550170 163014 550226
rect 163082 550170 163138 550226
rect 163206 550170 163262 550226
rect 162834 550046 162890 550102
rect 162958 550046 163014 550102
rect 163082 550046 163138 550102
rect 163206 550046 163262 550102
rect 162834 549922 162890 549978
rect 162958 549922 163014 549978
rect 163082 549922 163138 549978
rect 163206 549922 163262 549978
rect 162834 532294 162890 532350
rect 162958 532294 163014 532350
rect 163082 532294 163138 532350
rect 163206 532294 163262 532350
rect 162834 532170 162890 532226
rect 162958 532170 163014 532226
rect 163082 532170 163138 532226
rect 163206 532170 163262 532226
rect 162834 532046 162890 532102
rect 162958 532046 163014 532102
rect 163082 532046 163138 532102
rect 163206 532046 163262 532102
rect 162834 531922 162890 531978
rect 162958 531922 163014 531978
rect 163082 531922 163138 531978
rect 163206 531922 163262 531978
rect 162834 514294 162890 514350
rect 162958 514294 163014 514350
rect 163082 514294 163138 514350
rect 163206 514294 163262 514350
rect 162834 514170 162890 514226
rect 162958 514170 163014 514226
rect 163082 514170 163138 514226
rect 163206 514170 163262 514226
rect 162834 514046 162890 514102
rect 162958 514046 163014 514102
rect 163082 514046 163138 514102
rect 163206 514046 163262 514102
rect 162834 513922 162890 513978
rect 162958 513922 163014 513978
rect 163082 513922 163138 513978
rect 163206 513922 163262 513978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 174636 573722 174692 573778
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 159114 418294 159170 418350
rect 159238 418294 159294 418350
rect 159362 418294 159418 418350
rect 159486 418294 159542 418350
rect 159114 418170 159170 418226
rect 159238 418170 159294 418226
rect 159362 418170 159418 418226
rect 159486 418170 159542 418226
rect 159114 418046 159170 418102
rect 159238 418046 159294 418102
rect 159362 418046 159418 418102
rect 159486 418046 159542 418102
rect 159114 417922 159170 417978
rect 159238 417922 159294 417978
rect 159362 417922 159418 417978
rect 159486 417922 159542 417978
rect 159114 400294 159170 400350
rect 159238 400294 159294 400350
rect 159362 400294 159418 400350
rect 159486 400294 159542 400350
rect 159114 400170 159170 400226
rect 159238 400170 159294 400226
rect 159362 400170 159418 400226
rect 159486 400170 159542 400226
rect 159114 400046 159170 400102
rect 159238 400046 159294 400102
rect 159362 400046 159418 400102
rect 159486 400046 159542 400102
rect 159114 399922 159170 399978
rect 159238 399922 159294 399978
rect 159362 399922 159418 399978
rect 159486 399922 159542 399978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 134878 352294 134934 352350
rect 135002 352294 135058 352350
rect 134878 352170 134934 352226
rect 135002 352170 135058 352226
rect 134878 352046 134934 352102
rect 135002 352046 135058 352102
rect 134878 351922 134934 351978
rect 135002 351922 135058 351978
rect 128394 346294 128450 346350
rect 128518 346294 128574 346350
rect 128642 346294 128698 346350
rect 128766 346294 128822 346350
rect 128394 346170 128450 346226
rect 128518 346170 128574 346226
rect 128642 346170 128698 346226
rect 128766 346170 128822 346226
rect 128394 346046 128450 346102
rect 128518 346046 128574 346102
rect 128642 346046 128698 346102
rect 128766 346046 128822 346102
rect 128394 345922 128450 345978
rect 128518 345922 128574 345978
rect 128642 345922 128698 345978
rect 128766 345922 128822 345978
rect 119518 328294 119574 328350
rect 119642 328294 119698 328350
rect 119518 328170 119574 328226
rect 119642 328170 119698 328226
rect 119518 328046 119574 328102
rect 119642 328046 119698 328102
rect 119518 327922 119574 327978
rect 119642 327922 119698 327978
rect 150238 346294 150294 346350
rect 150362 346294 150418 346350
rect 150238 346170 150294 346226
rect 150362 346170 150418 346226
rect 150238 346046 150294 346102
rect 150362 346046 150418 346102
rect 150238 345922 150294 345978
rect 150362 345922 150418 345978
rect 134878 334294 134934 334350
rect 135002 334294 135058 334350
rect 134878 334170 134934 334226
rect 135002 334170 135058 334226
rect 134878 334046 134934 334102
rect 135002 334046 135058 334102
rect 134878 333922 134934 333978
rect 135002 333922 135058 333978
rect 128394 328294 128450 328350
rect 128518 328294 128574 328350
rect 128642 328294 128698 328350
rect 128766 328294 128822 328350
rect 128394 328170 128450 328226
rect 128518 328170 128574 328226
rect 128642 328170 128698 328226
rect 128766 328170 128822 328226
rect 128394 328046 128450 328102
rect 128518 328046 128574 328102
rect 128642 328046 128698 328102
rect 128766 328046 128822 328102
rect 128394 327922 128450 327978
rect 128518 327922 128574 327978
rect 128642 327922 128698 327978
rect 128766 327922 128822 327978
rect 150238 328294 150294 328350
rect 150362 328294 150418 328350
rect 150238 328170 150294 328226
rect 150362 328170 150418 328226
rect 150238 328046 150294 328102
rect 150362 328046 150418 328102
rect 150238 327922 150294 327978
rect 150362 327922 150418 327978
rect 128394 310294 128450 310350
rect 128518 310294 128574 310350
rect 128642 310294 128698 310350
rect 128766 310294 128822 310350
rect 128394 310170 128450 310226
rect 128518 310170 128574 310226
rect 128642 310170 128698 310226
rect 128766 310170 128822 310226
rect 128394 310046 128450 310102
rect 128518 310046 128574 310102
rect 128642 310046 128698 310102
rect 128766 310046 128822 310102
rect 128394 309922 128450 309978
rect 128518 309922 128574 309978
rect 128642 309922 128698 309978
rect 128766 309922 128822 309978
rect 128394 292294 128450 292350
rect 128518 292294 128574 292350
rect 128642 292294 128698 292350
rect 128766 292294 128822 292350
rect 128394 292170 128450 292226
rect 128518 292170 128574 292226
rect 128642 292170 128698 292226
rect 128766 292170 128822 292226
rect 128394 292046 128450 292102
rect 128518 292046 128574 292102
rect 128642 292046 128698 292102
rect 128766 292046 128822 292102
rect 128394 291922 128450 291978
rect 128518 291922 128574 291978
rect 128642 291922 128698 291978
rect 128766 291922 128822 291978
rect 101394 280294 101450 280350
rect 101518 280294 101574 280350
rect 101642 280294 101698 280350
rect 101766 280294 101822 280350
rect 101394 280170 101450 280226
rect 101518 280170 101574 280226
rect 101642 280170 101698 280226
rect 101766 280170 101822 280226
rect 101394 280046 101450 280102
rect 101518 280046 101574 280102
rect 101642 280046 101698 280102
rect 101766 280046 101822 280102
rect 101394 279922 101450 279978
rect 101518 279922 101574 279978
rect 101642 279922 101698 279978
rect 101766 279922 101822 279978
rect 101394 262294 101450 262350
rect 101518 262294 101574 262350
rect 101642 262294 101698 262350
rect 101766 262294 101822 262350
rect 101394 262170 101450 262226
rect 101518 262170 101574 262226
rect 101642 262170 101698 262226
rect 101766 262170 101822 262226
rect 101394 262046 101450 262102
rect 101518 262046 101574 262102
rect 101642 262046 101698 262102
rect 101766 262046 101822 262102
rect 101394 261922 101450 261978
rect 101518 261922 101574 261978
rect 101642 261922 101698 261978
rect 101766 261922 101822 261978
rect 101394 244294 101450 244350
rect 101518 244294 101574 244350
rect 101642 244294 101698 244350
rect 101766 244294 101822 244350
rect 101394 244170 101450 244226
rect 101518 244170 101574 244226
rect 101642 244170 101698 244226
rect 101766 244170 101822 244226
rect 101394 244046 101450 244102
rect 101518 244046 101574 244102
rect 101642 244046 101698 244102
rect 101766 244046 101822 244102
rect 101394 243922 101450 243978
rect 101518 243922 101574 243978
rect 101642 243922 101698 243978
rect 101766 243922 101822 243978
rect 101394 226294 101450 226350
rect 101518 226294 101574 226350
rect 101642 226294 101698 226350
rect 101766 226294 101822 226350
rect 101394 226170 101450 226226
rect 101518 226170 101574 226226
rect 101642 226170 101698 226226
rect 101766 226170 101822 226226
rect 101394 226046 101450 226102
rect 101518 226046 101574 226102
rect 101642 226046 101698 226102
rect 101766 226046 101822 226102
rect 101394 225922 101450 225978
rect 101518 225922 101574 225978
rect 101642 225922 101698 225978
rect 101766 225922 101822 225978
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 101394 208294 101450 208350
rect 101518 208294 101574 208350
rect 101642 208294 101698 208350
rect 101766 208294 101822 208350
rect 101394 208170 101450 208226
rect 101518 208170 101574 208226
rect 101642 208170 101698 208226
rect 101766 208170 101822 208226
rect 101394 208046 101450 208102
rect 101518 208046 101574 208102
rect 101642 208046 101698 208102
rect 101766 208046 101822 208102
rect 101394 207922 101450 207978
rect 101518 207922 101574 207978
rect 101642 207922 101698 207978
rect 101766 207922 101822 207978
rect 132114 316294 132170 316350
rect 132238 316294 132294 316350
rect 132362 316294 132418 316350
rect 132486 316294 132542 316350
rect 132114 316170 132170 316226
rect 132238 316170 132294 316226
rect 132362 316170 132418 316226
rect 132486 316170 132542 316226
rect 132114 316046 132170 316102
rect 132238 316046 132294 316102
rect 132362 316046 132418 316102
rect 132486 316046 132542 316102
rect 132114 315922 132170 315978
rect 132238 315922 132294 315978
rect 132362 315922 132418 315978
rect 132486 315922 132542 315978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 132114 298294 132170 298350
rect 132238 298294 132294 298350
rect 132362 298294 132418 298350
rect 132486 298294 132542 298350
rect 132114 298170 132170 298226
rect 132238 298170 132294 298226
rect 132362 298170 132418 298226
rect 132486 298170 132542 298226
rect 132114 298046 132170 298102
rect 132238 298046 132294 298102
rect 132362 298046 132418 298102
rect 132486 298046 132542 298102
rect 132114 297922 132170 297978
rect 132238 297922 132294 297978
rect 132362 297922 132418 297978
rect 132486 297922 132542 297978
rect 137788 290582 137844 290638
rect 139244 290582 139300 290638
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 162834 424294 162890 424350
rect 162958 424294 163014 424350
rect 163082 424294 163138 424350
rect 163206 424294 163262 424350
rect 162834 424170 162890 424226
rect 162958 424170 163014 424226
rect 163082 424170 163138 424226
rect 163206 424170 163262 424226
rect 162834 424046 162890 424102
rect 162958 424046 163014 424102
rect 163082 424046 163138 424102
rect 163206 424046 163262 424102
rect 162834 423922 162890 423978
rect 162958 423922 163014 423978
rect 163082 423922 163138 423978
rect 163206 423922 163262 423978
rect 162834 406294 162890 406350
rect 162958 406294 163014 406350
rect 163082 406294 163138 406350
rect 163206 406294 163262 406350
rect 162834 406170 162890 406226
rect 162958 406170 163014 406226
rect 163082 406170 163138 406226
rect 163206 406170 163262 406226
rect 162834 406046 162890 406102
rect 162958 406046 163014 406102
rect 163082 406046 163138 406102
rect 163206 406046 163262 406102
rect 162834 405922 162890 405978
rect 162958 405922 163014 405978
rect 163082 405922 163138 405978
rect 163206 405922 163262 405978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 162834 352294 162890 352350
rect 162958 352294 163014 352350
rect 163082 352294 163138 352350
rect 163206 352294 163262 352350
rect 162834 352170 162890 352226
rect 162958 352170 163014 352226
rect 163082 352170 163138 352226
rect 163206 352170 163262 352226
rect 162834 352046 162890 352102
rect 162958 352046 163014 352102
rect 163082 352046 163138 352102
rect 163206 352046 163262 352102
rect 162834 351922 162890 351978
rect 162958 351922 163014 351978
rect 163082 351922 163138 351978
rect 163206 351922 163262 351978
rect 162834 334294 162890 334350
rect 162958 334294 163014 334350
rect 163082 334294 163138 334350
rect 163206 334294 163262 334350
rect 162834 334170 162890 334226
rect 162958 334170 163014 334226
rect 163082 334170 163138 334226
rect 163206 334170 163262 334226
rect 162834 334046 162890 334102
rect 162958 334046 163014 334102
rect 163082 334046 163138 334102
rect 163206 334046 163262 334102
rect 162834 333922 162890 333978
rect 162958 333922 163014 333978
rect 163082 333922 163138 333978
rect 163206 333922 163262 333978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 142078 280294 142134 280350
rect 142202 280294 142258 280350
rect 142078 280170 142134 280226
rect 142202 280170 142258 280226
rect 142078 280046 142134 280102
rect 142202 280046 142258 280102
rect 142078 279922 142134 279978
rect 142202 279922 142258 279978
rect 147902 280294 147958 280350
rect 148026 280294 148082 280350
rect 147902 280170 147958 280226
rect 148026 280170 148082 280226
rect 147902 280046 147958 280102
rect 148026 280046 148082 280102
rect 147902 279922 147958 279978
rect 148026 279922 148082 279978
rect 153726 280294 153782 280350
rect 153850 280294 153906 280350
rect 153726 280170 153782 280226
rect 153850 280170 153906 280226
rect 153726 280046 153782 280102
rect 153850 280046 153906 280102
rect 153726 279922 153782 279978
rect 153850 279922 153906 279978
rect 159550 280294 159606 280350
rect 159674 280294 159730 280350
rect 159550 280170 159606 280226
rect 159674 280170 159730 280226
rect 159550 280046 159606 280102
rect 159674 280046 159730 280102
rect 159550 279922 159606 279978
rect 159674 279922 159730 279978
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 138684 275642 138740 275698
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 138572 270602 138628 270658
rect 139166 274294 139222 274350
rect 139290 274294 139346 274350
rect 139166 274170 139222 274226
rect 139290 274170 139346 274226
rect 139166 274046 139222 274102
rect 139290 274046 139346 274102
rect 139166 273922 139222 273978
rect 139290 273922 139346 273978
rect 144990 274294 145046 274350
rect 145114 274294 145170 274350
rect 144990 274170 145046 274226
rect 145114 274170 145170 274226
rect 144990 274046 145046 274102
rect 145114 274046 145170 274102
rect 144990 273922 145046 273978
rect 145114 273922 145170 273978
rect 150814 274294 150870 274350
rect 150938 274294 150994 274350
rect 150814 274170 150870 274226
rect 150938 274170 150994 274226
rect 150814 274046 150870 274102
rect 150938 274046 150994 274102
rect 150814 273922 150870 273978
rect 150938 273922 150994 273978
rect 156638 274294 156694 274350
rect 156762 274294 156818 274350
rect 156638 274170 156694 274226
rect 156762 274170 156818 274226
rect 156638 274046 156694 274102
rect 156762 274046 156818 274102
rect 156638 273922 156694 273978
rect 156762 273922 156818 273978
rect 163436 280682 163492 280738
rect 164108 284642 164164 284698
rect 163884 278882 163940 278938
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 132114 208294 132170 208350
rect 132238 208294 132294 208350
rect 132362 208294 132418 208350
rect 132486 208294 132542 208350
rect 132114 208170 132170 208226
rect 132238 208170 132294 208226
rect 132362 208170 132418 208226
rect 132486 208170 132542 208226
rect 132114 208046 132170 208102
rect 132238 208046 132294 208102
rect 132362 208046 132418 208102
rect 132486 208046 132542 208102
rect 132114 207922 132170 207978
rect 132238 207922 132294 207978
rect 132362 207922 132418 207978
rect 132486 207922 132542 207978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 163996 277982 164052 278038
rect 165564 283022 165620 283078
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 167244 281402 167300 281458
rect 168924 286442 168980 286498
rect 169036 283202 169092 283258
rect 168476 277262 168532 277318
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 179676 571922 179732 571978
rect 176316 569582 176372 569638
rect 176988 234242 177044 234298
rect 177548 211742 177604 211798
rect 180012 569762 180068 569818
rect 179900 279602 179956 279658
rect 180460 288782 180516 288838
rect 184716 397322 184772 397378
rect 184518 364294 184574 364350
rect 184642 364294 184698 364350
rect 184518 364170 184574 364226
rect 184642 364170 184698 364226
rect 184518 364046 184574 364102
rect 184642 364046 184698 364102
rect 184518 363922 184574 363978
rect 184642 363922 184698 363978
rect 184518 346294 184574 346350
rect 184642 346294 184698 346350
rect 184518 346170 184574 346226
rect 184642 346170 184698 346226
rect 184518 346046 184574 346102
rect 184642 346046 184698 346102
rect 184518 345922 184574 345978
rect 184642 345922 184698 345978
rect 184518 328294 184574 328350
rect 184642 328294 184698 328350
rect 184518 328170 184574 328226
rect 184642 328170 184698 328226
rect 184518 328046 184574 328102
rect 184642 328046 184698 328102
rect 184518 327922 184574 327978
rect 184642 327922 184698 327978
rect 184518 310294 184574 310350
rect 184642 310294 184698 310350
rect 184518 310170 184574 310226
rect 184642 310170 184698 310226
rect 184518 310046 184574 310102
rect 184642 310046 184698 310102
rect 184518 309922 184574 309978
rect 184642 309922 184698 309978
rect 184518 292294 184574 292350
rect 184642 292294 184698 292350
rect 184518 292170 184574 292226
rect 184642 292170 184698 292226
rect 184518 292046 184574 292102
rect 184642 292046 184698 292102
rect 184518 291922 184574 291978
rect 184642 291922 184698 291978
rect 184828 290582 184884 290638
rect 183932 287162 183988 287218
rect 183932 279602 183988 279658
rect 180572 265382 180628 265438
rect 180684 261100 180740 261118
rect 180684 261062 180740 261100
rect 180684 260036 180740 260038
rect 180684 259982 180740 260036
rect 180684 258916 180740 258958
rect 180684 258902 180740 258916
rect 180572 257102 180628 257158
rect 180572 252242 180628 252298
rect 180684 252062 180740 252118
rect 184518 274294 184574 274350
rect 184642 274294 184698 274350
rect 184518 274170 184574 274226
rect 184642 274170 184698 274226
rect 184518 274046 184574 274102
rect 184642 274046 184698 274102
rect 184518 273922 184574 273978
rect 184642 273922 184698 273978
rect 184518 256294 184574 256350
rect 184642 256294 184698 256350
rect 184518 256170 184574 256226
rect 184642 256170 184698 256226
rect 184518 256046 184574 256102
rect 184642 256046 184698 256102
rect 184518 255922 184574 255978
rect 184642 255922 184698 255978
rect 185612 290582 185668 290638
rect 187292 287162 187348 287218
rect 187180 285722 187236 285778
rect 187292 283742 187348 283798
rect 187292 283022 187348 283078
rect 186396 282122 186452 282178
rect 187404 282122 187460 282178
rect 186396 280682 186452 280738
rect 186284 279602 186340 279658
rect 186284 278882 186340 278938
rect 187852 283742 187908 283798
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 188076 286442 188132 286498
rect 188076 285722 188132 285778
rect 188076 284642 188132 284698
rect 187964 283202 188020 283258
rect 187740 281402 187796 281458
rect 187628 279602 187684 279658
rect 187516 277982 187572 278038
rect 187404 261062 187460 261118
rect 187292 258902 187348 258958
rect 188076 277262 188132 277318
rect 187628 259982 187684 260038
rect 189196 404162 189252 404218
rect 189420 390482 189476 390538
rect 189084 277262 189140 277318
rect 189308 288962 189364 289018
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 189834 544294 189890 544350
rect 189958 544294 190014 544350
rect 190082 544294 190138 544350
rect 190206 544294 190262 544350
rect 189834 544170 189890 544226
rect 189958 544170 190014 544226
rect 190082 544170 190138 544226
rect 190206 544170 190262 544226
rect 189834 544046 189890 544102
rect 189958 544046 190014 544102
rect 190082 544046 190138 544102
rect 190206 544046 190262 544102
rect 189834 543922 189890 543978
rect 189958 543922 190014 543978
rect 190082 543922 190138 543978
rect 190206 543922 190262 543978
rect 189834 526294 189890 526350
rect 189958 526294 190014 526350
rect 190082 526294 190138 526350
rect 190206 526294 190262 526350
rect 189834 526170 189890 526226
rect 189958 526170 190014 526226
rect 190082 526170 190138 526226
rect 190206 526170 190262 526226
rect 189834 526046 189890 526102
rect 189958 526046 190014 526102
rect 190082 526046 190138 526102
rect 190206 526046 190262 526102
rect 189834 525922 189890 525978
rect 189958 525922 190014 525978
rect 190082 525922 190138 525978
rect 190206 525922 190262 525978
rect 189834 508294 189890 508350
rect 189958 508294 190014 508350
rect 190082 508294 190138 508350
rect 190206 508294 190262 508350
rect 189834 508170 189890 508226
rect 189958 508170 190014 508226
rect 190082 508170 190138 508226
rect 190206 508170 190262 508226
rect 189834 508046 189890 508102
rect 189958 508046 190014 508102
rect 190082 508046 190138 508102
rect 190206 508046 190262 508102
rect 189834 507922 189890 507978
rect 189958 507922 190014 507978
rect 190082 507922 190138 507978
rect 190206 507922 190262 507978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 189834 418294 189890 418350
rect 189958 418294 190014 418350
rect 190082 418294 190138 418350
rect 190206 418294 190262 418350
rect 189834 418170 189890 418226
rect 189958 418170 190014 418226
rect 190082 418170 190138 418226
rect 190206 418170 190262 418226
rect 189834 418046 189890 418102
rect 189958 418046 190014 418102
rect 190082 418046 190138 418102
rect 190206 418046 190262 418102
rect 189834 417922 189890 417978
rect 189958 417922 190014 417978
rect 190082 417922 190138 417978
rect 190206 417922 190262 417978
rect 189834 400294 189890 400350
rect 189958 400294 190014 400350
rect 190082 400294 190138 400350
rect 190206 400294 190262 400350
rect 189834 400170 189890 400226
rect 189958 400170 190014 400226
rect 190082 400170 190138 400226
rect 190206 400170 190262 400226
rect 189834 400046 189890 400102
rect 189958 400046 190014 400102
rect 190082 400046 190138 400102
rect 190206 400046 190262 400102
rect 189834 399922 189890 399978
rect 189958 399922 190014 399978
rect 190082 399922 190138 399978
rect 190206 399922 190262 399978
rect 191548 391562 191604 391618
rect 189834 382294 189890 382350
rect 189958 382294 190014 382350
rect 190082 382294 190138 382350
rect 190206 382294 190262 382350
rect 189834 382170 189890 382226
rect 189958 382170 190014 382226
rect 190082 382170 190138 382226
rect 190206 382170 190262 382226
rect 189834 382046 189890 382102
rect 189958 382046 190014 382102
rect 190082 382046 190138 382102
rect 190206 382046 190262 382102
rect 189834 381922 189890 381978
rect 189958 381922 190014 381978
rect 190082 381922 190138 381978
rect 190206 381922 190262 381978
rect 187628 231002 187684 231058
rect 189834 364294 189890 364350
rect 189958 364294 190014 364350
rect 190082 364294 190138 364350
rect 190206 364294 190262 364350
rect 189834 364170 189890 364226
rect 189958 364170 190014 364226
rect 190082 364170 190138 364226
rect 190206 364170 190262 364226
rect 189834 364046 189890 364102
rect 189958 364046 190014 364102
rect 190082 364046 190138 364102
rect 190206 364046 190262 364102
rect 189834 363922 189890 363978
rect 189958 363922 190014 363978
rect 190082 363922 190138 363978
rect 190206 363922 190262 363978
rect 189834 346294 189890 346350
rect 189958 346294 190014 346350
rect 190082 346294 190138 346350
rect 190206 346294 190262 346350
rect 189834 346170 189890 346226
rect 189958 346170 190014 346226
rect 190082 346170 190138 346226
rect 190206 346170 190262 346226
rect 189834 346046 189890 346102
rect 189958 346046 190014 346102
rect 190082 346046 190138 346102
rect 190206 346046 190262 346102
rect 189834 345922 189890 345978
rect 189958 345922 190014 345978
rect 190082 345922 190138 345978
rect 190206 345922 190262 345978
rect 189834 328294 189890 328350
rect 189958 328294 190014 328350
rect 190082 328294 190138 328350
rect 190206 328294 190262 328350
rect 189834 328170 189890 328226
rect 189958 328170 190014 328226
rect 190082 328170 190138 328226
rect 190206 328170 190262 328226
rect 189834 328046 189890 328102
rect 189958 328046 190014 328102
rect 190082 328046 190138 328102
rect 190206 328046 190262 328102
rect 189834 327922 189890 327978
rect 189958 327922 190014 327978
rect 190082 327922 190138 327978
rect 190206 327922 190262 327978
rect 189834 310294 189890 310350
rect 189958 310294 190014 310350
rect 190082 310294 190138 310350
rect 190206 310294 190262 310350
rect 189834 310170 189890 310226
rect 189958 310170 190014 310226
rect 190082 310170 190138 310226
rect 190206 310170 190262 310226
rect 189834 310046 189890 310102
rect 189958 310046 190014 310102
rect 190082 310046 190138 310102
rect 190206 310046 190262 310102
rect 189834 309922 189890 309978
rect 189958 309922 190014 309978
rect 190082 309922 190138 309978
rect 190206 309922 190262 309978
rect 189834 292294 189890 292350
rect 189958 292294 190014 292350
rect 190082 292294 190138 292350
rect 190206 292294 190262 292350
rect 189834 292170 189890 292226
rect 189958 292170 190014 292226
rect 190082 292170 190138 292226
rect 190206 292170 190262 292226
rect 189834 292046 189890 292102
rect 189958 292046 190014 292102
rect 190082 292046 190138 292102
rect 190206 292046 190262 292102
rect 189834 291922 189890 291978
rect 189958 291922 190014 291978
rect 190082 291922 190138 291978
rect 190206 291922 190262 291978
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 162834 208294 162890 208350
rect 162958 208294 163014 208350
rect 163082 208294 163138 208350
rect 163206 208294 163262 208350
rect 162834 208170 162890 208226
rect 162958 208170 163014 208226
rect 163082 208170 163138 208226
rect 163206 208170 163262 208226
rect 162834 208046 162890 208102
rect 162958 208046 163014 208102
rect 163082 208046 163138 208102
rect 163206 208046 163262 208102
rect 162834 207922 162890 207978
rect 162958 207922 163014 207978
rect 163082 207922 163138 207978
rect 163206 207922 163262 207978
rect 193554 568294 193610 568350
rect 193678 568294 193734 568350
rect 193802 568294 193858 568350
rect 193926 568294 193982 568350
rect 193554 568170 193610 568226
rect 193678 568170 193734 568226
rect 193802 568170 193858 568226
rect 193926 568170 193982 568226
rect 193554 568046 193610 568102
rect 193678 568046 193734 568102
rect 193802 568046 193858 568102
rect 193926 568046 193982 568102
rect 193554 567922 193610 567978
rect 193678 567922 193734 567978
rect 193802 567922 193858 567978
rect 193926 567922 193982 567978
rect 194518 562294 194574 562350
rect 194642 562294 194698 562350
rect 194518 562170 194574 562226
rect 194642 562170 194698 562226
rect 194518 562046 194574 562102
rect 194642 562046 194698 562102
rect 194518 561922 194574 561978
rect 194642 561922 194698 561978
rect 193554 550294 193610 550350
rect 193678 550294 193734 550350
rect 193802 550294 193858 550350
rect 193926 550294 193982 550350
rect 193554 550170 193610 550226
rect 193678 550170 193734 550226
rect 193802 550170 193858 550226
rect 193926 550170 193982 550226
rect 193554 550046 193610 550102
rect 193678 550046 193734 550102
rect 193802 550046 193858 550102
rect 193926 550046 193982 550102
rect 193554 549922 193610 549978
rect 193678 549922 193734 549978
rect 193802 549922 193858 549978
rect 193926 549922 193982 549978
rect 194518 544294 194574 544350
rect 194642 544294 194698 544350
rect 194518 544170 194574 544226
rect 194642 544170 194698 544226
rect 194518 544046 194574 544102
rect 194642 544046 194698 544102
rect 194518 543922 194574 543978
rect 194642 543922 194698 543978
rect 193554 532294 193610 532350
rect 193678 532294 193734 532350
rect 193802 532294 193858 532350
rect 193926 532294 193982 532350
rect 193554 532170 193610 532226
rect 193678 532170 193734 532226
rect 193802 532170 193858 532226
rect 193926 532170 193982 532226
rect 193554 532046 193610 532102
rect 193678 532046 193734 532102
rect 193802 532046 193858 532102
rect 193926 532046 193982 532102
rect 193554 531922 193610 531978
rect 193678 531922 193734 531978
rect 193802 531922 193858 531978
rect 193926 531922 193982 531978
rect 194518 526294 194574 526350
rect 194642 526294 194698 526350
rect 194518 526170 194574 526226
rect 194642 526170 194698 526226
rect 194518 526046 194574 526102
rect 194642 526046 194698 526102
rect 194518 525922 194574 525978
rect 194642 525922 194698 525978
rect 193554 514294 193610 514350
rect 193678 514294 193734 514350
rect 193802 514294 193858 514350
rect 193926 514294 193982 514350
rect 193554 514170 193610 514226
rect 193678 514170 193734 514226
rect 193802 514170 193858 514226
rect 193926 514170 193982 514226
rect 193554 514046 193610 514102
rect 193678 514046 193734 514102
rect 193802 514046 193858 514102
rect 193926 514046 193982 514102
rect 193554 513922 193610 513978
rect 193678 513922 193734 513978
rect 193802 513922 193858 513978
rect 193926 513922 193982 513978
rect 194518 508294 194574 508350
rect 194642 508294 194698 508350
rect 194518 508170 194574 508226
rect 194642 508170 194698 508226
rect 194518 508046 194574 508102
rect 194642 508046 194698 508102
rect 194518 507922 194574 507978
rect 194642 507922 194698 507978
rect 193554 496294 193610 496350
rect 193678 496294 193734 496350
rect 193802 496294 193858 496350
rect 193926 496294 193982 496350
rect 193554 496170 193610 496226
rect 193678 496170 193734 496226
rect 193802 496170 193858 496226
rect 193926 496170 193982 496226
rect 193554 496046 193610 496102
rect 193678 496046 193734 496102
rect 193802 496046 193858 496102
rect 193926 496046 193982 496102
rect 193554 495922 193610 495978
rect 193678 495922 193734 495978
rect 193802 495922 193858 495978
rect 193926 495922 193982 495978
rect 194518 490294 194574 490350
rect 194642 490294 194698 490350
rect 194518 490170 194574 490226
rect 194642 490170 194698 490226
rect 194518 490046 194574 490102
rect 194642 490046 194698 490102
rect 194518 489922 194574 489978
rect 194642 489922 194698 489978
rect 193554 478294 193610 478350
rect 193678 478294 193734 478350
rect 193802 478294 193858 478350
rect 193926 478294 193982 478350
rect 193554 478170 193610 478226
rect 193678 478170 193734 478226
rect 193802 478170 193858 478226
rect 193926 478170 193982 478226
rect 193554 478046 193610 478102
rect 193678 478046 193734 478102
rect 193802 478046 193858 478102
rect 193926 478046 193982 478102
rect 193554 477922 193610 477978
rect 193678 477922 193734 477978
rect 193802 477922 193858 477978
rect 193926 477922 193982 477978
rect 194518 472294 194574 472350
rect 194642 472294 194698 472350
rect 194518 472170 194574 472226
rect 194642 472170 194698 472226
rect 194518 472046 194574 472102
rect 194642 472046 194698 472102
rect 194518 471922 194574 471978
rect 194642 471922 194698 471978
rect 193554 460294 193610 460350
rect 193678 460294 193734 460350
rect 193802 460294 193858 460350
rect 193926 460294 193982 460350
rect 193554 460170 193610 460226
rect 193678 460170 193734 460226
rect 193802 460170 193858 460226
rect 193926 460170 193982 460226
rect 193554 460046 193610 460102
rect 193678 460046 193734 460102
rect 193802 460046 193858 460102
rect 193926 460046 193982 460102
rect 193554 459922 193610 459978
rect 193678 459922 193734 459978
rect 193802 459922 193858 459978
rect 193926 459922 193982 459978
rect 194518 454294 194574 454350
rect 194642 454294 194698 454350
rect 194518 454170 194574 454226
rect 194642 454170 194698 454226
rect 194518 454046 194574 454102
rect 194642 454046 194698 454102
rect 194518 453922 194574 453978
rect 194642 453922 194698 453978
rect 193554 442294 193610 442350
rect 193678 442294 193734 442350
rect 193802 442294 193858 442350
rect 193926 442294 193982 442350
rect 193554 442170 193610 442226
rect 193678 442170 193734 442226
rect 193802 442170 193858 442226
rect 193926 442170 193982 442226
rect 193554 442046 193610 442102
rect 193678 442046 193734 442102
rect 193802 442046 193858 442102
rect 193926 442046 193982 442102
rect 193554 441922 193610 441978
rect 193678 441922 193734 441978
rect 193802 441922 193858 441978
rect 193926 441922 193982 441978
rect 194518 436294 194574 436350
rect 194642 436294 194698 436350
rect 194518 436170 194574 436226
rect 194642 436170 194698 436226
rect 194518 436046 194574 436102
rect 194642 436046 194698 436102
rect 194518 435922 194574 435978
rect 194642 435922 194698 435978
rect 193554 424294 193610 424350
rect 193678 424294 193734 424350
rect 193802 424294 193858 424350
rect 193926 424294 193982 424350
rect 193554 424170 193610 424226
rect 193678 424170 193734 424226
rect 193802 424170 193858 424226
rect 193926 424170 193982 424226
rect 193554 424046 193610 424102
rect 193678 424046 193734 424102
rect 193802 424046 193858 424102
rect 193926 424046 193982 424102
rect 193554 423922 193610 423978
rect 193678 423922 193734 423978
rect 193802 423922 193858 423978
rect 193926 423922 193982 423978
rect 194518 418294 194574 418350
rect 194642 418294 194698 418350
rect 194518 418170 194574 418226
rect 194642 418170 194698 418226
rect 194518 418046 194574 418102
rect 194642 418046 194698 418102
rect 194518 417922 194574 417978
rect 194642 417922 194698 417978
rect 193554 406294 193610 406350
rect 193678 406294 193734 406350
rect 193802 406294 193858 406350
rect 193926 406294 193982 406350
rect 193554 406170 193610 406226
rect 193678 406170 193734 406226
rect 193802 406170 193858 406226
rect 193926 406170 193982 406226
rect 193554 406046 193610 406102
rect 193678 406046 193734 406102
rect 193802 406046 193858 406102
rect 193926 406046 193982 406102
rect 193554 405922 193610 405978
rect 193678 405922 193734 405978
rect 193802 405922 193858 405978
rect 193926 405922 193982 405978
rect 192892 391562 192948 391618
rect 197596 566162 197652 566218
rect 193554 388294 193610 388350
rect 193678 388294 193734 388350
rect 193802 388294 193858 388350
rect 193926 388294 193982 388350
rect 193554 388170 193610 388226
rect 193678 388170 193734 388226
rect 193802 388170 193858 388226
rect 193926 388170 193982 388226
rect 193554 388046 193610 388102
rect 193678 388046 193734 388102
rect 193802 388046 193858 388102
rect 193926 388046 193982 388102
rect 193554 387922 193610 387978
rect 193678 387922 193734 387978
rect 193802 387922 193858 387978
rect 193926 387922 193982 387978
rect 192668 219122 192724 219178
rect 192108 215882 192164 215938
rect 193554 370294 193610 370350
rect 193678 370294 193734 370350
rect 193802 370294 193858 370350
rect 193926 370294 193982 370350
rect 193554 370170 193610 370226
rect 193678 370170 193734 370226
rect 193802 370170 193858 370226
rect 193926 370170 193982 370226
rect 193554 370046 193610 370102
rect 193678 370046 193734 370102
rect 193802 370046 193858 370102
rect 193926 370046 193982 370102
rect 193554 369922 193610 369978
rect 193678 369922 193734 369978
rect 193802 369922 193858 369978
rect 193926 369922 193982 369978
rect 193554 352294 193610 352350
rect 193678 352294 193734 352350
rect 193802 352294 193858 352350
rect 193926 352294 193982 352350
rect 193554 352170 193610 352226
rect 193678 352170 193734 352226
rect 193802 352170 193858 352226
rect 193926 352170 193982 352226
rect 193554 352046 193610 352102
rect 193678 352046 193734 352102
rect 193802 352046 193858 352102
rect 193926 352046 193982 352102
rect 193554 351922 193610 351978
rect 193678 351922 193734 351978
rect 193802 351922 193858 351978
rect 193926 351922 193982 351978
rect 193554 334294 193610 334350
rect 193678 334294 193734 334350
rect 193802 334294 193858 334350
rect 193926 334294 193982 334350
rect 193554 334170 193610 334226
rect 193678 334170 193734 334226
rect 193802 334170 193858 334226
rect 193926 334170 193982 334226
rect 193554 334046 193610 334102
rect 193678 334046 193734 334102
rect 193802 334046 193858 334102
rect 193926 334046 193982 334102
rect 193554 333922 193610 333978
rect 193678 333922 193734 333978
rect 193802 333922 193858 333978
rect 193926 333922 193982 333978
rect 193554 316294 193610 316350
rect 193678 316294 193734 316350
rect 193802 316294 193858 316350
rect 193926 316294 193982 316350
rect 193554 316170 193610 316226
rect 193678 316170 193734 316226
rect 193802 316170 193858 316226
rect 193926 316170 193982 316226
rect 193554 316046 193610 316102
rect 193678 316046 193734 316102
rect 193802 316046 193858 316102
rect 193926 316046 193982 316102
rect 193554 315922 193610 315978
rect 193678 315922 193734 315978
rect 193802 315922 193858 315978
rect 193926 315922 193982 315978
rect 193554 298294 193610 298350
rect 193678 298294 193734 298350
rect 193802 298294 193858 298350
rect 193926 298294 193982 298350
rect 193554 298170 193610 298226
rect 193678 298170 193734 298226
rect 193802 298170 193858 298226
rect 193926 298170 193982 298226
rect 193554 298046 193610 298102
rect 193678 298046 193734 298102
rect 193802 298046 193858 298102
rect 193926 298046 193982 298102
rect 193554 297922 193610 297978
rect 193678 297922 193734 297978
rect 193802 297922 193858 297978
rect 193926 297922 193982 297978
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 191324 212462 191380 212518
rect 190764 211022 190820 211078
rect 195244 288962 195300 289018
rect 196028 288782 196084 288838
rect 195916 286442 195972 286498
rect 195692 285722 195748 285778
rect 195916 282302 195972 282358
rect 195804 257102 195860 257158
rect 195916 246842 195972 246898
rect 196252 239282 196308 239338
rect 193554 208294 193610 208350
rect 193678 208294 193734 208350
rect 193802 208294 193858 208350
rect 193926 208294 193982 208350
rect 193554 208170 193610 208226
rect 193678 208170 193734 208226
rect 193802 208170 193858 208226
rect 193926 208170 193982 208226
rect 193554 208046 193610 208102
rect 193678 208046 193734 208102
rect 193802 208046 193858 208102
rect 193926 208046 193982 208102
rect 193554 207922 193610 207978
rect 193678 207922 193734 207978
rect 193802 207922 193858 207978
rect 193926 207922 193982 207978
rect 197708 392282 197764 392338
rect 197820 386522 197876 386578
rect 199724 571202 199780 571258
rect 198156 380042 198212 380098
rect 198940 288782 198996 288838
rect 199164 379682 199220 379738
rect 199164 283742 199220 283798
rect 199388 282302 199444 282358
rect 199276 253682 199332 253738
rect 199276 252242 199332 252298
rect 199388 246842 199444 246898
rect 199612 389762 199668 389818
rect 199948 404162 200004 404218
rect 199878 370294 199934 370350
rect 200002 370294 200058 370350
rect 199878 370170 199934 370226
rect 200002 370170 200058 370226
rect 199878 370046 199934 370102
rect 200002 370046 200058 370102
rect 199878 369922 199934 369978
rect 200002 369922 200058 369978
rect 199878 352294 199934 352350
rect 200002 352294 200058 352350
rect 199878 352170 199934 352226
rect 200002 352170 200058 352226
rect 199878 352046 199934 352102
rect 200002 352046 200058 352102
rect 199878 351922 199934 351978
rect 200002 351922 200058 351978
rect 199878 334294 199934 334350
rect 200002 334294 200058 334350
rect 199878 334170 199934 334226
rect 200002 334170 200058 334226
rect 199878 334046 199934 334102
rect 200002 334046 200058 334102
rect 199878 333922 199934 333978
rect 200002 333922 200058 333978
rect 199878 316294 199934 316350
rect 200002 316294 200058 316350
rect 199878 316170 199934 316226
rect 200002 316170 200058 316226
rect 199878 316046 199934 316102
rect 200002 316046 200058 316102
rect 199878 315922 199934 315978
rect 200002 315922 200058 315978
rect 199878 298294 199934 298350
rect 200002 298294 200058 298350
rect 199878 298170 199934 298226
rect 200002 298170 200058 298226
rect 199878 298046 199934 298102
rect 200002 298046 200058 298102
rect 199878 297922 199934 297978
rect 200002 297922 200058 297978
rect 199878 280294 199934 280350
rect 200002 280294 200058 280350
rect 199878 280170 199934 280226
rect 200002 280170 200058 280226
rect 199878 280046 199934 280102
rect 200002 280046 200058 280102
rect 199878 279922 199934 279978
rect 200002 279922 200058 279978
rect 202412 570302 202468 570358
rect 201068 389942 201124 389998
rect 200732 265382 200788 265438
rect 200844 383102 200900 383158
rect 199878 262294 199934 262350
rect 200002 262294 200058 262350
rect 199878 262170 199934 262226
rect 200002 262170 200058 262226
rect 199878 262046 199934 262102
rect 200002 262046 200058 262102
rect 199878 261922 199934 261978
rect 200002 261922 200058 261978
rect 200732 253682 200788 253738
rect 199878 244294 199934 244350
rect 200002 244294 200058 244350
rect 199878 244170 199934 244226
rect 200002 244170 200058 244226
rect 199878 244046 199934 244102
rect 200002 244046 200058 244102
rect 199878 243922 199934 243978
rect 200002 243922 200058 243978
rect 201068 351062 201124 351118
rect 201068 307322 201124 307378
rect 201068 305882 201124 305938
rect 201180 300842 201236 300898
rect 201180 265562 201236 265618
rect 201292 224162 201348 224218
rect 200844 222542 200900 222598
rect 199612 217502 199668 217558
rect 202300 410642 202356 410698
rect 201628 351062 201684 351118
rect 201740 300842 201796 300898
rect 201740 265562 201796 265618
rect 201516 227582 201572 227638
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 203308 406682 203364 406738
rect 202524 387242 202580 387298
rect 202748 384902 202804 384958
rect 202524 376262 202580 376318
rect 202636 377882 202692 377938
rect 202636 372122 202692 372178
rect 202412 307322 202468 307378
rect 202524 283202 202580 283258
rect 202412 281402 202468 281458
rect 202636 252062 202692 252118
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 253708 570302 253764 570358
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 341068 571922 341124 571978
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 225238 562294 225294 562350
rect 225362 562294 225418 562350
rect 225238 562170 225294 562226
rect 225362 562170 225418 562226
rect 225238 562046 225294 562102
rect 225362 562046 225418 562102
rect 225238 561922 225294 561978
rect 225362 561922 225418 561978
rect 255958 562294 256014 562350
rect 256082 562294 256138 562350
rect 255958 562170 256014 562226
rect 256082 562170 256138 562226
rect 255958 562046 256014 562102
rect 256082 562046 256138 562102
rect 255958 561922 256014 561978
rect 256082 561922 256138 561978
rect 286678 562294 286734 562350
rect 286802 562294 286858 562350
rect 286678 562170 286734 562226
rect 286802 562170 286858 562226
rect 286678 562046 286734 562102
rect 286802 562046 286858 562102
rect 286678 561922 286734 561978
rect 286802 561922 286858 561978
rect 317398 562294 317454 562350
rect 317522 562294 317578 562350
rect 317398 562170 317454 562226
rect 317522 562170 317578 562226
rect 317398 562046 317454 562102
rect 317522 562046 317578 562102
rect 317398 561922 317454 561978
rect 317522 561922 317578 561978
rect 348118 562294 348174 562350
rect 348242 562294 348298 562350
rect 348118 562170 348174 562226
rect 348242 562170 348298 562226
rect 348118 562046 348174 562102
rect 348242 562046 348298 562102
rect 348118 561922 348174 561978
rect 348242 561922 348298 561978
rect 378838 562294 378894 562350
rect 378962 562294 379018 562350
rect 378838 562170 378894 562226
rect 378962 562170 379018 562226
rect 378838 562046 378894 562102
rect 378962 562046 379018 562102
rect 378838 561922 378894 561978
rect 378962 561922 379018 561978
rect 409558 562294 409614 562350
rect 409682 562294 409738 562350
rect 409558 562170 409614 562226
rect 409682 562170 409738 562226
rect 409558 562046 409614 562102
rect 409682 562046 409738 562102
rect 409558 561922 409614 561978
rect 409682 561922 409738 561978
rect 440278 562294 440334 562350
rect 440402 562294 440458 562350
rect 440278 562170 440334 562226
rect 440402 562170 440458 562226
rect 440278 562046 440334 562102
rect 440402 562046 440458 562102
rect 440278 561922 440334 561978
rect 440402 561922 440458 561978
rect 470998 562294 471054 562350
rect 471122 562294 471178 562350
rect 470998 562170 471054 562226
rect 471122 562170 471178 562226
rect 470998 562046 471054 562102
rect 471122 562046 471178 562102
rect 470998 561922 471054 561978
rect 471122 561922 471178 561978
rect 209878 550294 209934 550350
rect 210002 550294 210058 550350
rect 209878 550170 209934 550226
rect 210002 550170 210058 550226
rect 209878 550046 209934 550102
rect 210002 550046 210058 550102
rect 209878 549922 209934 549978
rect 210002 549922 210058 549978
rect 240598 550294 240654 550350
rect 240722 550294 240778 550350
rect 240598 550170 240654 550226
rect 240722 550170 240778 550226
rect 240598 550046 240654 550102
rect 240722 550046 240778 550102
rect 240598 549922 240654 549978
rect 240722 549922 240778 549978
rect 271318 550294 271374 550350
rect 271442 550294 271498 550350
rect 271318 550170 271374 550226
rect 271442 550170 271498 550226
rect 271318 550046 271374 550102
rect 271442 550046 271498 550102
rect 271318 549922 271374 549978
rect 271442 549922 271498 549978
rect 302038 550294 302094 550350
rect 302162 550294 302218 550350
rect 302038 550170 302094 550226
rect 302162 550170 302218 550226
rect 302038 550046 302094 550102
rect 302162 550046 302218 550102
rect 302038 549922 302094 549978
rect 302162 549922 302218 549978
rect 332758 550294 332814 550350
rect 332882 550294 332938 550350
rect 332758 550170 332814 550226
rect 332882 550170 332938 550226
rect 332758 550046 332814 550102
rect 332882 550046 332938 550102
rect 332758 549922 332814 549978
rect 332882 549922 332938 549978
rect 363478 550294 363534 550350
rect 363602 550294 363658 550350
rect 363478 550170 363534 550226
rect 363602 550170 363658 550226
rect 363478 550046 363534 550102
rect 363602 550046 363658 550102
rect 363478 549922 363534 549978
rect 363602 549922 363658 549978
rect 394198 550294 394254 550350
rect 394322 550294 394378 550350
rect 394198 550170 394254 550226
rect 394322 550170 394378 550226
rect 394198 550046 394254 550102
rect 394322 550046 394378 550102
rect 394198 549922 394254 549978
rect 394322 549922 394378 549978
rect 424918 550294 424974 550350
rect 425042 550294 425098 550350
rect 424918 550170 424974 550226
rect 425042 550170 425098 550226
rect 424918 550046 424974 550102
rect 425042 550046 425098 550102
rect 424918 549922 424974 549978
rect 425042 549922 425098 549978
rect 455638 550294 455694 550350
rect 455762 550294 455818 550350
rect 455638 550170 455694 550226
rect 455762 550170 455818 550226
rect 455638 550046 455694 550102
rect 455762 550046 455818 550102
rect 455638 549922 455694 549978
rect 455762 549922 455818 549978
rect 225238 544294 225294 544350
rect 225362 544294 225418 544350
rect 225238 544170 225294 544226
rect 225362 544170 225418 544226
rect 225238 544046 225294 544102
rect 225362 544046 225418 544102
rect 225238 543922 225294 543978
rect 225362 543922 225418 543978
rect 255958 544294 256014 544350
rect 256082 544294 256138 544350
rect 255958 544170 256014 544226
rect 256082 544170 256138 544226
rect 255958 544046 256014 544102
rect 256082 544046 256138 544102
rect 255958 543922 256014 543978
rect 256082 543922 256138 543978
rect 286678 544294 286734 544350
rect 286802 544294 286858 544350
rect 286678 544170 286734 544226
rect 286802 544170 286858 544226
rect 286678 544046 286734 544102
rect 286802 544046 286858 544102
rect 286678 543922 286734 543978
rect 286802 543922 286858 543978
rect 317398 544294 317454 544350
rect 317522 544294 317578 544350
rect 317398 544170 317454 544226
rect 317522 544170 317578 544226
rect 317398 544046 317454 544102
rect 317522 544046 317578 544102
rect 317398 543922 317454 543978
rect 317522 543922 317578 543978
rect 348118 544294 348174 544350
rect 348242 544294 348298 544350
rect 348118 544170 348174 544226
rect 348242 544170 348298 544226
rect 348118 544046 348174 544102
rect 348242 544046 348298 544102
rect 348118 543922 348174 543978
rect 348242 543922 348298 543978
rect 378838 544294 378894 544350
rect 378962 544294 379018 544350
rect 378838 544170 378894 544226
rect 378962 544170 379018 544226
rect 378838 544046 378894 544102
rect 378962 544046 379018 544102
rect 378838 543922 378894 543978
rect 378962 543922 379018 543978
rect 409558 544294 409614 544350
rect 409682 544294 409738 544350
rect 409558 544170 409614 544226
rect 409682 544170 409738 544226
rect 409558 544046 409614 544102
rect 409682 544046 409738 544102
rect 409558 543922 409614 543978
rect 409682 543922 409738 543978
rect 440278 544294 440334 544350
rect 440402 544294 440458 544350
rect 440278 544170 440334 544226
rect 440402 544170 440458 544226
rect 440278 544046 440334 544102
rect 440402 544046 440458 544102
rect 440278 543922 440334 543978
rect 440402 543922 440458 543978
rect 470998 544294 471054 544350
rect 471122 544294 471178 544350
rect 470998 544170 471054 544226
rect 471122 544170 471178 544226
rect 470998 544046 471054 544102
rect 471122 544046 471178 544102
rect 470998 543922 471054 543978
rect 471122 543922 471178 543978
rect 209878 532294 209934 532350
rect 210002 532294 210058 532350
rect 209878 532170 209934 532226
rect 210002 532170 210058 532226
rect 209878 532046 209934 532102
rect 210002 532046 210058 532102
rect 209878 531922 209934 531978
rect 210002 531922 210058 531978
rect 240598 532294 240654 532350
rect 240722 532294 240778 532350
rect 240598 532170 240654 532226
rect 240722 532170 240778 532226
rect 240598 532046 240654 532102
rect 240722 532046 240778 532102
rect 240598 531922 240654 531978
rect 240722 531922 240778 531978
rect 271318 532294 271374 532350
rect 271442 532294 271498 532350
rect 271318 532170 271374 532226
rect 271442 532170 271498 532226
rect 271318 532046 271374 532102
rect 271442 532046 271498 532102
rect 271318 531922 271374 531978
rect 271442 531922 271498 531978
rect 302038 532294 302094 532350
rect 302162 532294 302218 532350
rect 302038 532170 302094 532226
rect 302162 532170 302218 532226
rect 302038 532046 302094 532102
rect 302162 532046 302218 532102
rect 302038 531922 302094 531978
rect 302162 531922 302218 531978
rect 332758 532294 332814 532350
rect 332882 532294 332938 532350
rect 332758 532170 332814 532226
rect 332882 532170 332938 532226
rect 332758 532046 332814 532102
rect 332882 532046 332938 532102
rect 332758 531922 332814 531978
rect 332882 531922 332938 531978
rect 363478 532294 363534 532350
rect 363602 532294 363658 532350
rect 363478 532170 363534 532226
rect 363602 532170 363658 532226
rect 363478 532046 363534 532102
rect 363602 532046 363658 532102
rect 363478 531922 363534 531978
rect 363602 531922 363658 531978
rect 394198 532294 394254 532350
rect 394322 532294 394378 532350
rect 394198 532170 394254 532226
rect 394322 532170 394378 532226
rect 394198 532046 394254 532102
rect 394322 532046 394378 532102
rect 394198 531922 394254 531978
rect 394322 531922 394378 531978
rect 424918 532294 424974 532350
rect 425042 532294 425098 532350
rect 424918 532170 424974 532226
rect 425042 532170 425098 532226
rect 424918 532046 424974 532102
rect 425042 532046 425098 532102
rect 424918 531922 424974 531978
rect 425042 531922 425098 531978
rect 455638 532294 455694 532350
rect 455762 532294 455818 532350
rect 455638 532170 455694 532226
rect 455762 532170 455818 532226
rect 455638 532046 455694 532102
rect 455762 532046 455818 532102
rect 455638 531922 455694 531978
rect 455762 531922 455818 531978
rect 225238 526294 225294 526350
rect 225362 526294 225418 526350
rect 225238 526170 225294 526226
rect 225362 526170 225418 526226
rect 225238 526046 225294 526102
rect 225362 526046 225418 526102
rect 225238 525922 225294 525978
rect 225362 525922 225418 525978
rect 255958 526294 256014 526350
rect 256082 526294 256138 526350
rect 255958 526170 256014 526226
rect 256082 526170 256138 526226
rect 255958 526046 256014 526102
rect 256082 526046 256138 526102
rect 255958 525922 256014 525978
rect 256082 525922 256138 525978
rect 286678 526294 286734 526350
rect 286802 526294 286858 526350
rect 286678 526170 286734 526226
rect 286802 526170 286858 526226
rect 286678 526046 286734 526102
rect 286802 526046 286858 526102
rect 286678 525922 286734 525978
rect 286802 525922 286858 525978
rect 317398 526294 317454 526350
rect 317522 526294 317578 526350
rect 317398 526170 317454 526226
rect 317522 526170 317578 526226
rect 317398 526046 317454 526102
rect 317522 526046 317578 526102
rect 317398 525922 317454 525978
rect 317522 525922 317578 525978
rect 348118 526294 348174 526350
rect 348242 526294 348298 526350
rect 348118 526170 348174 526226
rect 348242 526170 348298 526226
rect 348118 526046 348174 526102
rect 348242 526046 348298 526102
rect 348118 525922 348174 525978
rect 348242 525922 348298 525978
rect 378838 526294 378894 526350
rect 378962 526294 379018 526350
rect 378838 526170 378894 526226
rect 378962 526170 379018 526226
rect 378838 526046 378894 526102
rect 378962 526046 379018 526102
rect 378838 525922 378894 525978
rect 378962 525922 379018 525978
rect 409558 526294 409614 526350
rect 409682 526294 409738 526350
rect 409558 526170 409614 526226
rect 409682 526170 409738 526226
rect 409558 526046 409614 526102
rect 409682 526046 409738 526102
rect 409558 525922 409614 525978
rect 409682 525922 409738 525978
rect 440278 526294 440334 526350
rect 440402 526294 440458 526350
rect 440278 526170 440334 526226
rect 440402 526170 440458 526226
rect 440278 526046 440334 526102
rect 440402 526046 440458 526102
rect 440278 525922 440334 525978
rect 440402 525922 440458 525978
rect 470998 526294 471054 526350
rect 471122 526294 471178 526350
rect 470998 526170 471054 526226
rect 471122 526170 471178 526226
rect 470998 526046 471054 526102
rect 471122 526046 471178 526102
rect 470998 525922 471054 525978
rect 471122 525922 471178 525978
rect 209878 514294 209934 514350
rect 210002 514294 210058 514350
rect 209878 514170 209934 514226
rect 210002 514170 210058 514226
rect 209878 514046 209934 514102
rect 210002 514046 210058 514102
rect 209878 513922 209934 513978
rect 210002 513922 210058 513978
rect 240598 514294 240654 514350
rect 240722 514294 240778 514350
rect 240598 514170 240654 514226
rect 240722 514170 240778 514226
rect 240598 514046 240654 514102
rect 240722 514046 240778 514102
rect 240598 513922 240654 513978
rect 240722 513922 240778 513978
rect 271318 514294 271374 514350
rect 271442 514294 271498 514350
rect 271318 514170 271374 514226
rect 271442 514170 271498 514226
rect 271318 514046 271374 514102
rect 271442 514046 271498 514102
rect 271318 513922 271374 513978
rect 271442 513922 271498 513978
rect 302038 514294 302094 514350
rect 302162 514294 302218 514350
rect 302038 514170 302094 514226
rect 302162 514170 302218 514226
rect 302038 514046 302094 514102
rect 302162 514046 302218 514102
rect 302038 513922 302094 513978
rect 302162 513922 302218 513978
rect 332758 514294 332814 514350
rect 332882 514294 332938 514350
rect 332758 514170 332814 514226
rect 332882 514170 332938 514226
rect 332758 514046 332814 514102
rect 332882 514046 332938 514102
rect 332758 513922 332814 513978
rect 332882 513922 332938 513978
rect 363478 514294 363534 514350
rect 363602 514294 363658 514350
rect 363478 514170 363534 514226
rect 363602 514170 363658 514226
rect 363478 514046 363534 514102
rect 363602 514046 363658 514102
rect 363478 513922 363534 513978
rect 363602 513922 363658 513978
rect 394198 514294 394254 514350
rect 394322 514294 394378 514350
rect 394198 514170 394254 514226
rect 394322 514170 394378 514226
rect 394198 514046 394254 514102
rect 394322 514046 394378 514102
rect 394198 513922 394254 513978
rect 394322 513922 394378 513978
rect 424918 514294 424974 514350
rect 425042 514294 425098 514350
rect 424918 514170 424974 514226
rect 425042 514170 425098 514226
rect 424918 514046 424974 514102
rect 425042 514046 425098 514102
rect 424918 513922 424974 513978
rect 425042 513922 425098 513978
rect 455638 514294 455694 514350
rect 455762 514294 455818 514350
rect 455638 514170 455694 514226
rect 455762 514170 455818 514226
rect 455638 514046 455694 514102
rect 455762 514046 455818 514102
rect 455638 513922 455694 513978
rect 455762 513922 455818 513978
rect 225238 508294 225294 508350
rect 225362 508294 225418 508350
rect 225238 508170 225294 508226
rect 225362 508170 225418 508226
rect 225238 508046 225294 508102
rect 225362 508046 225418 508102
rect 225238 507922 225294 507978
rect 225362 507922 225418 507978
rect 255958 508294 256014 508350
rect 256082 508294 256138 508350
rect 255958 508170 256014 508226
rect 256082 508170 256138 508226
rect 255958 508046 256014 508102
rect 256082 508046 256138 508102
rect 255958 507922 256014 507978
rect 256082 507922 256138 507978
rect 286678 508294 286734 508350
rect 286802 508294 286858 508350
rect 286678 508170 286734 508226
rect 286802 508170 286858 508226
rect 286678 508046 286734 508102
rect 286802 508046 286858 508102
rect 286678 507922 286734 507978
rect 286802 507922 286858 507978
rect 317398 508294 317454 508350
rect 317522 508294 317578 508350
rect 317398 508170 317454 508226
rect 317522 508170 317578 508226
rect 317398 508046 317454 508102
rect 317522 508046 317578 508102
rect 317398 507922 317454 507978
rect 317522 507922 317578 507978
rect 348118 508294 348174 508350
rect 348242 508294 348298 508350
rect 348118 508170 348174 508226
rect 348242 508170 348298 508226
rect 348118 508046 348174 508102
rect 348242 508046 348298 508102
rect 348118 507922 348174 507978
rect 348242 507922 348298 507978
rect 378838 508294 378894 508350
rect 378962 508294 379018 508350
rect 378838 508170 378894 508226
rect 378962 508170 379018 508226
rect 378838 508046 378894 508102
rect 378962 508046 379018 508102
rect 378838 507922 378894 507978
rect 378962 507922 379018 507978
rect 409558 508294 409614 508350
rect 409682 508294 409738 508350
rect 409558 508170 409614 508226
rect 409682 508170 409738 508226
rect 409558 508046 409614 508102
rect 409682 508046 409738 508102
rect 409558 507922 409614 507978
rect 409682 507922 409738 507978
rect 440278 508294 440334 508350
rect 440402 508294 440458 508350
rect 440278 508170 440334 508226
rect 440402 508170 440458 508226
rect 440278 508046 440334 508102
rect 440402 508046 440458 508102
rect 440278 507922 440334 507978
rect 440402 507922 440458 507978
rect 470998 508294 471054 508350
rect 471122 508294 471178 508350
rect 470998 508170 471054 508226
rect 471122 508170 471178 508226
rect 470998 508046 471054 508102
rect 471122 508046 471178 508102
rect 470998 507922 471054 507978
rect 471122 507922 471178 507978
rect 209878 496294 209934 496350
rect 210002 496294 210058 496350
rect 209878 496170 209934 496226
rect 210002 496170 210058 496226
rect 209878 496046 209934 496102
rect 210002 496046 210058 496102
rect 209878 495922 209934 495978
rect 210002 495922 210058 495978
rect 240598 496294 240654 496350
rect 240722 496294 240778 496350
rect 240598 496170 240654 496226
rect 240722 496170 240778 496226
rect 240598 496046 240654 496102
rect 240722 496046 240778 496102
rect 240598 495922 240654 495978
rect 240722 495922 240778 495978
rect 271318 496294 271374 496350
rect 271442 496294 271498 496350
rect 271318 496170 271374 496226
rect 271442 496170 271498 496226
rect 271318 496046 271374 496102
rect 271442 496046 271498 496102
rect 271318 495922 271374 495978
rect 271442 495922 271498 495978
rect 302038 496294 302094 496350
rect 302162 496294 302218 496350
rect 302038 496170 302094 496226
rect 302162 496170 302218 496226
rect 302038 496046 302094 496102
rect 302162 496046 302218 496102
rect 302038 495922 302094 495978
rect 302162 495922 302218 495978
rect 332758 496294 332814 496350
rect 332882 496294 332938 496350
rect 332758 496170 332814 496226
rect 332882 496170 332938 496226
rect 332758 496046 332814 496102
rect 332882 496046 332938 496102
rect 332758 495922 332814 495978
rect 332882 495922 332938 495978
rect 363478 496294 363534 496350
rect 363602 496294 363658 496350
rect 363478 496170 363534 496226
rect 363602 496170 363658 496226
rect 363478 496046 363534 496102
rect 363602 496046 363658 496102
rect 363478 495922 363534 495978
rect 363602 495922 363658 495978
rect 394198 496294 394254 496350
rect 394322 496294 394378 496350
rect 394198 496170 394254 496226
rect 394322 496170 394378 496226
rect 394198 496046 394254 496102
rect 394322 496046 394378 496102
rect 394198 495922 394254 495978
rect 394322 495922 394378 495978
rect 424918 496294 424974 496350
rect 425042 496294 425098 496350
rect 424918 496170 424974 496226
rect 425042 496170 425098 496226
rect 424918 496046 424974 496102
rect 425042 496046 425098 496102
rect 424918 495922 424974 495978
rect 425042 495922 425098 495978
rect 455638 496294 455694 496350
rect 455762 496294 455818 496350
rect 455638 496170 455694 496226
rect 455762 496170 455818 496226
rect 455638 496046 455694 496102
rect 455762 496046 455818 496102
rect 455638 495922 455694 495978
rect 455762 495922 455818 495978
rect 225238 490294 225294 490350
rect 225362 490294 225418 490350
rect 225238 490170 225294 490226
rect 225362 490170 225418 490226
rect 225238 490046 225294 490102
rect 225362 490046 225418 490102
rect 225238 489922 225294 489978
rect 225362 489922 225418 489978
rect 255958 490294 256014 490350
rect 256082 490294 256138 490350
rect 255958 490170 256014 490226
rect 256082 490170 256138 490226
rect 255958 490046 256014 490102
rect 256082 490046 256138 490102
rect 255958 489922 256014 489978
rect 256082 489922 256138 489978
rect 286678 490294 286734 490350
rect 286802 490294 286858 490350
rect 286678 490170 286734 490226
rect 286802 490170 286858 490226
rect 286678 490046 286734 490102
rect 286802 490046 286858 490102
rect 286678 489922 286734 489978
rect 286802 489922 286858 489978
rect 317398 490294 317454 490350
rect 317522 490294 317578 490350
rect 317398 490170 317454 490226
rect 317522 490170 317578 490226
rect 317398 490046 317454 490102
rect 317522 490046 317578 490102
rect 317398 489922 317454 489978
rect 317522 489922 317578 489978
rect 348118 490294 348174 490350
rect 348242 490294 348298 490350
rect 348118 490170 348174 490226
rect 348242 490170 348298 490226
rect 348118 490046 348174 490102
rect 348242 490046 348298 490102
rect 348118 489922 348174 489978
rect 348242 489922 348298 489978
rect 378838 490294 378894 490350
rect 378962 490294 379018 490350
rect 378838 490170 378894 490226
rect 378962 490170 379018 490226
rect 378838 490046 378894 490102
rect 378962 490046 379018 490102
rect 378838 489922 378894 489978
rect 378962 489922 379018 489978
rect 409558 490294 409614 490350
rect 409682 490294 409738 490350
rect 409558 490170 409614 490226
rect 409682 490170 409738 490226
rect 409558 490046 409614 490102
rect 409682 490046 409738 490102
rect 409558 489922 409614 489978
rect 409682 489922 409738 489978
rect 440278 490294 440334 490350
rect 440402 490294 440458 490350
rect 440278 490170 440334 490226
rect 440402 490170 440458 490226
rect 440278 490046 440334 490102
rect 440402 490046 440458 490102
rect 440278 489922 440334 489978
rect 440402 489922 440458 489978
rect 470998 490294 471054 490350
rect 471122 490294 471178 490350
rect 470998 490170 471054 490226
rect 471122 490170 471178 490226
rect 470998 490046 471054 490102
rect 471122 490046 471178 490102
rect 470998 489922 471054 489978
rect 471122 489922 471178 489978
rect 209878 478294 209934 478350
rect 210002 478294 210058 478350
rect 209878 478170 209934 478226
rect 210002 478170 210058 478226
rect 209878 478046 209934 478102
rect 210002 478046 210058 478102
rect 209878 477922 209934 477978
rect 210002 477922 210058 477978
rect 240598 478294 240654 478350
rect 240722 478294 240778 478350
rect 240598 478170 240654 478226
rect 240722 478170 240778 478226
rect 240598 478046 240654 478102
rect 240722 478046 240778 478102
rect 240598 477922 240654 477978
rect 240722 477922 240778 477978
rect 271318 478294 271374 478350
rect 271442 478294 271498 478350
rect 271318 478170 271374 478226
rect 271442 478170 271498 478226
rect 271318 478046 271374 478102
rect 271442 478046 271498 478102
rect 271318 477922 271374 477978
rect 271442 477922 271498 477978
rect 302038 478294 302094 478350
rect 302162 478294 302218 478350
rect 302038 478170 302094 478226
rect 302162 478170 302218 478226
rect 302038 478046 302094 478102
rect 302162 478046 302218 478102
rect 302038 477922 302094 477978
rect 302162 477922 302218 477978
rect 332758 478294 332814 478350
rect 332882 478294 332938 478350
rect 332758 478170 332814 478226
rect 332882 478170 332938 478226
rect 332758 478046 332814 478102
rect 332882 478046 332938 478102
rect 332758 477922 332814 477978
rect 332882 477922 332938 477978
rect 363478 478294 363534 478350
rect 363602 478294 363658 478350
rect 363478 478170 363534 478226
rect 363602 478170 363658 478226
rect 363478 478046 363534 478102
rect 363602 478046 363658 478102
rect 363478 477922 363534 477978
rect 363602 477922 363658 477978
rect 394198 478294 394254 478350
rect 394322 478294 394378 478350
rect 394198 478170 394254 478226
rect 394322 478170 394378 478226
rect 394198 478046 394254 478102
rect 394322 478046 394378 478102
rect 394198 477922 394254 477978
rect 394322 477922 394378 477978
rect 424918 478294 424974 478350
rect 425042 478294 425098 478350
rect 424918 478170 424974 478226
rect 425042 478170 425098 478226
rect 424918 478046 424974 478102
rect 425042 478046 425098 478102
rect 424918 477922 424974 477978
rect 425042 477922 425098 477978
rect 455638 478294 455694 478350
rect 455762 478294 455818 478350
rect 455638 478170 455694 478226
rect 455762 478170 455818 478226
rect 455638 478046 455694 478102
rect 455762 478046 455818 478102
rect 455638 477922 455694 477978
rect 455762 477922 455818 477978
rect 225238 472294 225294 472350
rect 225362 472294 225418 472350
rect 225238 472170 225294 472226
rect 225362 472170 225418 472226
rect 225238 472046 225294 472102
rect 225362 472046 225418 472102
rect 225238 471922 225294 471978
rect 225362 471922 225418 471978
rect 255958 472294 256014 472350
rect 256082 472294 256138 472350
rect 255958 472170 256014 472226
rect 256082 472170 256138 472226
rect 255958 472046 256014 472102
rect 256082 472046 256138 472102
rect 255958 471922 256014 471978
rect 256082 471922 256138 471978
rect 286678 472294 286734 472350
rect 286802 472294 286858 472350
rect 286678 472170 286734 472226
rect 286802 472170 286858 472226
rect 286678 472046 286734 472102
rect 286802 472046 286858 472102
rect 286678 471922 286734 471978
rect 286802 471922 286858 471978
rect 317398 472294 317454 472350
rect 317522 472294 317578 472350
rect 317398 472170 317454 472226
rect 317522 472170 317578 472226
rect 317398 472046 317454 472102
rect 317522 472046 317578 472102
rect 317398 471922 317454 471978
rect 317522 471922 317578 471978
rect 348118 472294 348174 472350
rect 348242 472294 348298 472350
rect 348118 472170 348174 472226
rect 348242 472170 348298 472226
rect 348118 472046 348174 472102
rect 348242 472046 348298 472102
rect 348118 471922 348174 471978
rect 348242 471922 348298 471978
rect 378838 472294 378894 472350
rect 378962 472294 379018 472350
rect 378838 472170 378894 472226
rect 378962 472170 379018 472226
rect 378838 472046 378894 472102
rect 378962 472046 379018 472102
rect 378838 471922 378894 471978
rect 378962 471922 379018 471978
rect 409558 472294 409614 472350
rect 409682 472294 409738 472350
rect 409558 472170 409614 472226
rect 409682 472170 409738 472226
rect 409558 472046 409614 472102
rect 409682 472046 409738 472102
rect 409558 471922 409614 471978
rect 409682 471922 409738 471978
rect 440278 472294 440334 472350
rect 440402 472294 440458 472350
rect 440278 472170 440334 472226
rect 440402 472170 440458 472226
rect 440278 472046 440334 472102
rect 440402 472046 440458 472102
rect 440278 471922 440334 471978
rect 440402 471922 440458 471978
rect 470998 472294 471054 472350
rect 471122 472294 471178 472350
rect 470998 472170 471054 472226
rect 471122 472170 471178 472226
rect 470998 472046 471054 472102
rect 471122 472046 471178 472102
rect 470998 471922 471054 471978
rect 471122 471922 471178 471978
rect 209878 460294 209934 460350
rect 210002 460294 210058 460350
rect 209878 460170 209934 460226
rect 210002 460170 210058 460226
rect 209878 460046 209934 460102
rect 210002 460046 210058 460102
rect 209878 459922 209934 459978
rect 210002 459922 210058 459978
rect 240598 460294 240654 460350
rect 240722 460294 240778 460350
rect 240598 460170 240654 460226
rect 240722 460170 240778 460226
rect 240598 460046 240654 460102
rect 240722 460046 240778 460102
rect 240598 459922 240654 459978
rect 240722 459922 240778 459978
rect 271318 460294 271374 460350
rect 271442 460294 271498 460350
rect 271318 460170 271374 460226
rect 271442 460170 271498 460226
rect 271318 460046 271374 460102
rect 271442 460046 271498 460102
rect 271318 459922 271374 459978
rect 271442 459922 271498 459978
rect 302038 460294 302094 460350
rect 302162 460294 302218 460350
rect 302038 460170 302094 460226
rect 302162 460170 302218 460226
rect 302038 460046 302094 460102
rect 302162 460046 302218 460102
rect 302038 459922 302094 459978
rect 302162 459922 302218 459978
rect 332758 460294 332814 460350
rect 332882 460294 332938 460350
rect 332758 460170 332814 460226
rect 332882 460170 332938 460226
rect 332758 460046 332814 460102
rect 332882 460046 332938 460102
rect 332758 459922 332814 459978
rect 332882 459922 332938 459978
rect 363478 460294 363534 460350
rect 363602 460294 363658 460350
rect 363478 460170 363534 460226
rect 363602 460170 363658 460226
rect 363478 460046 363534 460102
rect 363602 460046 363658 460102
rect 363478 459922 363534 459978
rect 363602 459922 363658 459978
rect 394198 460294 394254 460350
rect 394322 460294 394378 460350
rect 394198 460170 394254 460226
rect 394322 460170 394378 460226
rect 394198 460046 394254 460102
rect 394322 460046 394378 460102
rect 394198 459922 394254 459978
rect 394322 459922 394378 459978
rect 424918 460294 424974 460350
rect 425042 460294 425098 460350
rect 424918 460170 424974 460226
rect 425042 460170 425098 460226
rect 424918 460046 424974 460102
rect 425042 460046 425098 460102
rect 424918 459922 424974 459978
rect 425042 459922 425098 459978
rect 455638 460294 455694 460350
rect 455762 460294 455818 460350
rect 455638 460170 455694 460226
rect 455762 460170 455818 460226
rect 455638 460046 455694 460102
rect 455762 460046 455818 460102
rect 455638 459922 455694 459978
rect 455762 459922 455818 459978
rect 225238 454294 225294 454350
rect 225362 454294 225418 454350
rect 225238 454170 225294 454226
rect 225362 454170 225418 454226
rect 225238 454046 225294 454102
rect 225362 454046 225418 454102
rect 225238 453922 225294 453978
rect 225362 453922 225418 453978
rect 255958 454294 256014 454350
rect 256082 454294 256138 454350
rect 255958 454170 256014 454226
rect 256082 454170 256138 454226
rect 255958 454046 256014 454102
rect 256082 454046 256138 454102
rect 255958 453922 256014 453978
rect 256082 453922 256138 453978
rect 286678 454294 286734 454350
rect 286802 454294 286858 454350
rect 286678 454170 286734 454226
rect 286802 454170 286858 454226
rect 286678 454046 286734 454102
rect 286802 454046 286858 454102
rect 286678 453922 286734 453978
rect 286802 453922 286858 453978
rect 317398 454294 317454 454350
rect 317522 454294 317578 454350
rect 317398 454170 317454 454226
rect 317522 454170 317578 454226
rect 317398 454046 317454 454102
rect 317522 454046 317578 454102
rect 317398 453922 317454 453978
rect 317522 453922 317578 453978
rect 348118 454294 348174 454350
rect 348242 454294 348298 454350
rect 348118 454170 348174 454226
rect 348242 454170 348298 454226
rect 348118 454046 348174 454102
rect 348242 454046 348298 454102
rect 348118 453922 348174 453978
rect 348242 453922 348298 453978
rect 378838 454294 378894 454350
rect 378962 454294 379018 454350
rect 378838 454170 378894 454226
rect 378962 454170 379018 454226
rect 378838 454046 378894 454102
rect 378962 454046 379018 454102
rect 378838 453922 378894 453978
rect 378962 453922 379018 453978
rect 409558 454294 409614 454350
rect 409682 454294 409738 454350
rect 409558 454170 409614 454226
rect 409682 454170 409738 454226
rect 409558 454046 409614 454102
rect 409682 454046 409738 454102
rect 409558 453922 409614 453978
rect 409682 453922 409738 453978
rect 440278 454294 440334 454350
rect 440402 454294 440458 454350
rect 440278 454170 440334 454226
rect 440402 454170 440458 454226
rect 440278 454046 440334 454102
rect 440402 454046 440458 454102
rect 440278 453922 440334 453978
rect 440402 453922 440458 453978
rect 470998 454294 471054 454350
rect 471122 454294 471178 454350
rect 470998 454170 471054 454226
rect 471122 454170 471178 454226
rect 470998 454046 471054 454102
rect 471122 454046 471178 454102
rect 470998 453922 471054 453978
rect 471122 453922 471178 453978
rect 209878 442294 209934 442350
rect 210002 442294 210058 442350
rect 209878 442170 209934 442226
rect 210002 442170 210058 442226
rect 209878 442046 209934 442102
rect 210002 442046 210058 442102
rect 209878 441922 209934 441978
rect 210002 441922 210058 441978
rect 240598 442294 240654 442350
rect 240722 442294 240778 442350
rect 240598 442170 240654 442226
rect 240722 442170 240778 442226
rect 240598 442046 240654 442102
rect 240722 442046 240778 442102
rect 240598 441922 240654 441978
rect 240722 441922 240778 441978
rect 271318 442294 271374 442350
rect 271442 442294 271498 442350
rect 271318 442170 271374 442226
rect 271442 442170 271498 442226
rect 271318 442046 271374 442102
rect 271442 442046 271498 442102
rect 271318 441922 271374 441978
rect 271442 441922 271498 441978
rect 302038 442294 302094 442350
rect 302162 442294 302218 442350
rect 302038 442170 302094 442226
rect 302162 442170 302218 442226
rect 302038 442046 302094 442102
rect 302162 442046 302218 442102
rect 302038 441922 302094 441978
rect 302162 441922 302218 441978
rect 332758 442294 332814 442350
rect 332882 442294 332938 442350
rect 332758 442170 332814 442226
rect 332882 442170 332938 442226
rect 332758 442046 332814 442102
rect 332882 442046 332938 442102
rect 332758 441922 332814 441978
rect 332882 441922 332938 441978
rect 363478 442294 363534 442350
rect 363602 442294 363658 442350
rect 363478 442170 363534 442226
rect 363602 442170 363658 442226
rect 363478 442046 363534 442102
rect 363602 442046 363658 442102
rect 363478 441922 363534 441978
rect 363602 441922 363658 441978
rect 394198 442294 394254 442350
rect 394322 442294 394378 442350
rect 394198 442170 394254 442226
rect 394322 442170 394378 442226
rect 394198 442046 394254 442102
rect 394322 442046 394378 442102
rect 394198 441922 394254 441978
rect 394322 441922 394378 441978
rect 424918 442294 424974 442350
rect 425042 442294 425098 442350
rect 424918 442170 424974 442226
rect 425042 442170 425098 442226
rect 424918 442046 424974 442102
rect 425042 442046 425098 442102
rect 424918 441922 424974 441978
rect 425042 441922 425098 441978
rect 455638 442294 455694 442350
rect 455762 442294 455818 442350
rect 455638 442170 455694 442226
rect 455762 442170 455818 442226
rect 455638 442046 455694 442102
rect 455762 442046 455818 442102
rect 455638 441922 455694 441978
rect 455762 441922 455818 441978
rect 225238 436294 225294 436350
rect 225362 436294 225418 436350
rect 225238 436170 225294 436226
rect 225362 436170 225418 436226
rect 225238 436046 225294 436102
rect 225362 436046 225418 436102
rect 225238 435922 225294 435978
rect 225362 435922 225418 435978
rect 255958 436294 256014 436350
rect 256082 436294 256138 436350
rect 255958 436170 256014 436226
rect 256082 436170 256138 436226
rect 255958 436046 256014 436102
rect 256082 436046 256138 436102
rect 255958 435922 256014 435978
rect 256082 435922 256138 435978
rect 286678 436294 286734 436350
rect 286802 436294 286858 436350
rect 286678 436170 286734 436226
rect 286802 436170 286858 436226
rect 286678 436046 286734 436102
rect 286802 436046 286858 436102
rect 286678 435922 286734 435978
rect 286802 435922 286858 435978
rect 317398 436294 317454 436350
rect 317522 436294 317578 436350
rect 317398 436170 317454 436226
rect 317522 436170 317578 436226
rect 317398 436046 317454 436102
rect 317522 436046 317578 436102
rect 317398 435922 317454 435978
rect 317522 435922 317578 435978
rect 348118 436294 348174 436350
rect 348242 436294 348298 436350
rect 348118 436170 348174 436226
rect 348242 436170 348298 436226
rect 348118 436046 348174 436102
rect 348242 436046 348298 436102
rect 348118 435922 348174 435978
rect 348242 435922 348298 435978
rect 378838 436294 378894 436350
rect 378962 436294 379018 436350
rect 378838 436170 378894 436226
rect 378962 436170 379018 436226
rect 378838 436046 378894 436102
rect 378962 436046 379018 436102
rect 378838 435922 378894 435978
rect 378962 435922 379018 435978
rect 409558 436294 409614 436350
rect 409682 436294 409738 436350
rect 409558 436170 409614 436226
rect 409682 436170 409738 436226
rect 409558 436046 409614 436102
rect 409682 436046 409738 436102
rect 409558 435922 409614 435978
rect 409682 435922 409738 435978
rect 440278 436294 440334 436350
rect 440402 436294 440458 436350
rect 440278 436170 440334 436226
rect 440402 436170 440458 436226
rect 440278 436046 440334 436102
rect 440402 436046 440458 436102
rect 440278 435922 440334 435978
rect 440402 435922 440458 435978
rect 470998 436294 471054 436350
rect 471122 436294 471178 436350
rect 470998 436170 471054 436226
rect 471122 436170 471178 436226
rect 470998 436046 471054 436102
rect 471122 436046 471178 436102
rect 470998 435922 471054 435978
rect 471122 435922 471178 435978
rect 209878 424294 209934 424350
rect 210002 424294 210058 424350
rect 209878 424170 209934 424226
rect 210002 424170 210058 424226
rect 209878 424046 209934 424102
rect 210002 424046 210058 424102
rect 209878 423922 209934 423978
rect 210002 423922 210058 423978
rect 240598 424294 240654 424350
rect 240722 424294 240778 424350
rect 240598 424170 240654 424226
rect 240722 424170 240778 424226
rect 240598 424046 240654 424102
rect 240722 424046 240778 424102
rect 240598 423922 240654 423978
rect 240722 423922 240778 423978
rect 271318 424294 271374 424350
rect 271442 424294 271498 424350
rect 271318 424170 271374 424226
rect 271442 424170 271498 424226
rect 271318 424046 271374 424102
rect 271442 424046 271498 424102
rect 271318 423922 271374 423978
rect 271442 423922 271498 423978
rect 302038 424294 302094 424350
rect 302162 424294 302218 424350
rect 302038 424170 302094 424226
rect 302162 424170 302218 424226
rect 302038 424046 302094 424102
rect 302162 424046 302218 424102
rect 302038 423922 302094 423978
rect 302162 423922 302218 423978
rect 332758 424294 332814 424350
rect 332882 424294 332938 424350
rect 332758 424170 332814 424226
rect 332882 424170 332938 424226
rect 332758 424046 332814 424102
rect 332882 424046 332938 424102
rect 332758 423922 332814 423978
rect 332882 423922 332938 423978
rect 363478 424294 363534 424350
rect 363602 424294 363658 424350
rect 363478 424170 363534 424226
rect 363602 424170 363658 424226
rect 363478 424046 363534 424102
rect 363602 424046 363658 424102
rect 363478 423922 363534 423978
rect 363602 423922 363658 423978
rect 394198 424294 394254 424350
rect 394322 424294 394378 424350
rect 394198 424170 394254 424226
rect 394322 424170 394378 424226
rect 394198 424046 394254 424102
rect 394322 424046 394378 424102
rect 394198 423922 394254 423978
rect 394322 423922 394378 423978
rect 424918 424294 424974 424350
rect 425042 424294 425098 424350
rect 424918 424170 424974 424226
rect 425042 424170 425098 424226
rect 424918 424046 424974 424102
rect 425042 424046 425098 424102
rect 424918 423922 424974 423978
rect 425042 423922 425098 423978
rect 455638 424294 455694 424350
rect 455762 424294 455818 424350
rect 455638 424170 455694 424226
rect 455762 424170 455818 424226
rect 455638 424046 455694 424102
rect 455762 424046 455818 424102
rect 455638 423922 455694 423978
rect 455762 423922 455818 423978
rect 225238 418294 225294 418350
rect 225362 418294 225418 418350
rect 225238 418170 225294 418226
rect 225362 418170 225418 418226
rect 225238 418046 225294 418102
rect 225362 418046 225418 418102
rect 225238 417922 225294 417978
rect 225362 417922 225418 417978
rect 255958 418294 256014 418350
rect 256082 418294 256138 418350
rect 255958 418170 256014 418226
rect 256082 418170 256138 418226
rect 255958 418046 256014 418102
rect 256082 418046 256138 418102
rect 255958 417922 256014 417978
rect 256082 417922 256138 417978
rect 286678 418294 286734 418350
rect 286802 418294 286858 418350
rect 286678 418170 286734 418226
rect 286802 418170 286858 418226
rect 286678 418046 286734 418102
rect 286802 418046 286858 418102
rect 286678 417922 286734 417978
rect 286802 417922 286858 417978
rect 317398 418294 317454 418350
rect 317522 418294 317578 418350
rect 317398 418170 317454 418226
rect 317522 418170 317578 418226
rect 317398 418046 317454 418102
rect 317522 418046 317578 418102
rect 317398 417922 317454 417978
rect 317522 417922 317578 417978
rect 348118 418294 348174 418350
rect 348242 418294 348298 418350
rect 348118 418170 348174 418226
rect 348242 418170 348298 418226
rect 348118 418046 348174 418102
rect 348242 418046 348298 418102
rect 348118 417922 348174 417978
rect 348242 417922 348298 417978
rect 378838 418294 378894 418350
rect 378962 418294 379018 418350
rect 378838 418170 378894 418226
rect 378962 418170 379018 418226
rect 378838 418046 378894 418102
rect 378962 418046 379018 418102
rect 378838 417922 378894 417978
rect 378962 417922 379018 417978
rect 409558 418294 409614 418350
rect 409682 418294 409738 418350
rect 409558 418170 409614 418226
rect 409682 418170 409738 418226
rect 409558 418046 409614 418102
rect 409682 418046 409738 418102
rect 409558 417922 409614 417978
rect 409682 417922 409738 417978
rect 440278 418294 440334 418350
rect 440402 418294 440458 418350
rect 440278 418170 440334 418226
rect 440402 418170 440458 418226
rect 440278 418046 440334 418102
rect 440402 418046 440458 418102
rect 440278 417922 440334 417978
rect 440402 417922 440458 417978
rect 470998 418294 471054 418350
rect 471122 418294 471178 418350
rect 470998 418170 471054 418226
rect 471122 418170 471178 418226
rect 470998 418046 471054 418102
rect 471122 418046 471178 418102
rect 470998 417922 471054 417978
rect 471122 417922 471178 417978
rect 336924 410462 336980 410518
rect 297276 410282 297332 410338
rect 261996 409562 262052 409618
rect 206668 403982 206724 404038
rect 203308 390482 203364 390538
rect 203084 383462 203140 383518
rect 201404 214082 201460 214138
rect 196476 206522 196532 206578
rect 204092 302462 204148 302518
rect 204652 379322 204708 379378
rect 208348 402362 208404 402418
rect 220554 400294 220610 400350
rect 220678 400294 220734 400350
rect 220802 400294 220858 400350
rect 220926 400294 220982 400350
rect 220554 400170 220610 400226
rect 220678 400170 220734 400226
rect 220802 400170 220858 400226
rect 220926 400170 220982 400226
rect 220554 400046 220610 400102
rect 220678 400046 220734 400102
rect 220802 400046 220858 400102
rect 220926 400046 220982 400102
rect 220554 399922 220610 399978
rect 220678 399922 220734 399978
rect 220802 399922 220858 399978
rect 220926 399922 220982 399978
rect 214508 383282 214564 383338
rect 216524 383102 216580 383158
rect 220554 382294 220610 382350
rect 220678 382294 220734 382350
rect 220802 382294 220858 382350
rect 220926 382294 220982 382350
rect 220554 382170 220610 382226
rect 220678 382170 220734 382226
rect 220802 382170 220858 382226
rect 220926 382170 220982 382226
rect 220554 382046 220610 382102
rect 220678 382046 220734 382102
rect 220802 382046 220858 382102
rect 220926 382046 220982 382102
rect 220554 381922 220610 381978
rect 220678 381922 220734 381978
rect 220802 381922 220858 381978
rect 220926 381922 220982 381978
rect 215852 380222 215908 380278
rect 204876 379862 204932 379918
rect 218540 379862 218596 379918
rect 213164 379142 213220 379198
rect 217196 379322 217252 379378
rect 240268 407402 240324 407458
rect 243516 409022 243572 409078
rect 232316 406682 232372 406738
rect 224274 406294 224330 406350
rect 224398 406294 224454 406350
rect 224522 406294 224578 406350
rect 224646 406294 224702 406350
rect 224274 406170 224330 406226
rect 224398 406170 224454 406226
rect 224522 406170 224578 406226
rect 224646 406170 224702 406226
rect 224274 406046 224330 406102
rect 224398 406046 224454 406102
rect 224522 406046 224578 406102
rect 224646 406046 224702 406102
rect 224274 405922 224330 405978
rect 224398 405922 224454 405978
rect 224522 405922 224578 405978
rect 224646 405922 224702 405978
rect 224274 388294 224330 388350
rect 224398 388294 224454 388350
rect 224522 388294 224578 388350
rect 224646 388294 224702 388350
rect 224274 388170 224330 388226
rect 224398 388170 224454 388226
rect 224522 388170 224578 388226
rect 224646 388170 224702 388226
rect 224274 388046 224330 388102
rect 224398 388046 224454 388102
rect 224522 388046 224578 388102
rect 224646 388046 224702 388102
rect 224274 387922 224330 387978
rect 224398 387922 224454 387978
rect 224522 387922 224578 387978
rect 224646 387922 224702 387978
rect 246876 407222 246932 407278
rect 251274 400294 251330 400350
rect 251398 400294 251454 400350
rect 251522 400294 251578 400350
rect 251646 400294 251702 400350
rect 251274 400170 251330 400226
rect 251398 400170 251454 400226
rect 251522 400170 251578 400226
rect 251646 400170 251702 400226
rect 251274 400046 251330 400102
rect 251398 400046 251454 400102
rect 251522 400046 251578 400102
rect 251646 400046 251702 400102
rect 251274 399922 251330 399978
rect 251398 399922 251454 399978
rect 251522 399922 251578 399978
rect 251646 399922 251702 399978
rect 251274 382294 251330 382350
rect 251398 382294 251454 382350
rect 251522 382294 251578 382350
rect 251646 382294 251702 382350
rect 251274 382170 251330 382226
rect 251398 382170 251454 382226
rect 251522 382170 251578 382226
rect 251646 382170 251702 382226
rect 251274 382046 251330 382102
rect 251398 382046 251454 382102
rect 251522 382046 251578 382102
rect 251646 382046 251702 382102
rect 251274 381922 251330 381978
rect 251398 381922 251454 381978
rect 251522 381922 251578 381978
rect 251646 381922 251702 381978
rect 254994 406294 255050 406350
rect 255118 406294 255174 406350
rect 255242 406294 255298 406350
rect 255366 406294 255422 406350
rect 254994 406170 255050 406226
rect 255118 406170 255174 406226
rect 255242 406170 255298 406226
rect 255366 406170 255422 406226
rect 254994 406046 255050 406102
rect 255118 406046 255174 406102
rect 255242 406046 255298 406102
rect 255366 406046 255422 406102
rect 254994 405922 255050 405978
rect 255118 405922 255174 405978
rect 255242 405922 255298 405978
rect 255366 405922 255422 405978
rect 254994 388294 255050 388350
rect 255118 388294 255174 388350
rect 255242 388294 255298 388350
rect 255366 388294 255422 388350
rect 254994 388170 255050 388226
rect 255118 388170 255174 388226
rect 255242 388170 255298 388226
rect 255366 388170 255422 388226
rect 254994 388046 255050 388102
rect 255118 388046 255174 388102
rect 255242 388046 255298 388102
rect 255366 388046 255422 388102
rect 254994 387922 255050 387978
rect 255118 387922 255174 387978
rect 255242 387922 255298 387978
rect 255366 387922 255422 387978
rect 278908 409382 278964 409438
rect 288092 409202 288148 409258
rect 278796 402362 278852 402418
rect 263676 400562 263732 400618
rect 281994 400294 282050 400350
rect 282118 400294 282174 400350
rect 282242 400294 282298 400350
rect 282366 400294 282422 400350
rect 281994 400170 282050 400226
rect 282118 400170 282174 400226
rect 282242 400170 282298 400226
rect 282366 400170 282422 400226
rect 281994 400046 282050 400102
rect 282118 400046 282174 400102
rect 282242 400046 282298 400102
rect 282366 400046 282422 400102
rect 281994 399922 282050 399978
rect 282118 399922 282174 399978
rect 282242 399922 282298 399978
rect 282366 399922 282422 399978
rect 281994 382294 282050 382350
rect 282118 382294 282174 382350
rect 282242 382294 282298 382350
rect 282366 382294 282422 382350
rect 281994 382170 282050 382226
rect 282118 382170 282174 382226
rect 282242 382170 282298 382226
rect 282366 382170 282422 382226
rect 281994 382046 282050 382102
rect 282118 382046 282174 382102
rect 282242 382046 282298 382102
rect 282366 382046 282422 382102
rect 281994 381922 282050 381978
rect 282118 381922 282174 381978
rect 282242 381922 282298 381978
rect 282366 381922 282422 381978
rect 295596 408662 295652 408718
rect 285714 406294 285770 406350
rect 285838 406294 285894 406350
rect 285962 406294 286018 406350
rect 286086 406294 286142 406350
rect 285714 406170 285770 406226
rect 285838 406170 285894 406226
rect 285962 406170 286018 406226
rect 286086 406170 286142 406226
rect 285714 406046 285770 406102
rect 285838 406046 285894 406102
rect 285962 406046 286018 406102
rect 286086 406046 286142 406102
rect 285714 405922 285770 405978
rect 285838 405922 285894 405978
rect 285962 405922 286018 405978
rect 286086 405922 286142 405978
rect 285714 388294 285770 388350
rect 285838 388294 285894 388350
rect 285962 388294 286018 388350
rect 286086 388294 286142 388350
rect 285714 388170 285770 388226
rect 285838 388170 285894 388226
rect 285962 388170 286018 388226
rect 286086 388170 286142 388226
rect 285714 388046 285770 388102
rect 285838 388046 285894 388102
rect 285962 388046 286018 388102
rect 286086 388046 286142 388102
rect 285714 387922 285770 387978
rect 285838 387922 285894 387978
rect 285962 387922 286018 387978
rect 286086 387922 286142 387978
rect 293916 402722 293972 402778
rect 298956 408302 299012 408358
rect 305676 407582 305732 407638
rect 302316 407042 302372 407098
rect 302204 406862 302260 406918
rect 300636 403982 300692 404038
rect 303996 405602 304052 405658
rect 303884 400742 303940 400798
rect 312714 400294 312770 400350
rect 312838 400294 312894 400350
rect 312962 400294 313018 400350
rect 313086 400294 313142 400350
rect 312714 400170 312770 400226
rect 312838 400170 312894 400226
rect 312962 400170 313018 400226
rect 313086 400170 313142 400226
rect 312714 400046 312770 400102
rect 312838 400046 312894 400102
rect 312962 400046 313018 400102
rect 313086 400046 313142 400102
rect 312714 399922 312770 399978
rect 312838 399922 312894 399978
rect 312962 399922 313018 399978
rect 313086 399922 313142 399978
rect 316434 406294 316490 406350
rect 316558 406294 316614 406350
rect 316682 406294 316738 406350
rect 316806 406294 316862 406350
rect 316434 406170 316490 406226
rect 316558 406170 316614 406226
rect 316682 406170 316738 406226
rect 316806 406170 316862 406226
rect 316434 406046 316490 406102
rect 316558 406046 316614 406102
rect 316682 406046 316738 406102
rect 316806 406046 316862 406102
rect 316434 405922 316490 405978
rect 316558 405922 316614 405978
rect 316682 405922 316738 405978
rect 316806 405922 316862 405978
rect 312714 382294 312770 382350
rect 312838 382294 312894 382350
rect 312962 382294 313018 382350
rect 313086 382294 313142 382350
rect 312714 382170 312770 382226
rect 312838 382170 312894 382226
rect 312962 382170 313018 382226
rect 313086 382170 313142 382226
rect 312714 382046 312770 382102
rect 312838 382046 312894 382102
rect 312962 382046 313018 382102
rect 313086 382046 313142 382102
rect 312714 381922 312770 381978
rect 312838 381922 312894 381978
rect 312962 381922 313018 381978
rect 313086 381922 313142 381978
rect 313404 395522 313460 395578
rect 316434 388294 316490 388350
rect 316558 388294 316614 388350
rect 316682 388294 316738 388350
rect 316806 388294 316862 388350
rect 316434 388170 316490 388226
rect 316558 388170 316614 388226
rect 316682 388170 316738 388226
rect 316806 388170 316862 388226
rect 316434 388046 316490 388102
rect 316558 388046 316614 388102
rect 316682 388046 316738 388102
rect 316806 388046 316862 388102
rect 316434 387922 316490 387978
rect 316558 387922 316614 387978
rect 316682 387922 316738 387978
rect 316806 387922 316862 387978
rect 317436 387242 317492 387298
rect 215180 378962 215236 379018
rect 213836 378782 213892 378838
rect 230598 370294 230654 370350
rect 230722 370294 230778 370350
rect 230598 370170 230654 370226
rect 230722 370170 230778 370226
rect 230598 370046 230654 370102
rect 230722 370046 230778 370102
rect 230598 369922 230654 369978
rect 230722 369922 230778 369978
rect 261318 370294 261374 370350
rect 261442 370294 261498 370350
rect 261318 370170 261374 370226
rect 261442 370170 261498 370226
rect 261318 370046 261374 370102
rect 261442 370046 261498 370102
rect 261318 369922 261374 369978
rect 261442 369922 261498 369978
rect 292038 370294 292094 370350
rect 292162 370294 292218 370350
rect 292038 370170 292094 370226
rect 292162 370170 292218 370226
rect 292038 370046 292094 370102
rect 292162 370046 292218 370102
rect 292038 369922 292094 369978
rect 292162 369922 292218 369978
rect 322758 370294 322814 370350
rect 322882 370294 322938 370350
rect 322758 370170 322814 370226
rect 322882 370170 322938 370226
rect 322758 370046 322814 370102
rect 322882 370046 322938 370102
rect 322758 369922 322814 369978
rect 322882 369922 322938 369978
rect 215238 364294 215294 364350
rect 215362 364294 215418 364350
rect 215238 364170 215294 364226
rect 215362 364170 215418 364226
rect 215238 364046 215294 364102
rect 215362 364046 215418 364102
rect 215238 363922 215294 363978
rect 215362 363922 215418 363978
rect 245958 364294 246014 364350
rect 246082 364294 246138 364350
rect 245958 364170 246014 364226
rect 246082 364170 246138 364226
rect 245958 364046 246014 364102
rect 246082 364046 246138 364102
rect 245958 363922 246014 363978
rect 246082 363922 246138 363978
rect 276678 364294 276734 364350
rect 276802 364294 276858 364350
rect 276678 364170 276734 364226
rect 276802 364170 276858 364226
rect 276678 364046 276734 364102
rect 276802 364046 276858 364102
rect 276678 363922 276734 363978
rect 276802 363922 276858 363978
rect 307398 364294 307454 364350
rect 307522 364294 307578 364350
rect 307398 364170 307454 364226
rect 307522 364170 307578 364226
rect 307398 364046 307454 364102
rect 307522 364046 307578 364102
rect 307398 363922 307454 363978
rect 307522 363922 307578 363978
rect 327404 360782 327460 360838
rect 328412 379682 328468 379738
rect 230598 352294 230654 352350
rect 230722 352294 230778 352350
rect 230598 352170 230654 352226
rect 230722 352170 230778 352226
rect 230598 352046 230654 352102
rect 230722 352046 230778 352102
rect 230598 351922 230654 351978
rect 230722 351922 230778 351978
rect 261318 352294 261374 352350
rect 261442 352294 261498 352350
rect 261318 352170 261374 352226
rect 261442 352170 261498 352226
rect 261318 352046 261374 352102
rect 261442 352046 261498 352102
rect 261318 351922 261374 351978
rect 261442 351922 261498 351978
rect 292038 352294 292094 352350
rect 292162 352294 292218 352350
rect 292038 352170 292094 352226
rect 292162 352170 292218 352226
rect 292038 352046 292094 352102
rect 292162 352046 292218 352102
rect 292038 351922 292094 351978
rect 292162 351922 292218 351978
rect 322758 352294 322814 352350
rect 322882 352294 322938 352350
rect 322758 352170 322814 352226
rect 322882 352170 322938 352226
rect 322758 352046 322814 352102
rect 322882 352046 322938 352102
rect 322758 351922 322814 351978
rect 322882 351922 322938 351978
rect 215238 346294 215294 346350
rect 215362 346294 215418 346350
rect 215238 346170 215294 346226
rect 215362 346170 215418 346226
rect 215238 346046 215294 346102
rect 215362 346046 215418 346102
rect 215238 345922 215294 345978
rect 215362 345922 215418 345978
rect 245958 346294 246014 346350
rect 246082 346294 246138 346350
rect 245958 346170 246014 346226
rect 246082 346170 246138 346226
rect 245958 346046 246014 346102
rect 246082 346046 246138 346102
rect 245958 345922 246014 345978
rect 246082 345922 246138 345978
rect 276678 346294 276734 346350
rect 276802 346294 276858 346350
rect 276678 346170 276734 346226
rect 276802 346170 276858 346226
rect 276678 346046 276734 346102
rect 276802 346046 276858 346102
rect 276678 345922 276734 345978
rect 276802 345922 276858 345978
rect 307398 346294 307454 346350
rect 307522 346294 307578 346350
rect 307398 346170 307454 346226
rect 307522 346170 307578 346226
rect 307398 346046 307454 346102
rect 307522 346046 307578 346102
rect 307398 345922 307454 345978
rect 307522 345922 307578 345978
rect 230598 334294 230654 334350
rect 230722 334294 230778 334350
rect 230598 334170 230654 334226
rect 230722 334170 230778 334226
rect 230598 334046 230654 334102
rect 230722 334046 230778 334102
rect 230598 333922 230654 333978
rect 230722 333922 230778 333978
rect 261318 334294 261374 334350
rect 261442 334294 261498 334350
rect 261318 334170 261374 334226
rect 261442 334170 261498 334226
rect 261318 334046 261374 334102
rect 261442 334046 261498 334102
rect 261318 333922 261374 333978
rect 261442 333922 261498 333978
rect 292038 334294 292094 334350
rect 292162 334294 292218 334350
rect 292038 334170 292094 334226
rect 292162 334170 292218 334226
rect 292038 334046 292094 334102
rect 292162 334046 292218 334102
rect 292038 333922 292094 333978
rect 292162 333922 292218 333978
rect 322758 334294 322814 334350
rect 322882 334294 322938 334350
rect 322758 334170 322814 334226
rect 322882 334170 322938 334226
rect 322758 334046 322814 334102
rect 322882 334046 322938 334102
rect 322758 333922 322814 333978
rect 322882 333922 322938 333978
rect 215238 328294 215294 328350
rect 215362 328294 215418 328350
rect 215238 328170 215294 328226
rect 215362 328170 215418 328226
rect 215238 328046 215294 328102
rect 215362 328046 215418 328102
rect 215238 327922 215294 327978
rect 215362 327922 215418 327978
rect 245958 328294 246014 328350
rect 246082 328294 246138 328350
rect 245958 328170 246014 328226
rect 246082 328170 246138 328226
rect 245958 328046 246014 328102
rect 246082 328046 246138 328102
rect 245958 327922 246014 327978
rect 246082 327922 246138 327978
rect 276678 328294 276734 328350
rect 276802 328294 276858 328350
rect 276678 328170 276734 328226
rect 276802 328170 276858 328226
rect 276678 328046 276734 328102
rect 276802 328046 276858 328102
rect 276678 327922 276734 327978
rect 276802 327922 276858 327978
rect 307398 328294 307454 328350
rect 307522 328294 307578 328350
rect 307398 328170 307454 328226
rect 307522 328170 307578 328226
rect 307398 328046 307454 328102
rect 307522 328046 307578 328102
rect 307398 327922 307454 327978
rect 307522 327922 307578 327978
rect 230598 316294 230654 316350
rect 230722 316294 230778 316350
rect 230598 316170 230654 316226
rect 230722 316170 230778 316226
rect 230598 316046 230654 316102
rect 230722 316046 230778 316102
rect 230598 315922 230654 315978
rect 230722 315922 230778 315978
rect 261318 316294 261374 316350
rect 261442 316294 261498 316350
rect 261318 316170 261374 316226
rect 261442 316170 261498 316226
rect 261318 316046 261374 316102
rect 261442 316046 261498 316102
rect 261318 315922 261374 315978
rect 261442 315922 261498 315978
rect 292038 316294 292094 316350
rect 292162 316294 292218 316350
rect 292038 316170 292094 316226
rect 292162 316170 292218 316226
rect 292038 316046 292094 316102
rect 292162 316046 292218 316102
rect 292038 315922 292094 315978
rect 292162 315922 292218 315978
rect 322758 316294 322814 316350
rect 322882 316294 322938 316350
rect 322758 316170 322814 316226
rect 322882 316170 322938 316226
rect 322758 316046 322814 316102
rect 322882 316046 322938 316102
rect 322758 315922 322814 315978
rect 322882 315922 322938 315978
rect 328076 311642 328132 311698
rect 215238 310294 215294 310350
rect 215362 310294 215418 310350
rect 215238 310170 215294 310226
rect 215362 310170 215418 310226
rect 215238 310046 215294 310102
rect 215362 310046 215418 310102
rect 215238 309922 215294 309978
rect 215362 309922 215418 309978
rect 245958 310294 246014 310350
rect 246082 310294 246138 310350
rect 245958 310170 246014 310226
rect 246082 310170 246138 310226
rect 245958 310046 246014 310102
rect 246082 310046 246138 310102
rect 245958 309922 246014 309978
rect 246082 309922 246138 309978
rect 276678 310294 276734 310350
rect 276802 310294 276858 310350
rect 276678 310170 276734 310226
rect 276802 310170 276858 310226
rect 276678 310046 276734 310102
rect 276802 310046 276858 310102
rect 276678 309922 276734 309978
rect 276802 309922 276858 309978
rect 307398 310294 307454 310350
rect 307522 310294 307578 310350
rect 307398 310170 307454 310226
rect 307522 310170 307578 310226
rect 307398 310046 307454 310102
rect 307522 310046 307578 310102
rect 307398 309922 307454 309978
rect 307522 309922 307578 309978
rect 230598 298294 230654 298350
rect 230722 298294 230778 298350
rect 230598 298170 230654 298226
rect 230722 298170 230778 298226
rect 230598 298046 230654 298102
rect 230722 298046 230778 298102
rect 230598 297922 230654 297978
rect 230722 297922 230778 297978
rect 261318 298294 261374 298350
rect 261442 298294 261498 298350
rect 261318 298170 261374 298226
rect 261442 298170 261498 298226
rect 261318 298046 261374 298102
rect 261442 298046 261498 298102
rect 261318 297922 261374 297978
rect 261442 297922 261498 297978
rect 292038 298294 292094 298350
rect 292162 298294 292218 298350
rect 292038 298170 292094 298226
rect 292162 298170 292218 298226
rect 292038 298046 292094 298102
rect 292162 298046 292218 298102
rect 292038 297922 292094 297978
rect 292162 297922 292218 297978
rect 322758 298294 322814 298350
rect 322882 298294 322938 298350
rect 322758 298170 322814 298226
rect 322882 298170 322938 298226
rect 322758 298046 322814 298102
rect 322882 298046 322938 298102
rect 322758 297922 322814 297978
rect 322882 297922 322938 297978
rect 215238 292294 215294 292350
rect 215362 292294 215418 292350
rect 215238 292170 215294 292226
rect 215362 292170 215418 292226
rect 215238 292046 215294 292102
rect 215362 292046 215418 292102
rect 215238 291922 215294 291978
rect 215362 291922 215418 291978
rect 245958 292294 246014 292350
rect 246082 292294 246138 292350
rect 245958 292170 246014 292226
rect 246082 292170 246138 292226
rect 245958 292046 246014 292102
rect 246082 292046 246138 292102
rect 245958 291922 246014 291978
rect 246082 291922 246138 291978
rect 276678 292294 276734 292350
rect 276802 292294 276858 292350
rect 276678 292170 276734 292226
rect 276802 292170 276858 292226
rect 276678 292046 276734 292102
rect 276802 292046 276858 292102
rect 276678 291922 276734 291978
rect 276802 291922 276858 291978
rect 307398 292294 307454 292350
rect 307522 292294 307578 292350
rect 307398 292170 307454 292226
rect 307522 292170 307578 292226
rect 307398 292046 307454 292102
rect 307522 292046 307578 292102
rect 307398 291922 307454 291978
rect 307522 291922 307578 291978
rect 230598 280294 230654 280350
rect 230722 280294 230778 280350
rect 230598 280170 230654 280226
rect 230722 280170 230778 280226
rect 230598 280046 230654 280102
rect 230722 280046 230778 280102
rect 230598 279922 230654 279978
rect 230722 279922 230778 279978
rect 261318 280294 261374 280350
rect 261442 280294 261498 280350
rect 261318 280170 261374 280226
rect 261442 280170 261498 280226
rect 261318 280046 261374 280102
rect 261442 280046 261498 280102
rect 261318 279922 261374 279978
rect 261442 279922 261498 279978
rect 292038 280294 292094 280350
rect 292162 280294 292218 280350
rect 292038 280170 292094 280226
rect 292162 280170 292218 280226
rect 292038 280046 292094 280102
rect 292162 280046 292218 280102
rect 292038 279922 292094 279978
rect 292162 279922 292218 279978
rect 322758 280294 322814 280350
rect 322882 280294 322938 280350
rect 322758 280170 322814 280226
rect 322882 280170 322938 280226
rect 322758 280046 322814 280102
rect 322882 280046 322938 280102
rect 322758 279922 322814 279978
rect 322882 279922 322938 279978
rect 215238 274294 215294 274350
rect 215362 274294 215418 274350
rect 215238 274170 215294 274226
rect 215362 274170 215418 274226
rect 215238 274046 215294 274102
rect 215362 274046 215418 274102
rect 215238 273922 215294 273978
rect 215362 273922 215418 273978
rect 245958 274294 246014 274350
rect 246082 274294 246138 274350
rect 245958 274170 246014 274226
rect 246082 274170 246138 274226
rect 245958 274046 246014 274102
rect 246082 274046 246138 274102
rect 245958 273922 246014 273978
rect 246082 273922 246138 273978
rect 276678 274294 276734 274350
rect 276802 274294 276858 274350
rect 276678 274170 276734 274226
rect 276802 274170 276858 274226
rect 276678 274046 276734 274102
rect 276802 274046 276858 274102
rect 276678 273922 276734 273978
rect 276802 273922 276858 273978
rect 307398 274294 307454 274350
rect 307522 274294 307578 274350
rect 307398 274170 307454 274226
rect 307522 274170 307578 274226
rect 307398 274046 307454 274102
rect 307522 274046 307578 274102
rect 307398 273922 307454 273978
rect 307522 273922 307578 273978
rect 230598 262294 230654 262350
rect 230722 262294 230778 262350
rect 230598 262170 230654 262226
rect 230722 262170 230778 262226
rect 230598 262046 230654 262102
rect 230722 262046 230778 262102
rect 230598 261922 230654 261978
rect 230722 261922 230778 261978
rect 261318 262294 261374 262350
rect 261442 262294 261498 262350
rect 261318 262170 261374 262226
rect 261442 262170 261498 262226
rect 261318 262046 261374 262102
rect 261442 262046 261498 262102
rect 261318 261922 261374 261978
rect 261442 261922 261498 261978
rect 292038 262294 292094 262350
rect 292162 262294 292218 262350
rect 292038 262170 292094 262226
rect 292162 262170 292218 262226
rect 292038 262046 292094 262102
rect 292162 262046 292218 262102
rect 292038 261922 292094 261978
rect 292162 261922 292218 261978
rect 322758 262294 322814 262350
rect 322882 262294 322938 262350
rect 322758 262170 322814 262226
rect 322882 262170 322938 262226
rect 322758 262046 322814 262102
rect 322882 262046 322938 262102
rect 322758 261922 322814 261978
rect 322882 261922 322938 261978
rect 327964 260342 328020 260398
rect 215238 256294 215294 256350
rect 215362 256294 215418 256350
rect 215238 256170 215294 256226
rect 215362 256170 215418 256226
rect 215238 256046 215294 256102
rect 215362 256046 215418 256102
rect 215238 255922 215294 255978
rect 215362 255922 215418 255978
rect 245958 256294 246014 256350
rect 246082 256294 246138 256350
rect 245958 256170 246014 256226
rect 246082 256170 246138 256226
rect 245958 256046 246014 256102
rect 246082 256046 246138 256102
rect 245958 255922 246014 255978
rect 246082 255922 246138 255978
rect 276678 256294 276734 256350
rect 276802 256294 276858 256350
rect 276678 256170 276734 256226
rect 276802 256170 276858 256226
rect 276678 256046 276734 256102
rect 276802 256046 276858 256102
rect 276678 255922 276734 255978
rect 276802 255922 276858 255978
rect 307398 256294 307454 256350
rect 307522 256294 307578 256350
rect 307398 256170 307454 256226
rect 307522 256170 307578 256226
rect 307398 256046 307454 256102
rect 307522 256046 307578 256102
rect 307398 255922 307454 255978
rect 307522 255922 307578 255978
rect 327404 248102 327460 248158
rect 230598 244294 230654 244350
rect 230722 244294 230778 244350
rect 230598 244170 230654 244226
rect 230722 244170 230778 244226
rect 230598 244046 230654 244102
rect 230722 244046 230778 244102
rect 230598 243922 230654 243978
rect 230722 243922 230778 243978
rect 261318 244294 261374 244350
rect 261442 244294 261498 244350
rect 261318 244170 261374 244226
rect 261442 244170 261498 244226
rect 261318 244046 261374 244102
rect 261442 244046 261498 244102
rect 261318 243922 261374 243978
rect 261442 243922 261498 243978
rect 292038 244294 292094 244350
rect 292162 244294 292218 244350
rect 292038 244170 292094 244226
rect 292162 244170 292218 244226
rect 292038 244046 292094 244102
rect 292162 244046 292218 244102
rect 292038 243922 292094 243978
rect 292162 243922 292218 243978
rect 322758 244294 322814 244350
rect 322882 244294 322938 244350
rect 322758 244170 322814 244226
rect 322882 244170 322938 244226
rect 322758 244046 322814 244102
rect 322882 244046 322938 244102
rect 322758 243922 322814 243978
rect 322882 243922 322938 243978
rect 326732 240902 326788 240958
rect 326620 240722 326676 240778
rect 220554 238294 220610 238350
rect 220678 238294 220734 238350
rect 220802 238294 220858 238350
rect 220926 238294 220982 238350
rect 220554 238170 220610 238226
rect 220678 238170 220734 238226
rect 220802 238170 220858 238226
rect 220926 238170 220982 238226
rect 220554 238046 220610 238102
rect 220678 238046 220734 238102
rect 220802 238046 220858 238102
rect 220926 238046 220982 238102
rect 220554 237922 220610 237978
rect 220678 237922 220734 237978
rect 220802 237922 220858 237978
rect 220926 237922 220982 237978
rect 220554 220294 220610 220350
rect 220678 220294 220734 220350
rect 220802 220294 220858 220350
rect 220926 220294 220982 220350
rect 220554 220170 220610 220226
rect 220678 220170 220734 220226
rect 220802 220170 220858 220226
rect 220926 220170 220982 220226
rect 220554 220046 220610 220102
rect 220678 220046 220734 220102
rect 220802 220046 220858 220102
rect 220926 220046 220982 220102
rect 203084 205802 203140 205858
rect 220554 219922 220610 219978
rect 220678 219922 220734 219978
rect 220802 219922 220858 219978
rect 220926 219922 220982 219978
rect 251274 238294 251330 238350
rect 251398 238294 251454 238350
rect 251522 238294 251578 238350
rect 251646 238294 251702 238350
rect 251274 238170 251330 238226
rect 251398 238170 251454 238226
rect 251522 238170 251578 238226
rect 251646 238170 251702 238226
rect 251274 238046 251330 238102
rect 251398 238046 251454 238102
rect 251522 238046 251578 238102
rect 251646 238046 251702 238102
rect 251274 237922 251330 237978
rect 251398 237922 251454 237978
rect 251522 237922 251578 237978
rect 251646 237922 251702 237978
rect 235116 237132 235172 237178
rect 235116 237122 235172 237132
rect 224274 226294 224330 226350
rect 224398 226294 224454 226350
rect 224522 226294 224578 226350
rect 224646 226294 224702 226350
rect 224274 226170 224330 226226
rect 224398 226170 224454 226226
rect 224522 226170 224578 226226
rect 224646 226170 224702 226226
rect 224274 226046 224330 226102
rect 224398 226046 224454 226102
rect 224522 226046 224578 226102
rect 224646 226046 224702 226102
rect 224274 225922 224330 225978
rect 224398 225922 224454 225978
rect 224522 225922 224578 225978
rect 224646 225922 224702 225978
rect 224274 208294 224330 208350
rect 224398 208294 224454 208350
rect 224522 208294 224578 208350
rect 224646 208294 224702 208350
rect 224274 208170 224330 208226
rect 224398 208170 224454 208226
rect 224522 208170 224578 208226
rect 224646 208170 224702 208226
rect 224274 208046 224330 208102
rect 224398 208046 224454 208102
rect 224522 208046 224578 208102
rect 224646 208046 224702 208102
rect 224274 207922 224330 207978
rect 224398 207922 224454 207978
rect 224522 207922 224578 207978
rect 224646 207922 224702 207978
rect 234220 236942 234276 236998
rect 251274 220294 251330 220350
rect 251398 220294 251454 220350
rect 251522 220294 251578 220350
rect 251646 220294 251702 220350
rect 251274 220170 251330 220226
rect 251398 220170 251454 220226
rect 251522 220170 251578 220226
rect 251646 220170 251702 220226
rect 251274 220046 251330 220102
rect 251398 220046 251454 220102
rect 251522 220046 251578 220102
rect 251646 220046 251702 220102
rect 251274 219922 251330 219978
rect 251398 219922 251454 219978
rect 251522 219922 251578 219978
rect 251646 219922 251702 219978
rect 233436 207422 233492 207478
rect 231756 206522 231812 206578
rect 267148 237122 267204 237178
rect 254994 226294 255050 226350
rect 255118 226294 255174 226350
rect 255242 226294 255298 226350
rect 255366 226294 255422 226350
rect 254994 226170 255050 226226
rect 255118 226170 255174 226226
rect 255242 226170 255298 226226
rect 255366 226170 255422 226226
rect 254994 226046 255050 226102
rect 255118 226046 255174 226102
rect 255242 226046 255298 226102
rect 255366 226046 255422 226102
rect 254994 225922 255050 225978
rect 255118 225922 255174 225978
rect 255242 225922 255298 225978
rect 255366 225922 255422 225978
rect 254994 208294 255050 208350
rect 255118 208294 255174 208350
rect 255242 208294 255298 208350
rect 255366 208294 255422 208350
rect 254994 208170 255050 208226
rect 255118 208170 255174 208226
rect 255242 208170 255298 208226
rect 255366 208170 255422 208226
rect 254994 208046 255050 208102
rect 255118 208046 255174 208102
rect 255242 208046 255298 208102
rect 255366 208046 255422 208102
rect 254994 207922 255050 207978
rect 255118 207922 255174 207978
rect 255242 207922 255298 207978
rect 255366 207922 255422 207978
rect 265244 206522 265300 206578
rect 266812 206162 266868 206218
rect 265356 204362 265412 204418
rect 254492 204182 254548 204238
rect 226716 204002 226772 204058
rect 44518 202294 44574 202350
rect 44642 202294 44698 202350
rect 44518 202170 44574 202226
rect 44642 202170 44698 202226
rect 44518 202046 44574 202102
rect 44642 202046 44698 202102
rect 44518 201922 44574 201978
rect 44642 201922 44698 201978
rect 75238 202294 75294 202350
rect 75362 202294 75418 202350
rect 75238 202170 75294 202226
rect 75362 202170 75418 202226
rect 75238 202046 75294 202102
rect 75362 202046 75418 202102
rect 75238 201922 75294 201978
rect 75362 201922 75418 201978
rect 105958 202294 106014 202350
rect 106082 202294 106138 202350
rect 105958 202170 106014 202226
rect 106082 202170 106138 202226
rect 105958 202046 106014 202102
rect 106082 202046 106138 202102
rect 105958 201922 106014 201978
rect 106082 201922 106138 201978
rect 136678 202294 136734 202350
rect 136802 202294 136858 202350
rect 136678 202170 136734 202226
rect 136802 202170 136858 202226
rect 136678 202046 136734 202102
rect 136802 202046 136858 202102
rect 136678 201922 136734 201978
rect 136802 201922 136858 201978
rect 167398 202294 167454 202350
rect 167522 202294 167578 202350
rect 167398 202170 167454 202226
rect 167522 202170 167578 202226
rect 167398 202046 167454 202102
rect 167522 202046 167578 202102
rect 167398 201922 167454 201978
rect 167522 201922 167578 201978
rect 198118 202294 198174 202350
rect 198242 202294 198298 202350
rect 198118 202170 198174 202226
rect 198242 202170 198298 202226
rect 198118 202046 198174 202102
rect 198242 202046 198298 202102
rect 198118 201922 198174 201978
rect 198242 201922 198298 201978
rect 228838 202294 228894 202350
rect 228962 202294 229018 202350
rect 228838 202170 228894 202226
rect 228962 202170 229018 202226
rect 228838 202046 228894 202102
rect 228962 202046 229018 202102
rect 228838 201922 228894 201978
rect 228962 201922 229018 201978
rect 259558 202294 259614 202350
rect 259682 202294 259738 202350
rect 259558 202170 259614 202226
rect 259682 202170 259738 202226
rect 259558 202046 259614 202102
rect 259682 202046 259738 202102
rect 259558 201922 259614 201978
rect 259682 201922 259738 201978
rect 59878 190294 59934 190350
rect 60002 190294 60058 190350
rect 59878 190170 59934 190226
rect 60002 190170 60058 190226
rect 59878 190046 59934 190102
rect 60002 190046 60058 190102
rect 59878 189922 59934 189978
rect 60002 189922 60058 189978
rect 90598 190294 90654 190350
rect 90722 190294 90778 190350
rect 90598 190170 90654 190226
rect 90722 190170 90778 190226
rect 90598 190046 90654 190102
rect 90722 190046 90778 190102
rect 90598 189922 90654 189978
rect 90722 189922 90778 189978
rect 121318 190294 121374 190350
rect 121442 190294 121498 190350
rect 121318 190170 121374 190226
rect 121442 190170 121498 190226
rect 121318 190046 121374 190102
rect 121442 190046 121498 190102
rect 121318 189922 121374 189978
rect 121442 189922 121498 189978
rect 152038 190294 152094 190350
rect 152162 190294 152218 190350
rect 152038 190170 152094 190226
rect 152162 190170 152218 190226
rect 152038 190046 152094 190102
rect 152162 190046 152218 190102
rect 152038 189922 152094 189978
rect 152162 189922 152218 189978
rect 182758 190294 182814 190350
rect 182882 190294 182938 190350
rect 182758 190170 182814 190226
rect 182882 190170 182938 190226
rect 182758 190046 182814 190102
rect 182882 190046 182938 190102
rect 182758 189922 182814 189978
rect 182882 189922 182938 189978
rect 213478 190294 213534 190350
rect 213602 190294 213658 190350
rect 213478 190170 213534 190226
rect 213602 190170 213658 190226
rect 213478 190046 213534 190102
rect 213602 190046 213658 190102
rect 213478 189922 213534 189978
rect 213602 189922 213658 189978
rect 244198 190294 244254 190350
rect 244322 190294 244378 190350
rect 244198 190170 244254 190226
rect 244322 190170 244378 190226
rect 244198 190046 244254 190102
rect 244322 190046 244378 190102
rect 244198 189922 244254 189978
rect 244322 189922 244378 189978
rect 44518 184294 44574 184350
rect 44642 184294 44698 184350
rect 44518 184170 44574 184226
rect 44642 184170 44698 184226
rect 44518 184046 44574 184102
rect 44642 184046 44698 184102
rect 44518 183922 44574 183978
rect 44642 183922 44698 183978
rect 75238 184294 75294 184350
rect 75362 184294 75418 184350
rect 75238 184170 75294 184226
rect 75362 184170 75418 184226
rect 75238 184046 75294 184102
rect 75362 184046 75418 184102
rect 75238 183922 75294 183978
rect 75362 183922 75418 183978
rect 105958 184294 106014 184350
rect 106082 184294 106138 184350
rect 105958 184170 106014 184226
rect 106082 184170 106138 184226
rect 105958 184046 106014 184102
rect 106082 184046 106138 184102
rect 105958 183922 106014 183978
rect 106082 183922 106138 183978
rect 136678 184294 136734 184350
rect 136802 184294 136858 184350
rect 136678 184170 136734 184226
rect 136802 184170 136858 184226
rect 136678 184046 136734 184102
rect 136802 184046 136858 184102
rect 136678 183922 136734 183978
rect 136802 183922 136858 183978
rect 167398 184294 167454 184350
rect 167522 184294 167578 184350
rect 167398 184170 167454 184226
rect 167522 184170 167578 184226
rect 167398 184046 167454 184102
rect 167522 184046 167578 184102
rect 167398 183922 167454 183978
rect 167522 183922 167578 183978
rect 198118 184294 198174 184350
rect 198242 184294 198298 184350
rect 198118 184170 198174 184226
rect 198242 184170 198298 184226
rect 198118 184046 198174 184102
rect 198242 184046 198298 184102
rect 198118 183922 198174 183978
rect 198242 183922 198298 183978
rect 228838 184294 228894 184350
rect 228962 184294 229018 184350
rect 228838 184170 228894 184226
rect 228962 184170 229018 184226
rect 228838 184046 228894 184102
rect 228962 184046 229018 184102
rect 228838 183922 228894 183978
rect 228962 183922 229018 183978
rect 259558 184294 259614 184350
rect 259682 184294 259738 184350
rect 259558 184170 259614 184226
rect 259682 184170 259738 184226
rect 259558 184046 259614 184102
rect 259682 184046 259738 184102
rect 259558 183922 259614 183978
rect 259682 183922 259738 183978
rect 59878 172294 59934 172350
rect 60002 172294 60058 172350
rect 59878 172170 59934 172226
rect 60002 172170 60058 172226
rect 59878 172046 59934 172102
rect 60002 172046 60058 172102
rect 59878 171922 59934 171978
rect 60002 171922 60058 171978
rect 90598 172294 90654 172350
rect 90722 172294 90778 172350
rect 90598 172170 90654 172226
rect 90722 172170 90778 172226
rect 90598 172046 90654 172102
rect 90722 172046 90778 172102
rect 90598 171922 90654 171978
rect 90722 171922 90778 171978
rect 121318 172294 121374 172350
rect 121442 172294 121498 172350
rect 121318 172170 121374 172226
rect 121442 172170 121498 172226
rect 121318 172046 121374 172102
rect 121442 172046 121498 172102
rect 121318 171922 121374 171978
rect 121442 171922 121498 171978
rect 152038 172294 152094 172350
rect 152162 172294 152218 172350
rect 152038 172170 152094 172226
rect 152162 172170 152218 172226
rect 152038 172046 152094 172102
rect 152162 172046 152218 172102
rect 152038 171922 152094 171978
rect 152162 171922 152218 171978
rect 182758 172294 182814 172350
rect 182882 172294 182938 172350
rect 182758 172170 182814 172226
rect 182882 172170 182938 172226
rect 182758 172046 182814 172102
rect 182882 172046 182938 172102
rect 182758 171922 182814 171978
rect 182882 171922 182938 171978
rect 213478 172294 213534 172350
rect 213602 172294 213658 172350
rect 213478 172170 213534 172226
rect 213602 172170 213658 172226
rect 213478 172046 213534 172102
rect 213602 172046 213658 172102
rect 213478 171922 213534 171978
rect 213602 171922 213658 171978
rect 244198 172294 244254 172350
rect 244322 172294 244378 172350
rect 244198 172170 244254 172226
rect 244322 172170 244378 172226
rect 244198 172046 244254 172102
rect 244322 172046 244378 172102
rect 244198 171922 244254 171978
rect 244322 171922 244378 171978
rect 44518 166294 44574 166350
rect 44642 166294 44698 166350
rect 44518 166170 44574 166226
rect 44642 166170 44698 166226
rect 44518 166046 44574 166102
rect 44642 166046 44698 166102
rect 44518 165922 44574 165978
rect 44642 165922 44698 165978
rect 75238 166294 75294 166350
rect 75362 166294 75418 166350
rect 75238 166170 75294 166226
rect 75362 166170 75418 166226
rect 75238 166046 75294 166102
rect 75362 166046 75418 166102
rect 75238 165922 75294 165978
rect 75362 165922 75418 165978
rect 105958 166294 106014 166350
rect 106082 166294 106138 166350
rect 105958 166170 106014 166226
rect 106082 166170 106138 166226
rect 105958 166046 106014 166102
rect 106082 166046 106138 166102
rect 105958 165922 106014 165978
rect 106082 165922 106138 165978
rect 136678 166294 136734 166350
rect 136802 166294 136858 166350
rect 136678 166170 136734 166226
rect 136802 166170 136858 166226
rect 136678 166046 136734 166102
rect 136802 166046 136858 166102
rect 136678 165922 136734 165978
rect 136802 165922 136858 165978
rect 167398 166294 167454 166350
rect 167522 166294 167578 166350
rect 167398 166170 167454 166226
rect 167522 166170 167578 166226
rect 167398 166046 167454 166102
rect 167522 166046 167578 166102
rect 167398 165922 167454 165978
rect 167522 165922 167578 165978
rect 198118 166294 198174 166350
rect 198242 166294 198298 166350
rect 198118 166170 198174 166226
rect 198242 166170 198298 166226
rect 198118 166046 198174 166102
rect 198242 166046 198298 166102
rect 198118 165922 198174 165978
rect 198242 165922 198298 165978
rect 228838 166294 228894 166350
rect 228962 166294 229018 166350
rect 228838 166170 228894 166226
rect 228962 166170 229018 166226
rect 228838 166046 228894 166102
rect 228962 166046 229018 166102
rect 228838 165922 228894 165978
rect 228962 165922 229018 165978
rect 259558 166294 259614 166350
rect 259682 166294 259738 166350
rect 259558 166170 259614 166226
rect 259682 166170 259738 166226
rect 259558 166046 259614 166102
rect 259682 166046 259738 166102
rect 259558 165922 259614 165978
rect 259682 165922 259738 165978
rect 59878 154294 59934 154350
rect 60002 154294 60058 154350
rect 59878 154170 59934 154226
rect 60002 154170 60058 154226
rect 59878 154046 59934 154102
rect 60002 154046 60058 154102
rect 59878 153922 59934 153978
rect 60002 153922 60058 153978
rect 90598 154294 90654 154350
rect 90722 154294 90778 154350
rect 90598 154170 90654 154226
rect 90722 154170 90778 154226
rect 90598 154046 90654 154102
rect 90722 154046 90778 154102
rect 90598 153922 90654 153978
rect 90722 153922 90778 153978
rect 121318 154294 121374 154350
rect 121442 154294 121498 154350
rect 121318 154170 121374 154226
rect 121442 154170 121498 154226
rect 121318 154046 121374 154102
rect 121442 154046 121498 154102
rect 121318 153922 121374 153978
rect 121442 153922 121498 153978
rect 152038 154294 152094 154350
rect 152162 154294 152218 154350
rect 152038 154170 152094 154226
rect 152162 154170 152218 154226
rect 152038 154046 152094 154102
rect 152162 154046 152218 154102
rect 152038 153922 152094 153978
rect 152162 153922 152218 153978
rect 182758 154294 182814 154350
rect 182882 154294 182938 154350
rect 182758 154170 182814 154226
rect 182882 154170 182938 154226
rect 182758 154046 182814 154102
rect 182882 154046 182938 154102
rect 182758 153922 182814 153978
rect 182882 153922 182938 153978
rect 213478 154294 213534 154350
rect 213602 154294 213658 154350
rect 213478 154170 213534 154226
rect 213602 154170 213658 154226
rect 213478 154046 213534 154102
rect 213602 154046 213658 154102
rect 213478 153922 213534 153978
rect 213602 153922 213658 153978
rect 244198 154294 244254 154350
rect 244322 154294 244378 154350
rect 244198 154170 244254 154226
rect 244322 154170 244378 154226
rect 244198 154046 244254 154102
rect 244322 154046 244378 154102
rect 244198 153922 244254 153978
rect 244322 153922 244378 153978
rect 44518 148294 44574 148350
rect 44642 148294 44698 148350
rect 44518 148170 44574 148226
rect 44642 148170 44698 148226
rect 44518 148046 44574 148102
rect 44642 148046 44698 148102
rect 44518 147922 44574 147978
rect 44642 147922 44698 147978
rect 75238 148294 75294 148350
rect 75362 148294 75418 148350
rect 75238 148170 75294 148226
rect 75362 148170 75418 148226
rect 75238 148046 75294 148102
rect 75362 148046 75418 148102
rect 75238 147922 75294 147978
rect 75362 147922 75418 147978
rect 105958 148294 106014 148350
rect 106082 148294 106138 148350
rect 105958 148170 106014 148226
rect 106082 148170 106138 148226
rect 105958 148046 106014 148102
rect 106082 148046 106138 148102
rect 105958 147922 106014 147978
rect 106082 147922 106138 147978
rect 136678 148294 136734 148350
rect 136802 148294 136858 148350
rect 136678 148170 136734 148226
rect 136802 148170 136858 148226
rect 136678 148046 136734 148102
rect 136802 148046 136858 148102
rect 136678 147922 136734 147978
rect 136802 147922 136858 147978
rect 167398 148294 167454 148350
rect 167522 148294 167578 148350
rect 167398 148170 167454 148226
rect 167522 148170 167578 148226
rect 167398 148046 167454 148102
rect 167522 148046 167578 148102
rect 167398 147922 167454 147978
rect 167522 147922 167578 147978
rect 198118 148294 198174 148350
rect 198242 148294 198298 148350
rect 198118 148170 198174 148226
rect 198242 148170 198298 148226
rect 198118 148046 198174 148102
rect 198242 148046 198298 148102
rect 198118 147922 198174 147978
rect 198242 147922 198298 147978
rect 228838 148294 228894 148350
rect 228962 148294 229018 148350
rect 228838 148170 228894 148226
rect 228962 148170 229018 148226
rect 228838 148046 228894 148102
rect 228962 148046 229018 148102
rect 228838 147922 228894 147978
rect 228962 147922 229018 147978
rect 259558 148294 259614 148350
rect 259682 148294 259738 148350
rect 259558 148170 259614 148226
rect 259682 148170 259738 148226
rect 259558 148046 259614 148102
rect 259682 148046 259738 148102
rect 259558 147922 259614 147978
rect 259682 147922 259738 147978
rect 59878 136294 59934 136350
rect 60002 136294 60058 136350
rect 59878 136170 59934 136226
rect 60002 136170 60058 136226
rect 59878 136046 59934 136102
rect 60002 136046 60058 136102
rect 59878 135922 59934 135978
rect 60002 135922 60058 135978
rect 90598 136294 90654 136350
rect 90722 136294 90778 136350
rect 90598 136170 90654 136226
rect 90722 136170 90778 136226
rect 90598 136046 90654 136102
rect 90722 136046 90778 136102
rect 90598 135922 90654 135978
rect 90722 135922 90778 135978
rect 121318 136294 121374 136350
rect 121442 136294 121498 136350
rect 121318 136170 121374 136226
rect 121442 136170 121498 136226
rect 121318 136046 121374 136102
rect 121442 136046 121498 136102
rect 121318 135922 121374 135978
rect 121442 135922 121498 135978
rect 152038 136294 152094 136350
rect 152162 136294 152218 136350
rect 152038 136170 152094 136226
rect 152162 136170 152218 136226
rect 152038 136046 152094 136102
rect 152162 136046 152218 136102
rect 152038 135922 152094 135978
rect 152162 135922 152218 135978
rect 182758 136294 182814 136350
rect 182882 136294 182938 136350
rect 182758 136170 182814 136226
rect 182882 136170 182938 136226
rect 182758 136046 182814 136102
rect 182882 136046 182938 136102
rect 182758 135922 182814 135978
rect 182882 135922 182938 135978
rect 213478 136294 213534 136350
rect 213602 136294 213658 136350
rect 213478 136170 213534 136226
rect 213602 136170 213658 136226
rect 213478 136046 213534 136102
rect 213602 136046 213658 136102
rect 213478 135922 213534 135978
rect 213602 135922 213658 135978
rect 244198 136294 244254 136350
rect 244322 136294 244378 136350
rect 244198 136170 244254 136226
rect 244322 136170 244378 136226
rect 244198 136046 244254 136102
rect 244322 136046 244378 136102
rect 244198 135922 244254 135978
rect 244322 135922 244378 135978
rect 44518 130294 44574 130350
rect 44642 130294 44698 130350
rect 44518 130170 44574 130226
rect 44642 130170 44698 130226
rect 44518 130046 44574 130102
rect 44642 130046 44698 130102
rect 44518 129922 44574 129978
rect 44642 129922 44698 129978
rect 75238 130294 75294 130350
rect 75362 130294 75418 130350
rect 75238 130170 75294 130226
rect 75362 130170 75418 130226
rect 75238 130046 75294 130102
rect 75362 130046 75418 130102
rect 75238 129922 75294 129978
rect 75362 129922 75418 129978
rect 105958 130294 106014 130350
rect 106082 130294 106138 130350
rect 105958 130170 106014 130226
rect 106082 130170 106138 130226
rect 105958 130046 106014 130102
rect 106082 130046 106138 130102
rect 105958 129922 106014 129978
rect 106082 129922 106138 129978
rect 136678 130294 136734 130350
rect 136802 130294 136858 130350
rect 136678 130170 136734 130226
rect 136802 130170 136858 130226
rect 136678 130046 136734 130102
rect 136802 130046 136858 130102
rect 136678 129922 136734 129978
rect 136802 129922 136858 129978
rect 167398 130294 167454 130350
rect 167522 130294 167578 130350
rect 167398 130170 167454 130226
rect 167522 130170 167578 130226
rect 167398 130046 167454 130102
rect 167522 130046 167578 130102
rect 167398 129922 167454 129978
rect 167522 129922 167578 129978
rect 198118 130294 198174 130350
rect 198242 130294 198298 130350
rect 198118 130170 198174 130226
rect 198242 130170 198298 130226
rect 198118 130046 198174 130102
rect 198242 130046 198298 130102
rect 198118 129922 198174 129978
rect 198242 129922 198298 129978
rect 228838 130294 228894 130350
rect 228962 130294 229018 130350
rect 228838 130170 228894 130226
rect 228962 130170 229018 130226
rect 228838 130046 228894 130102
rect 228962 130046 229018 130102
rect 228838 129922 228894 129978
rect 228962 129922 229018 129978
rect 259558 130294 259614 130350
rect 259682 130294 259738 130350
rect 259558 130170 259614 130226
rect 259682 130170 259738 130226
rect 259558 130046 259614 130102
rect 259682 130046 259738 130102
rect 259558 129922 259614 129978
rect 259682 129922 259738 129978
rect 59878 118294 59934 118350
rect 60002 118294 60058 118350
rect 59878 118170 59934 118226
rect 60002 118170 60058 118226
rect 59878 118046 59934 118102
rect 60002 118046 60058 118102
rect 59878 117922 59934 117978
rect 60002 117922 60058 117978
rect 90598 118294 90654 118350
rect 90722 118294 90778 118350
rect 90598 118170 90654 118226
rect 90722 118170 90778 118226
rect 90598 118046 90654 118102
rect 90722 118046 90778 118102
rect 90598 117922 90654 117978
rect 90722 117922 90778 117978
rect 121318 118294 121374 118350
rect 121442 118294 121498 118350
rect 121318 118170 121374 118226
rect 121442 118170 121498 118226
rect 121318 118046 121374 118102
rect 121442 118046 121498 118102
rect 121318 117922 121374 117978
rect 121442 117922 121498 117978
rect 152038 118294 152094 118350
rect 152162 118294 152218 118350
rect 152038 118170 152094 118226
rect 152162 118170 152218 118226
rect 152038 118046 152094 118102
rect 152162 118046 152218 118102
rect 152038 117922 152094 117978
rect 152162 117922 152218 117978
rect 182758 118294 182814 118350
rect 182882 118294 182938 118350
rect 182758 118170 182814 118226
rect 182882 118170 182938 118226
rect 182758 118046 182814 118102
rect 182882 118046 182938 118102
rect 182758 117922 182814 117978
rect 182882 117922 182938 117978
rect 213478 118294 213534 118350
rect 213602 118294 213658 118350
rect 213478 118170 213534 118226
rect 213602 118170 213658 118226
rect 213478 118046 213534 118102
rect 213602 118046 213658 118102
rect 213478 117922 213534 117978
rect 213602 117922 213658 117978
rect 244198 118294 244254 118350
rect 244322 118294 244378 118350
rect 244198 118170 244254 118226
rect 244322 118170 244378 118226
rect 244198 118046 244254 118102
rect 244322 118046 244378 118102
rect 244198 117922 244254 117978
rect 244322 117922 244378 117978
rect 44518 112294 44574 112350
rect 44642 112294 44698 112350
rect 44518 112170 44574 112226
rect 44642 112170 44698 112226
rect 44518 112046 44574 112102
rect 44642 112046 44698 112102
rect 44518 111922 44574 111978
rect 44642 111922 44698 111978
rect 75238 112294 75294 112350
rect 75362 112294 75418 112350
rect 75238 112170 75294 112226
rect 75362 112170 75418 112226
rect 75238 112046 75294 112102
rect 75362 112046 75418 112102
rect 75238 111922 75294 111978
rect 75362 111922 75418 111978
rect 105958 112294 106014 112350
rect 106082 112294 106138 112350
rect 105958 112170 106014 112226
rect 106082 112170 106138 112226
rect 105958 112046 106014 112102
rect 106082 112046 106138 112102
rect 105958 111922 106014 111978
rect 106082 111922 106138 111978
rect 136678 112294 136734 112350
rect 136802 112294 136858 112350
rect 136678 112170 136734 112226
rect 136802 112170 136858 112226
rect 136678 112046 136734 112102
rect 136802 112046 136858 112102
rect 136678 111922 136734 111978
rect 136802 111922 136858 111978
rect 167398 112294 167454 112350
rect 167522 112294 167578 112350
rect 167398 112170 167454 112226
rect 167522 112170 167578 112226
rect 167398 112046 167454 112102
rect 167522 112046 167578 112102
rect 167398 111922 167454 111978
rect 167522 111922 167578 111978
rect 198118 112294 198174 112350
rect 198242 112294 198298 112350
rect 198118 112170 198174 112226
rect 198242 112170 198298 112226
rect 198118 112046 198174 112102
rect 198242 112046 198298 112102
rect 198118 111922 198174 111978
rect 198242 111922 198298 111978
rect 228838 112294 228894 112350
rect 228962 112294 229018 112350
rect 228838 112170 228894 112226
rect 228962 112170 229018 112226
rect 228838 112046 228894 112102
rect 228962 112046 229018 112102
rect 228838 111922 228894 111978
rect 228962 111922 229018 111978
rect 259558 112294 259614 112350
rect 259682 112294 259738 112350
rect 259558 112170 259614 112226
rect 259682 112170 259738 112226
rect 259558 112046 259614 112102
rect 259682 112046 259738 112102
rect 259558 111922 259614 111978
rect 259682 111922 259738 111978
rect 59878 100294 59934 100350
rect 60002 100294 60058 100350
rect 59878 100170 59934 100226
rect 60002 100170 60058 100226
rect 59878 100046 59934 100102
rect 60002 100046 60058 100102
rect 59878 99922 59934 99978
rect 60002 99922 60058 99978
rect 90598 100294 90654 100350
rect 90722 100294 90778 100350
rect 90598 100170 90654 100226
rect 90722 100170 90778 100226
rect 90598 100046 90654 100102
rect 90722 100046 90778 100102
rect 90598 99922 90654 99978
rect 90722 99922 90778 99978
rect 121318 100294 121374 100350
rect 121442 100294 121498 100350
rect 121318 100170 121374 100226
rect 121442 100170 121498 100226
rect 121318 100046 121374 100102
rect 121442 100046 121498 100102
rect 121318 99922 121374 99978
rect 121442 99922 121498 99978
rect 152038 100294 152094 100350
rect 152162 100294 152218 100350
rect 152038 100170 152094 100226
rect 152162 100170 152218 100226
rect 152038 100046 152094 100102
rect 152162 100046 152218 100102
rect 152038 99922 152094 99978
rect 152162 99922 152218 99978
rect 182758 100294 182814 100350
rect 182882 100294 182938 100350
rect 182758 100170 182814 100226
rect 182882 100170 182938 100226
rect 182758 100046 182814 100102
rect 182882 100046 182938 100102
rect 182758 99922 182814 99978
rect 182882 99922 182938 99978
rect 213478 100294 213534 100350
rect 213602 100294 213658 100350
rect 213478 100170 213534 100226
rect 213602 100170 213658 100226
rect 213478 100046 213534 100102
rect 213602 100046 213658 100102
rect 213478 99922 213534 99978
rect 213602 99922 213658 99978
rect 244198 100294 244254 100350
rect 244322 100294 244378 100350
rect 244198 100170 244254 100226
rect 244322 100170 244378 100226
rect 244198 100046 244254 100102
rect 244322 100046 244378 100102
rect 244198 99922 244254 99978
rect 244322 99922 244378 99978
rect 44518 94294 44574 94350
rect 44642 94294 44698 94350
rect 44518 94170 44574 94226
rect 44642 94170 44698 94226
rect 44518 94046 44574 94102
rect 44642 94046 44698 94102
rect 44518 93922 44574 93978
rect 44642 93922 44698 93978
rect 75238 94294 75294 94350
rect 75362 94294 75418 94350
rect 75238 94170 75294 94226
rect 75362 94170 75418 94226
rect 75238 94046 75294 94102
rect 75362 94046 75418 94102
rect 75238 93922 75294 93978
rect 75362 93922 75418 93978
rect 105958 94294 106014 94350
rect 106082 94294 106138 94350
rect 105958 94170 106014 94226
rect 106082 94170 106138 94226
rect 105958 94046 106014 94102
rect 106082 94046 106138 94102
rect 105958 93922 106014 93978
rect 106082 93922 106138 93978
rect 136678 94294 136734 94350
rect 136802 94294 136858 94350
rect 136678 94170 136734 94226
rect 136802 94170 136858 94226
rect 136678 94046 136734 94102
rect 136802 94046 136858 94102
rect 136678 93922 136734 93978
rect 136802 93922 136858 93978
rect 167398 94294 167454 94350
rect 167522 94294 167578 94350
rect 167398 94170 167454 94226
rect 167522 94170 167578 94226
rect 167398 94046 167454 94102
rect 167522 94046 167578 94102
rect 167398 93922 167454 93978
rect 167522 93922 167578 93978
rect 198118 94294 198174 94350
rect 198242 94294 198298 94350
rect 198118 94170 198174 94226
rect 198242 94170 198298 94226
rect 198118 94046 198174 94102
rect 198242 94046 198298 94102
rect 198118 93922 198174 93978
rect 198242 93922 198298 93978
rect 228838 94294 228894 94350
rect 228962 94294 229018 94350
rect 228838 94170 228894 94226
rect 228962 94170 229018 94226
rect 228838 94046 228894 94102
rect 228962 94046 229018 94102
rect 228838 93922 228894 93978
rect 228962 93922 229018 93978
rect 259558 94294 259614 94350
rect 259682 94294 259738 94350
rect 259558 94170 259614 94226
rect 259682 94170 259738 94226
rect 259558 94046 259614 94102
rect 259682 94046 259738 94102
rect 259558 93922 259614 93978
rect 259682 93922 259738 93978
rect 59878 82294 59934 82350
rect 60002 82294 60058 82350
rect 59878 82170 59934 82226
rect 60002 82170 60058 82226
rect 59878 82046 59934 82102
rect 60002 82046 60058 82102
rect 59878 81922 59934 81978
rect 60002 81922 60058 81978
rect 90598 82294 90654 82350
rect 90722 82294 90778 82350
rect 90598 82170 90654 82226
rect 90722 82170 90778 82226
rect 90598 82046 90654 82102
rect 90722 82046 90778 82102
rect 90598 81922 90654 81978
rect 90722 81922 90778 81978
rect 121318 82294 121374 82350
rect 121442 82294 121498 82350
rect 121318 82170 121374 82226
rect 121442 82170 121498 82226
rect 121318 82046 121374 82102
rect 121442 82046 121498 82102
rect 121318 81922 121374 81978
rect 121442 81922 121498 81978
rect 152038 82294 152094 82350
rect 152162 82294 152218 82350
rect 152038 82170 152094 82226
rect 152162 82170 152218 82226
rect 152038 82046 152094 82102
rect 152162 82046 152218 82102
rect 152038 81922 152094 81978
rect 152162 81922 152218 81978
rect 182758 82294 182814 82350
rect 182882 82294 182938 82350
rect 182758 82170 182814 82226
rect 182882 82170 182938 82226
rect 182758 82046 182814 82102
rect 182882 82046 182938 82102
rect 182758 81922 182814 81978
rect 182882 81922 182938 81978
rect 213478 82294 213534 82350
rect 213602 82294 213658 82350
rect 213478 82170 213534 82226
rect 213602 82170 213658 82226
rect 213478 82046 213534 82102
rect 213602 82046 213658 82102
rect 213478 81922 213534 81978
rect 213602 81922 213658 81978
rect 244198 82294 244254 82350
rect 244322 82294 244378 82350
rect 244198 82170 244254 82226
rect 244322 82170 244378 82226
rect 244198 82046 244254 82102
rect 244322 82046 244378 82102
rect 244198 81922 244254 81978
rect 244322 81922 244378 81978
rect 44518 76294 44574 76350
rect 44642 76294 44698 76350
rect 44518 76170 44574 76226
rect 44642 76170 44698 76226
rect 44518 76046 44574 76102
rect 44642 76046 44698 76102
rect 44518 75922 44574 75978
rect 44642 75922 44698 75978
rect 75238 76294 75294 76350
rect 75362 76294 75418 76350
rect 75238 76170 75294 76226
rect 75362 76170 75418 76226
rect 75238 76046 75294 76102
rect 75362 76046 75418 76102
rect 75238 75922 75294 75978
rect 75362 75922 75418 75978
rect 105958 76294 106014 76350
rect 106082 76294 106138 76350
rect 105958 76170 106014 76226
rect 106082 76170 106138 76226
rect 105958 76046 106014 76102
rect 106082 76046 106138 76102
rect 105958 75922 106014 75978
rect 106082 75922 106138 75978
rect 136678 76294 136734 76350
rect 136802 76294 136858 76350
rect 136678 76170 136734 76226
rect 136802 76170 136858 76226
rect 136678 76046 136734 76102
rect 136802 76046 136858 76102
rect 136678 75922 136734 75978
rect 136802 75922 136858 75978
rect 167398 76294 167454 76350
rect 167522 76294 167578 76350
rect 167398 76170 167454 76226
rect 167522 76170 167578 76226
rect 167398 76046 167454 76102
rect 167522 76046 167578 76102
rect 167398 75922 167454 75978
rect 167522 75922 167578 75978
rect 198118 76294 198174 76350
rect 198242 76294 198298 76350
rect 198118 76170 198174 76226
rect 198242 76170 198298 76226
rect 198118 76046 198174 76102
rect 198242 76046 198298 76102
rect 198118 75922 198174 75978
rect 198242 75922 198298 75978
rect 228838 76294 228894 76350
rect 228962 76294 229018 76350
rect 228838 76170 228894 76226
rect 228962 76170 229018 76226
rect 228838 76046 228894 76102
rect 228962 76046 229018 76102
rect 228838 75922 228894 75978
rect 228962 75922 229018 75978
rect 259558 76294 259614 76350
rect 259682 76294 259738 76350
rect 259558 76170 259614 76226
rect 259682 76170 259738 76226
rect 259558 76046 259614 76102
rect 259682 76046 259738 76102
rect 259558 75922 259614 75978
rect 259682 75922 259738 75978
rect 59878 64294 59934 64350
rect 60002 64294 60058 64350
rect 59878 64170 59934 64226
rect 60002 64170 60058 64226
rect 59878 64046 59934 64102
rect 60002 64046 60058 64102
rect 59878 63922 59934 63978
rect 60002 63922 60058 63978
rect 90598 64294 90654 64350
rect 90722 64294 90778 64350
rect 90598 64170 90654 64226
rect 90722 64170 90778 64226
rect 90598 64046 90654 64102
rect 90722 64046 90778 64102
rect 90598 63922 90654 63978
rect 90722 63922 90778 63978
rect 121318 64294 121374 64350
rect 121442 64294 121498 64350
rect 121318 64170 121374 64226
rect 121442 64170 121498 64226
rect 121318 64046 121374 64102
rect 121442 64046 121498 64102
rect 121318 63922 121374 63978
rect 121442 63922 121498 63978
rect 152038 64294 152094 64350
rect 152162 64294 152218 64350
rect 152038 64170 152094 64226
rect 152162 64170 152218 64226
rect 152038 64046 152094 64102
rect 152162 64046 152218 64102
rect 152038 63922 152094 63978
rect 152162 63922 152218 63978
rect 182758 64294 182814 64350
rect 182882 64294 182938 64350
rect 182758 64170 182814 64226
rect 182882 64170 182938 64226
rect 182758 64046 182814 64102
rect 182882 64046 182938 64102
rect 182758 63922 182814 63978
rect 182882 63922 182938 63978
rect 213478 64294 213534 64350
rect 213602 64294 213658 64350
rect 213478 64170 213534 64226
rect 213602 64170 213658 64226
rect 213478 64046 213534 64102
rect 213602 64046 213658 64102
rect 213478 63922 213534 63978
rect 213602 63922 213658 63978
rect 244198 64294 244254 64350
rect 244322 64294 244378 64350
rect 244198 64170 244254 64226
rect 244322 64170 244378 64226
rect 244198 64046 244254 64102
rect 244322 64046 244378 64102
rect 244198 63922 244254 63978
rect 244322 63922 244378 63978
rect 44518 58294 44574 58350
rect 44642 58294 44698 58350
rect 44518 58170 44574 58226
rect 44642 58170 44698 58226
rect 44518 58046 44574 58102
rect 44642 58046 44698 58102
rect 44518 57922 44574 57978
rect 44642 57922 44698 57978
rect 75238 58294 75294 58350
rect 75362 58294 75418 58350
rect 75238 58170 75294 58226
rect 75362 58170 75418 58226
rect 75238 58046 75294 58102
rect 75362 58046 75418 58102
rect 75238 57922 75294 57978
rect 75362 57922 75418 57978
rect 105958 58294 106014 58350
rect 106082 58294 106138 58350
rect 105958 58170 106014 58226
rect 106082 58170 106138 58226
rect 105958 58046 106014 58102
rect 106082 58046 106138 58102
rect 105958 57922 106014 57978
rect 106082 57922 106138 57978
rect 136678 58294 136734 58350
rect 136802 58294 136858 58350
rect 136678 58170 136734 58226
rect 136802 58170 136858 58226
rect 136678 58046 136734 58102
rect 136802 58046 136858 58102
rect 136678 57922 136734 57978
rect 136802 57922 136858 57978
rect 167398 58294 167454 58350
rect 167522 58294 167578 58350
rect 167398 58170 167454 58226
rect 167522 58170 167578 58226
rect 167398 58046 167454 58102
rect 167522 58046 167578 58102
rect 167398 57922 167454 57978
rect 167522 57922 167578 57978
rect 198118 58294 198174 58350
rect 198242 58294 198298 58350
rect 198118 58170 198174 58226
rect 198242 58170 198298 58226
rect 198118 58046 198174 58102
rect 198242 58046 198298 58102
rect 198118 57922 198174 57978
rect 198242 57922 198298 57978
rect 228838 58294 228894 58350
rect 228962 58294 229018 58350
rect 228838 58170 228894 58226
rect 228962 58170 229018 58226
rect 228838 58046 228894 58102
rect 228962 58046 229018 58102
rect 228838 57922 228894 57978
rect 228962 57922 229018 57978
rect 259558 58294 259614 58350
rect 259682 58294 259738 58350
rect 259558 58170 259614 58226
rect 259682 58170 259738 58226
rect 259558 58046 259614 58102
rect 259682 58046 259738 58102
rect 259558 57922 259614 57978
rect 259682 57922 259738 57978
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 46294 101450 46350
rect 101518 46294 101574 46350
rect 101642 46294 101698 46350
rect 101766 46294 101822 46350
rect 101394 46170 101450 46226
rect 101518 46170 101574 46226
rect 101642 46170 101698 46226
rect 101766 46170 101822 46226
rect 101394 46046 101450 46102
rect 101518 46046 101574 46102
rect 101642 46046 101698 46102
rect 101766 46046 101822 46102
rect 101394 45922 101450 45978
rect 101518 45922 101574 45978
rect 101642 45922 101698 45978
rect 101766 45922 101822 45978
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 267036 204902 267092 204958
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 267372 236942 267428 236998
rect 267932 205802 267988 205858
rect 267596 204002 267652 204058
rect 268044 201482 268100 201538
rect 267932 143342 267988 143398
rect 268716 115262 268772 115318
rect 268604 115082 268660 115138
rect 269724 206522 269780 206578
rect 269612 201482 269668 201538
rect 269836 204902 269892 204958
rect 270620 55322 270676 55378
rect 271404 222542 271460 222598
rect 271628 206162 271684 206218
rect 271852 205982 271908 206038
rect 272300 204182 272356 204238
rect 272188 143342 272244 143398
rect 272188 142802 272244 142858
rect 273084 207422 273140 207478
rect 272972 206388 273028 206398
rect 272972 206342 273028 206388
rect 272972 143882 273028 143938
rect 273196 143522 273252 143578
rect 274764 212462 274820 212518
rect 274652 211022 274708 211078
rect 273756 143522 273812 143578
rect 274876 204362 274932 204418
rect 274988 161162 275044 161218
rect 274988 132542 275044 132598
rect 276332 211742 276388 211798
rect 276556 160982 276612 161038
rect 276332 35162 276388 35218
rect 278236 139382 278292 139438
rect 286412 239462 286468 239518
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 279692 236042 279748 236098
rect 281484 231002 281540 231058
rect 280140 143702 280196 143758
rect 280252 131822 280308 131878
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281708 159542 281764 159598
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281372 104102 281428 104158
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 283164 215882 283220 215938
rect 282604 132542 282660 132598
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 283164 150362 283220 150418
rect 283052 103922 283108 103978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 281994 76294 282050 76350
rect 282118 76294 282174 76350
rect 282242 76294 282298 76350
rect 282366 76294 282422 76350
rect 281994 76170 282050 76226
rect 282118 76170 282174 76226
rect 282242 76170 282298 76226
rect 282366 76170 282422 76226
rect 281994 76046 282050 76102
rect 282118 76046 282174 76102
rect 282242 76046 282298 76102
rect 282366 76046 282422 76102
rect 281994 75922 282050 75978
rect 282118 75922 282174 75978
rect 282242 75922 282298 75978
rect 282366 75922 282422 75978
rect 281994 58294 282050 58350
rect 282118 58294 282174 58350
rect 282242 58294 282298 58350
rect 282366 58294 282422 58350
rect 281994 58170 282050 58226
rect 282118 58170 282174 58226
rect 282242 58170 282298 58226
rect 282366 58170 282422 58226
rect 281994 58046 282050 58102
rect 282118 58046 282174 58102
rect 282242 58046 282298 58102
rect 282366 58046 282422 58102
rect 281994 57922 282050 57978
rect 282118 57922 282174 57978
rect 282242 57922 282298 57978
rect 282366 57922 282422 57978
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 285180 219122 285236 219178
rect 285292 151982 285348 152038
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285180 134342 285236 134398
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 285714 64294 285770 64350
rect 285838 64294 285894 64350
rect 285962 64294 286018 64350
rect 286086 64294 286142 64350
rect 285714 64170 285770 64226
rect 285838 64170 285894 64226
rect 285962 64170 286018 64226
rect 286086 64170 286142 64226
rect 285714 64046 285770 64102
rect 285838 64046 285894 64102
rect 285962 64046 286018 64102
rect 286086 64046 286142 64102
rect 285714 63922 285770 63978
rect 285838 63922 285894 63978
rect 285962 63922 286018 63978
rect 286086 63922 286142 63978
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 288316 231002 288372 231058
rect 290916 184294 290972 184350
rect 291040 184294 291096 184350
rect 290916 184170 290972 184226
rect 291040 184170 291096 184226
rect 290916 184046 290972 184102
rect 291040 184046 291096 184102
rect 290916 183922 290972 183978
rect 291040 183922 291096 183978
rect 290916 166294 290972 166350
rect 291040 166294 291096 166350
rect 290916 166170 290972 166226
rect 291040 166170 291096 166226
rect 290916 166046 290972 166102
rect 291040 166046 291096 166102
rect 290916 165922 290972 165978
rect 291040 165922 291096 165978
rect 290668 144422 290724 144478
rect 292348 224162 292404 224218
rect 293356 169802 293412 169858
rect 292348 132362 292404 132418
rect 293132 134522 293188 134578
rect 321692 239282 321748 239338
rect 294924 234242 294980 234298
rect 294924 152702 294980 152758
rect 295036 214082 295092 214138
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 295260 170522 295316 170578
rect 298956 198962 299012 199018
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 323372 236222 323428 236278
rect 321692 197342 321748 197398
rect 323148 191402 323204 191458
rect 295578 190294 295634 190350
rect 295702 190294 295758 190350
rect 295578 190170 295634 190226
rect 295702 190170 295758 190226
rect 295578 190046 295634 190102
rect 295702 190046 295758 190102
rect 295578 189922 295634 189978
rect 295702 189922 295758 189978
rect 304902 190294 304958 190350
rect 305026 190294 305082 190350
rect 304902 190170 304958 190226
rect 305026 190170 305082 190226
rect 304902 190046 304958 190102
rect 305026 190046 305082 190102
rect 304902 189922 304958 189978
rect 305026 189922 305082 189978
rect 314226 190294 314282 190350
rect 314350 190294 314406 190350
rect 314226 190170 314282 190226
rect 314350 190170 314406 190226
rect 314226 190046 314282 190102
rect 314350 190046 314406 190102
rect 314226 189922 314282 189978
rect 314350 189922 314406 189978
rect 300240 184294 300296 184350
rect 300364 184294 300420 184350
rect 300240 184170 300296 184226
rect 300364 184170 300420 184226
rect 300240 184046 300296 184102
rect 300364 184046 300420 184102
rect 300240 183922 300296 183978
rect 300364 183922 300420 183978
rect 309564 184294 309620 184350
rect 309688 184294 309744 184350
rect 309564 184170 309620 184226
rect 309688 184170 309744 184226
rect 309564 184046 309620 184102
rect 309688 184046 309744 184102
rect 309564 183922 309620 183978
rect 309688 183922 309744 183978
rect 318888 184294 318944 184350
rect 319012 184294 319068 184350
rect 318888 184170 318944 184226
rect 319012 184170 319068 184226
rect 318888 184046 318944 184102
rect 319012 184046 319068 184102
rect 318888 183922 318944 183978
rect 319012 183922 319068 183978
rect 295578 172294 295634 172350
rect 295702 172294 295758 172350
rect 295578 172170 295634 172226
rect 295702 172170 295758 172226
rect 295578 172046 295634 172102
rect 295702 172046 295758 172102
rect 295578 171922 295634 171978
rect 295702 171922 295758 171978
rect 304902 172294 304958 172350
rect 305026 172294 305082 172350
rect 304902 172170 304958 172226
rect 305026 172170 305082 172226
rect 304902 172046 304958 172102
rect 305026 172046 305082 172102
rect 304902 171922 304958 171978
rect 305026 171922 305082 171978
rect 314226 172294 314282 172350
rect 314350 172294 314406 172350
rect 314226 172170 314282 172226
rect 314350 172170 314406 172226
rect 314226 172046 314282 172102
rect 314350 172046 314406 172102
rect 314226 171922 314282 171978
rect 314350 171922 314406 171978
rect 297500 170522 297556 170578
rect 297388 169802 297444 169858
rect 300240 166294 300296 166350
rect 300364 166294 300420 166350
rect 300240 166170 300296 166226
rect 300364 166170 300420 166226
rect 300240 166046 300296 166102
rect 300364 166046 300420 166102
rect 300240 165922 300296 165978
rect 300364 165922 300420 165978
rect 309564 166294 309620 166350
rect 309688 166294 309744 166350
rect 309564 166170 309620 166226
rect 309688 166170 309744 166226
rect 309564 166046 309620 166102
rect 309688 166046 309744 166102
rect 309564 165922 309620 165978
rect 309688 165922 309744 165978
rect 312714 166294 312770 166350
rect 312838 166294 312894 166350
rect 312962 166294 313018 166350
rect 313086 166294 313142 166350
rect 312714 166170 312770 166226
rect 312838 166170 312894 166226
rect 312962 166170 313018 166226
rect 313086 166170 313142 166226
rect 312714 166046 312770 166102
rect 312838 166046 312894 166102
rect 312962 166046 313018 166102
rect 313086 166046 313142 166102
rect 312714 165922 312770 165978
rect 312838 165922 312894 165978
rect 312962 165922 313018 165978
rect 313086 165922 313142 165978
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 297388 135602 297444 135658
rect 297388 134522 297444 134578
rect 306572 136862 306628 136918
rect 304892 132722 304948 132778
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 299528 82091 299584 82147
rect 299632 82091 299688 82147
rect 299736 82091 299792 82147
rect 299528 81987 299584 82043
rect 299632 81987 299688 82043
rect 299736 81987 299792 82043
rect 299528 81883 299584 81939
rect 299632 81883 299688 81939
rect 299736 81883 299792 81939
rect 307844 82091 307900 82147
rect 307948 82091 308004 82147
rect 308052 82091 308108 82147
rect 307844 81987 307900 82043
rect 307948 81987 308004 82043
rect 308052 81987 308108 82043
rect 307844 81883 307900 81939
rect 307948 81883 308004 81939
rect 308052 81883 308108 81939
rect 318888 166294 318944 166350
rect 319012 166294 319068 166350
rect 318888 166170 318944 166226
rect 319012 166170 319068 166226
rect 318888 166046 318944 166102
rect 319012 166046 319068 166102
rect 318888 165922 318944 165978
rect 319012 165922 319068 165978
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 323550 190294 323606 190350
rect 323674 190294 323730 190350
rect 323550 190170 323606 190226
rect 323674 190170 323730 190226
rect 323550 190046 323606 190102
rect 323674 190046 323730 190102
rect 323550 189922 323606 189978
rect 323674 189922 323730 189978
rect 323550 172294 323606 172350
rect 323674 172294 323730 172350
rect 323550 172170 323606 172226
rect 323674 172170 323730 172226
rect 323550 172046 323606 172102
rect 323674 172046 323730 172102
rect 323550 171922 323606 171978
rect 323674 171922 323730 171978
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 316160 82091 316216 82147
rect 316264 82091 316320 82147
rect 316368 82091 316424 82147
rect 316160 81987 316216 82043
rect 316264 81987 316320 82043
rect 316368 81987 316424 82043
rect 316160 81883 316216 81939
rect 316264 81883 316320 81939
rect 316368 81883 316424 81939
rect 324476 82091 324532 82147
rect 324580 82091 324636 82147
rect 324684 82091 324740 82147
rect 324476 81987 324532 82043
rect 324580 81987 324636 82043
rect 324684 81987 324740 82043
rect 324476 81883 324532 81939
rect 324580 81883 324636 81939
rect 324684 81883 324740 81939
rect 295412 76294 295468 76350
rect 295536 76294 295592 76350
rect 295412 76170 295468 76226
rect 295536 76170 295592 76226
rect 295412 76046 295468 76102
rect 295536 76046 295592 76102
rect 295412 75922 295468 75978
rect 295536 75922 295592 75978
rect 303728 76294 303784 76350
rect 303852 76294 303908 76350
rect 303728 76170 303784 76226
rect 303852 76170 303908 76226
rect 303728 76046 303784 76102
rect 303852 76046 303908 76102
rect 303728 75922 303784 75978
rect 303852 75922 303908 75978
rect 312044 76294 312100 76350
rect 312168 76294 312224 76350
rect 312044 76170 312100 76226
rect 312168 76170 312224 76226
rect 312044 76046 312100 76102
rect 312168 76046 312224 76102
rect 312044 75922 312100 75978
rect 312168 75922 312224 75978
rect 320360 76294 320416 76350
rect 320484 76294 320540 76350
rect 320360 76170 320416 76226
rect 320484 76170 320540 76226
rect 320360 76046 320416 76102
rect 320484 76046 320540 76102
rect 320360 75922 320416 75978
rect 320484 75922 320540 75978
rect 299570 64294 299626 64350
rect 299694 64294 299750 64350
rect 299570 64170 299626 64226
rect 299694 64170 299750 64226
rect 299570 64046 299626 64102
rect 299694 64046 299750 64102
rect 299570 63922 299626 63978
rect 299694 63922 299750 63978
rect 307886 64294 307942 64350
rect 308010 64294 308066 64350
rect 307886 64170 307942 64226
rect 308010 64170 308066 64226
rect 307886 64046 307942 64102
rect 308010 64046 308066 64102
rect 307886 63922 307942 63978
rect 308010 63922 308066 63978
rect 316202 64294 316258 64350
rect 316326 64294 316382 64350
rect 316202 64170 316258 64226
rect 316326 64170 316382 64226
rect 316202 64046 316258 64102
rect 316326 64046 316382 64102
rect 316202 63922 316258 63978
rect 316326 63922 316382 63978
rect 324518 64294 324574 64350
rect 324642 64294 324698 64350
rect 324518 64170 324574 64226
rect 324642 64170 324698 64226
rect 324518 64046 324574 64102
rect 324642 64046 324698 64102
rect 324518 63922 324574 63978
rect 324642 63922 324698 63978
rect 295412 58294 295468 58350
rect 295536 58294 295592 58350
rect 295412 58170 295468 58226
rect 295536 58170 295592 58226
rect 295412 58046 295468 58102
rect 295536 58046 295592 58102
rect 295412 57922 295468 57978
rect 295536 57922 295592 57978
rect 303728 58294 303784 58350
rect 303852 58294 303908 58350
rect 303728 58170 303784 58226
rect 303852 58170 303908 58226
rect 303728 58046 303784 58102
rect 303852 58046 303908 58102
rect 303728 57922 303784 57978
rect 303852 57922 303908 57978
rect 312044 58294 312100 58350
rect 312168 58294 312224 58350
rect 312044 58170 312100 58226
rect 312168 58170 312224 58226
rect 312044 58046 312100 58102
rect 312168 58046 312224 58102
rect 312044 57922 312100 57978
rect 312168 57922 312224 57978
rect 320360 58294 320416 58350
rect 320484 58294 320540 58350
rect 320360 58170 320416 58226
rect 320484 58170 320540 58226
rect 320360 58046 320416 58102
rect 320484 58046 320540 58102
rect 320360 57922 320416 57978
rect 320484 57922 320540 57978
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 325276 210842 325332 210898
rect 325164 157742 325220 157798
rect 326844 240542 326900 240598
rect 326956 240362 327012 240418
rect 326620 162062 326676 162118
rect 327068 238562 327124 238618
rect 326844 198962 326900 199018
rect 327180 155402 327236 155458
rect 327628 239282 327684 239338
rect 326844 140282 326900 140338
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 335132 407402 335188 407458
rect 332780 397322 332836 397378
rect 329084 369602 329140 369658
rect 328524 313262 328580 313318
rect 328636 321002 328692 321058
rect 328412 282662 328468 282718
rect 328524 313082 328580 313138
rect 328412 258542 328468 258598
rect 328300 249182 328356 249238
rect 329308 321002 329364 321058
rect 328860 308222 328916 308278
rect 328748 283742 328804 283798
rect 328860 296522 328916 296578
rect 328636 249542 328692 249598
rect 328748 283022 328804 283078
rect 328748 249362 328804 249418
rect 328636 248282 328692 248338
rect 328748 242162 328804 242218
rect 329308 313124 329364 313138
rect 329308 313082 329364 313124
rect 329084 300842 329140 300898
rect 329084 285722 329140 285778
rect 329308 282662 329364 282718
rect 329084 272942 329140 272998
rect 329420 260342 329476 260398
rect 329196 253682 329252 253738
rect 329084 248462 329140 248518
rect 329196 247922 329252 247978
rect 329084 241982 329140 242038
rect 328972 158642 329028 158698
rect 329980 308222 330036 308278
rect 330204 285722 330260 285778
rect 331548 386522 331604 386578
rect 331772 383642 331828 383698
rect 330428 296522 330484 296578
rect 330540 272942 330596 272998
rect 329756 253682 329812 253738
rect 329756 236222 329812 236278
rect 330428 249542 330484 249598
rect 330988 248462 331044 248518
rect 330876 248102 330932 248158
rect 332668 376442 332724 376498
rect 331772 301562 331828 301618
rect 331212 248282 331268 248338
rect 331100 240362 331156 240418
rect 331660 241982 331716 242038
rect 331548 238588 331604 238618
rect 331548 238562 331604 238588
rect 333004 389942 333060 389998
rect 332892 389762 332948 389818
rect 331996 142622 332052 142678
rect 332332 240722 332388 240778
rect 332220 227582 332276 227638
rect 332332 146942 332388 146998
rect 332444 141902 332500 141958
rect 332668 258542 332724 258598
rect 333228 391562 333284 391618
rect 332892 283742 332948 283798
rect 334572 384722 334628 384778
rect 332668 249182 332724 249238
rect 333116 242162 333172 242218
rect 333340 240542 333396 240598
rect 333564 247922 333620 247978
rect 333004 231002 333060 231058
rect 333452 217502 333508 217558
rect 333340 135242 333396 135298
rect 333900 229202 333956 229258
rect 333788 155582 333844 155638
rect 333900 127502 333956 127558
rect 336028 407222 336084 407278
rect 335916 383516 335972 383518
rect 335916 383462 335972 383516
rect 335356 369602 335412 369658
rect 335132 243422 335188 243478
rect 335020 137582 335076 137638
rect 354620 410462 354676 410518
rect 359996 410462 360052 410518
rect 352828 410102 352884 410158
rect 340844 408842 340900 408898
rect 339612 407222 339668 407278
rect 337484 406682 337540 406738
rect 338492 404702 338548 404758
rect 337708 399662 337764 399718
rect 336028 300842 336084 300898
rect 336140 384902 336196 384958
rect 335580 283922 335636 283978
rect 336252 380042 336308 380098
rect 337708 378062 337764 378118
rect 336364 360782 336420 360838
rect 335692 283022 335748 283078
rect 336252 239462 336308 239518
rect 336028 191436 336084 191458
rect 336028 191402 336084 191436
rect 336028 173042 336084 173098
rect 336028 168002 336084 168058
rect 336140 162242 336196 162298
rect 336140 143882 336196 143938
rect 336924 313262 336980 313318
rect 336812 136862 336868 136918
rect 335916 133982 335972 134038
rect 336028 134162 336084 134218
rect 336812 134162 336868 134218
rect 336028 132722 336084 132778
rect 336812 132182 336868 132238
rect 337036 197342 337092 197398
rect 337148 143882 337204 143938
rect 338716 402902 338772 402958
rect 339500 404162 339556 404218
rect 339052 402542 339108 402598
rect 338716 392282 338772 392338
rect 340172 404882 340228 404938
rect 354508 408122 354564 408178
rect 340956 403262 341012 403318
rect 341516 403442 341572 403498
rect 346108 404342 346164 404398
rect 352156 406700 352212 406738
rect 352156 406682 352212 406700
rect 354732 409922 354788 409978
rect 359772 410102 359828 410158
rect 359660 409922 359716 409978
rect 359548 409562 359604 409618
rect 356188 408842 356244 408898
rect 356636 408482 356692 408538
rect 347900 403442 347956 403498
rect 350476 402902 350532 402958
rect 350700 402902 350756 402958
rect 350924 403082 350980 403138
rect 354508 404342 354564 404398
rect 350812 402722 350868 402778
rect 357308 404882 357364 404938
rect 352716 401462 352772 401518
rect 365932 410462 365988 410518
rect 358540 401462 358596 401518
rect 366268 410102 366324 410158
rect 371308 410102 371364 410158
rect 369628 409922 369684 409978
rect 366156 408662 366212 408718
rect 386204 410102 386260 410158
rect 386092 409922 386148 409978
rect 404908 410102 404964 410158
rect 366044 404702 366100 404758
rect 366156 403982 366212 404038
rect 365932 403802 365988 403858
rect 364812 403082 364868 403138
rect 366156 402902 366212 402958
rect 367948 402722 368004 402778
rect 361228 401462 361284 401518
rect 383068 405602 383124 405658
rect 383068 403262 383124 403318
rect 497034 562294 497090 562350
rect 497158 562294 497214 562350
rect 497282 562294 497338 562350
rect 497406 562294 497462 562350
rect 497034 562170 497090 562226
rect 497158 562170 497214 562226
rect 497282 562170 497338 562226
rect 497406 562170 497462 562226
rect 497034 562046 497090 562102
rect 497158 562046 497214 562102
rect 497282 562046 497338 562102
rect 497406 562046 497462 562102
rect 497034 561922 497090 561978
rect 497158 561922 497214 561978
rect 497282 561922 497338 561978
rect 497406 561922 497462 561978
rect 486358 550294 486414 550350
rect 486482 550294 486538 550350
rect 486358 550170 486414 550226
rect 486482 550170 486538 550226
rect 486358 550046 486414 550102
rect 486482 550046 486538 550102
rect 486358 549922 486414 549978
rect 486482 549922 486538 549978
rect 497034 544294 497090 544350
rect 497158 544294 497214 544350
rect 497282 544294 497338 544350
rect 497406 544294 497462 544350
rect 497034 544170 497090 544226
rect 497158 544170 497214 544226
rect 497282 544170 497338 544226
rect 497406 544170 497462 544226
rect 497034 544046 497090 544102
rect 497158 544046 497214 544102
rect 497282 544046 497338 544102
rect 497406 544046 497462 544102
rect 497034 543922 497090 543978
rect 497158 543922 497214 543978
rect 497282 543922 497338 543978
rect 497406 543922 497462 543978
rect 486358 532294 486414 532350
rect 486482 532294 486538 532350
rect 486358 532170 486414 532226
rect 486482 532170 486538 532226
rect 486358 532046 486414 532102
rect 486482 532046 486538 532102
rect 486358 531922 486414 531978
rect 486482 531922 486538 531978
rect 497034 526294 497090 526350
rect 497158 526294 497214 526350
rect 497282 526294 497338 526350
rect 497406 526294 497462 526350
rect 497034 526170 497090 526226
rect 497158 526170 497214 526226
rect 497282 526170 497338 526226
rect 497406 526170 497462 526226
rect 497034 526046 497090 526102
rect 497158 526046 497214 526102
rect 497282 526046 497338 526102
rect 497406 526046 497462 526102
rect 497034 525922 497090 525978
rect 497158 525922 497214 525978
rect 497282 525922 497338 525978
rect 497406 525922 497462 525978
rect 486358 514294 486414 514350
rect 486482 514294 486538 514350
rect 486358 514170 486414 514226
rect 486482 514170 486538 514226
rect 486358 514046 486414 514102
rect 486482 514046 486538 514102
rect 486358 513922 486414 513978
rect 486482 513922 486538 513978
rect 497034 508294 497090 508350
rect 497158 508294 497214 508350
rect 497282 508294 497338 508350
rect 497406 508294 497462 508350
rect 497034 508170 497090 508226
rect 497158 508170 497214 508226
rect 497282 508170 497338 508226
rect 497406 508170 497462 508226
rect 497034 508046 497090 508102
rect 497158 508046 497214 508102
rect 497282 508046 497338 508102
rect 497406 508046 497462 508102
rect 497034 507922 497090 507978
rect 497158 507922 497214 507978
rect 497282 507922 497338 507978
rect 497406 507922 497462 507978
rect 486358 496294 486414 496350
rect 486482 496294 486538 496350
rect 486358 496170 486414 496226
rect 486482 496170 486538 496226
rect 486358 496046 486414 496102
rect 486482 496046 486538 496102
rect 486358 495922 486414 495978
rect 486482 495922 486538 495978
rect 497034 490294 497090 490350
rect 497158 490294 497214 490350
rect 497282 490294 497338 490350
rect 497406 490294 497462 490350
rect 497034 490170 497090 490226
rect 497158 490170 497214 490226
rect 497282 490170 497338 490226
rect 497406 490170 497462 490226
rect 497034 490046 497090 490102
rect 497158 490046 497214 490102
rect 497282 490046 497338 490102
rect 497406 490046 497462 490102
rect 497034 489922 497090 489978
rect 497158 489922 497214 489978
rect 497282 489922 497338 489978
rect 497406 489922 497462 489978
rect 486358 478294 486414 478350
rect 486482 478294 486538 478350
rect 486358 478170 486414 478226
rect 486482 478170 486538 478226
rect 486358 478046 486414 478102
rect 486482 478046 486538 478102
rect 486358 477922 486414 477978
rect 486482 477922 486538 477978
rect 497034 472294 497090 472350
rect 497158 472294 497214 472350
rect 497282 472294 497338 472350
rect 497406 472294 497462 472350
rect 497034 472170 497090 472226
rect 497158 472170 497214 472226
rect 497282 472170 497338 472226
rect 497406 472170 497462 472226
rect 497034 472046 497090 472102
rect 497158 472046 497214 472102
rect 497282 472046 497338 472102
rect 497406 472046 497462 472102
rect 497034 471922 497090 471978
rect 497158 471922 497214 471978
rect 497282 471922 497338 471978
rect 497406 471922 497462 471978
rect 486358 460294 486414 460350
rect 486482 460294 486538 460350
rect 486358 460170 486414 460226
rect 486482 460170 486538 460226
rect 486358 460046 486414 460102
rect 486482 460046 486538 460102
rect 486358 459922 486414 459978
rect 486482 459922 486538 459978
rect 497034 454294 497090 454350
rect 497158 454294 497214 454350
rect 497282 454294 497338 454350
rect 497406 454294 497462 454350
rect 497034 454170 497090 454226
rect 497158 454170 497214 454226
rect 497282 454170 497338 454226
rect 497406 454170 497462 454226
rect 497034 454046 497090 454102
rect 497158 454046 497214 454102
rect 497282 454046 497338 454102
rect 497406 454046 497462 454102
rect 497034 453922 497090 453978
rect 497158 453922 497214 453978
rect 497282 453922 497338 453978
rect 497406 453922 497462 453978
rect 486358 442294 486414 442350
rect 486482 442294 486538 442350
rect 486358 442170 486414 442226
rect 486482 442170 486538 442226
rect 486358 442046 486414 442102
rect 486482 442046 486538 442102
rect 486358 441922 486414 441978
rect 486482 441922 486538 441978
rect 497034 436294 497090 436350
rect 497158 436294 497214 436350
rect 497282 436294 497338 436350
rect 497406 436294 497462 436350
rect 497034 436170 497090 436226
rect 497158 436170 497214 436226
rect 497282 436170 497338 436226
rect 497406 436170 497462 436226
rect 497034 436046 497090 436102
rect 497158 436046 497214 436102
rect 497282 436046 497338 436102
rect 497406 436046 497462 436102
rect 497034 435922 497090 435978
rect 497158 435922 497214 435978
rect 497282 435922 497338 435978
rect 497406 435922 497462 435978
rect 486358 424294 486414 424350
rect 486482 424294 486538 424350
rect 486358 424170 486414 424226
rect 486482 424170 486538 424226
rect 486358 424046 486414 424102
rect 486482 424046 486538 424102
rect 486358 423922 486414 423978
rect 486482 423922 486538 423978
rect 497034 418294 497090 418350
rect 497158 418294 497214 418350
rect 497282 418294 497338 418350
rect 497406 418294 497462 418350
rect 497034 418170 497090 418226
rect 497158 418170 497214 418226
rect 497282 418170 497338 418226
rect 497406 418170 497462 418226
rect 497034 418046 497090 418102
rect 497158 418046 497214 418102
rect 497282 418046 497338 418102
rect 497406 418046 497462 418102
rect 497034 417922 497090 417978
rect 497158 417922 497214 417978
rect 497282 417922 497338 417978
rect 497406 417922 497462 417978
rect 496412 408482 496468 408538
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 500754 568294 500810 568350
rect 500878 568294 500934 568350
rect 501002 568294 501058 568350
rect 501126 568294 501182 568350
rect 500754 568170 500810 568226
rect 500878 568170 500934 568226
rect 501002 568170 501058 568226
rect 501126 568170 501182 568226
rect 500754 568046 500810 568102
rect 500878 568046 500934 568102
rect 501002 568046 501058 568102
rect 501126 568046 501182 568102
rect 500754 567922 500810 567978
rect 500878 567922 500934 567978
rect 501002 567922 501058 567978
rect 501126 567922 501182 567978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 501718 562294 501774 562350
rect 501842 562294 501898 562350
rect 501718 562170 501774 562226
rect 501842 562170 501898 562226
rect 501718 562046 501774 562102
rect 501842 562046 501898 562102
rect 501718 561922 501774 561978
rect 501842 561922 501898 561978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 527754 562294 527810 562350
rect 527878 562294 527934 562350
rect 528002 562294 528058 562350
rect 528126 562294 528182 562350
rect 527754 562170 527810 562226
rect 527878 562170 527934 562226
rect 528002 562170 528058 562226
rect 528126 562170 528182 562226
rect 527754 562046 527810 562102
rect 527878 562046 527934 562102
rect 528002 562046 528058 562102
rect 528126 562046 528182 562102
rect 527754 561922 527810 561978
rect 527878 561922 527934 561978
rect 528002 561922 528058 561978
rect 528126 561922 528182 561978
rect 500754 550294 500810 550350
rect 500878 550294 500934 550350
rect 501002 550294 501058 550350
rect 501126 550294 501182 550350
rect 500754 550170 500810 550226
rect 500878 550170 500934 550226
rect 501002 550170 501058 550226
rect 501126 550170 501182 550226
rect 500754 550046 500810 550102
rect 500878 550046 500934 550102
rect 501002 550046 501058 550102
rect 501126 550046 501182 550102
rect 500754 549922 500810 549978
rect 500878 549922 500934 549978
rect 501002 549922 501058 549978
rect 501126 549922 501182 549978
rect 517078 550294 517134 550350
rect 517202 550294 517258 550350
rect 517078 550170 517134 550226
rect 517202 550170 517258 550226
rect 517078 550046 517134 550102
rect 517202 550046 517258 550102
rect 517078 549922 517134 549978
rect 517202 549922 517258 549978
rect 501718 544294 501774 544350
rect 501842 544294 501898 544350
rect 501718 544170 501774 544226
rect 501842 544170 501898 544226
rect 501718 544046 501774 544102
rect 501842 544046 501898 544102
rect 501718 543922 501774 543978
rect 501842 543922 501898 543978
rect 527754 544294 527810 544350
rect 527878 544294 527934 544350
rect 528002 544294 528058 544350
rect 528126 544294 528182 544350
rect 527754 544170 527810 544226
rect 527878 544170 527934 544226
rect 528002 544170 528058 544226
rect 528126 544170 528182 544226
rect 527754 544046 527810 544102
rect 527878 544046 527934 544102
rect 528002 544046 528058 544102
rect 528126 544046 528182 544102
rect 527754 543922 527810 543978
rect 527878 543922 527934 543978
rect 528002 543922 528058 543978
rect 528126 543922 528182 543978
rect 500754 532294 500810 532350
rect 500878 532294 500934 532350
rect 501002 532294 501058 532350
rect 501126 532294 501182 532350
rect 500754 532170 500810 532226
rect 500878 532170 500934 532226
rect 501002 532170 501058 532226
rect 501126 532170 501182 532226
rect 500754 532046 500810 532102
rect 500878 532046 500934 532102
rect 501002 532046 501058 532102
rect 501126 532046 501182 532102
rect 500754 531922 500810 531978
rect 500878 531922 500934 531978
rect 501002 531922 501058 531978
rect 501126 531922 501182 531978
rect 517078 532294 517134 532350
rect 517202 532294 517258 532350
rect 517078 532170 517134 532226
rect 517202 532170 517258 532226
rect 517078 532046 517134 532102
rect 517202 532046 517258 532102
rect 517078 531922 517134 531978
rect 517202 531922 517258 531978
rect 501718 526294 501774 526350
rect 501842 526294 501898 526350
rect 501718 526170 501774 526226
rect 501842 526170 501898 526226
rect 501718 526046 501774 526102
rect 501842 526046 501898 526102
rect 501718 525922 501774 525978
rect 501842 525922 501898 525978
rect 527754 526294 527810 526350
rect 527878 526294 527934 526350
rect 528002 526294 528058 526350
rect 528126 526294 528182 526350
rect 527754 526170 527810 526226
rect 527878 526170 527934 526226
rect 528002 526170 528058 526226
rect 528126 526170 528182 526226
rect 527754 526046 527810 526102
rect 527878 526046 527934 526102
rect 528002 526046 528058 526102
rect 528126 526046 528182 526102
rect 527754 525922 527810 525978
rect 527878 525922 527934 525978
rect 528002 525922 528058 525978
rect 528126 525922 528182 525978
rect 500754 514294 500810 514350
rect 500878 514294 500934 514350
rect 501002 514294 501058 514350
rect 501126 514294 501182 514350
rect 500754 514170 500810 514226
rect 500878 514170 500934 514226
rect 501002 514170 501058 514226
rect 501126 514170 501182 514226
rect 500754 514046 500810 514102
rect 500878 514046 500934 514102
rect 501002 514046 501058 514102
rect 501126 514046 501182 514102
rect 500754 513922 500810 513978
rect 500878 513922 500934 513978
rect 501002 513922 501058 513978
rect 501126 513922 501182 513978
rect 517078 514294 517134 514350
rect 517202 514294 517258 514350
rect 517078 514170 517134 514226
rect 517202 514170 517258 514226
rect 517078 514046 517134 514102
rect 517202 514046 517258 514102
rect 517078 513922 517134 513978
rect 517202 513922 517258 513978
rect 501718 508294 501774 508350
rect 501842 508294 501898 508350
rect 501718 508170 501774 508226
rect 501842 508170 501898 508226
rect 501718 508046 501774 508102
rect 501842 508046 501898 508102
rect 501718 507922 501774 507978
rect 501842 507922 501898 507978
rect 527754 508294 527810 508350
rect 527878 508294 527934 508350
rect 528002 508294 528058 508350
rect 528126 508294 528182 508350
rect 527754 508170 527810 508226
rect 527878 508170 527934 508226
rect 528002 508170 528058 508226
rect 528126 508170 528182 508226
rect 527754 508046 527810 508102
rect 527878 508046 527934 508102
rect 528002 508046 528058 508102
rect 528126 508046 528182 508102
rect 527754 507922 527810 507978
rect 527878 507922 527934 507978
rect 528002 507922 528058 507978
rect 528126 507922 528182 507978
rect 500754 496294 500810 496350
rect 500878 496294 500934 496350
rect 501002 496294 501058 496350
rect 501126 496294 501182 496350
rect 500754 496170 500810 496226
rect 500878 496170 500934 496226
rect 501002 496170 501058 496226
rect 501126 496170 501182 496226
rect 500754 496046 500810 496102
rect 500878 496046 500934 496102
rect 501002 496046 501058 496102
rect 501126 496046 501182 496102
rect 500754 495922 500810 495978
rect 500878 495922 500934 495978
rect 501002 495922 501058 495978
rect 501126 495922 501182 495978
rect 517078 496294 517134 496350
rect 517202 496294 517258 496350
rect 517078 496170 517134 496226
rect 517202 496170 517258 496226
rect 517078 496046 517134 496102
rect 517202 496046 517258 496102
rect 517078 495922 517134 495978
rect 517202 495922 517258 495978
rect 501718 490294 501774 490350
rect 501842 490294 501898 490350
rect 501718 490170 501774 490226
rect 501842 490170 501898 490226
rect 501718 490046 501774 490102
rect 501842 490046 501898 490102
rect 501718 489922 501774 489978
rect 501842 489922 501898 489978
rect 527754 490294 527810 490350
rect 527878 490294 527934 490350
rect 528002 490294 528058 490350
rect 528126 490294 528182 490350
rect 527754 490170 527810 490226
rect 527878 490170 527934 490226
rect 528002 490170 528058 490226
rect 528126 490170 528182 490226
rect 527754 490046 527810 490102
rect 527878 490046 527934 490102
rect 528002 490046 528058 490102
rect 528126 490046 528182 490102
rect 527754 489922 527810 489978
rect 527878 489922 527934 489978
rect 528002 489922 528058 489978
rect 528126 489922 528182 489978
rect 500754 478294 500810 478350
rect 500878 478294 500934 478350
rect 501002 478294 501058 478350
rect 501126 478294 501182 478350
rect 500754 478170 500810 478226
rect 500878 478170 500934 478226
rect 501002 478170 501058 478226
rect 501126 478170 501182 478226
rect 500754 478046 500810 478102
rect 500878 478046 500934 478102
rect 501002 478046 501058 478102
rect 501126 478046 501182 478102
rect 500754 477922 500810 477978
rect 500878 477922 500934 477978
rect 501002 477922 501058 477978
rect 501126 477922 501182 477978
rect 517078 478294 517134 478350
rect 517202 478294 517258 478350
rect 517078 478170 517134 478226
rect 517202 478170 517258 478226
rect 517078 478046 517134 478102
rect 517202 478046 517258 478102
rect 517078 477922 517134 477978
rect 517202 477922 517258 477978
rect 501718 472294 501774 472350
rect 501842 472294 501898 472350
rect 501718 472170 501774 472226
rect 501842 472170 501898 472226
rect 501718 472046 501774 472102
rect 501842 472046 501898 472102
rect 501718 471922 501774 471978
rect 501842 471922 501898 471978
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 531474 568294 531530 568350
rect 531598 568294 531654 568350
rect 531722 568294 531778 568350
rect 531846 568294 531902 568350
rect 531474 568170 531530 568226
rect 531598 568170 531654 568226
rect 531722 568170 531778 568226
rect 531846 568170 531902 568226
rect 531474 568046 531530 568102
rect 531598 568046 531654 568102
rect 531722 568046 531778 568102
rect 531846 568046 531902 568102
rect 531474 567922 531530 567978
rect 531598 567922 531654 567978
rect 531722 567922 531778 567978
rect 531846 567922 531902 567978
rect 531474 550294 531530 550350
rect 531598 550294 531654 550350
rect 531722 550294 531778 550350
rect 531846 550294 531902 550350
rect 531474 550170 531530 550226
rect 531598 550170 531654 550226
rect 531722 550170 531778 550226
rect 531846 550170 531902 550226
rect 531474 550046 531530 550102
rect 531598 550046 531654 550102
rect 531722 550046 531778 550102
rect 531846 550046 531902 550102
rect 531474 549922 531530 549978
rect 531598 549922 531654 549978
rect 531722 549922 531778 549978
rect 531846 549922 531902 549978
rect 533148 566162 533204 566218
rect 531474 532294 531530 532350
rect 531598 532294 531654 532350
rect 531722 532294 531778 532350
rect 531846 532294 531902 532350
rect 531474 532170 531530 532226
rect 531598 532170 531654 532226
rect 531722 532170 531778 532226
rect 531846 532170 531902 532226
rect 531474 532046 531530 532102
rect 531598 532046 531654 532102
rect 531722 532046 531778 532102
rect 531846 532046 531902 532102
rect 531474 531922 531530 531978
rect 531598 531922 531654 531978
rect 531722 531922 531778 531978
rect 531846 531922 531902 531978
rect 531474 514294 531530 514350
rect 531598 514294 531654 514350
rect 531722 514294 531778 514350
rect 531846 514294 531902 514350
rect 531474 514170 531530 514226
rect 531598 514170 531654 514226
rect 531722 514170 531778 514226
rect 531846 514170 531902 514226
rect 531474 514046 531530 514102
rect 531598 514046 531654 514102
rect 531722 514046 531778 514102
rect 531846 514046 531902 514102
rect 531474 513922 531530 513978
rect 531598 513922 531654 513978
rect 531722 513922 531778 513978
rect 531846 513922 531902 513978
rect 531474 496294 531530 496350
rect 531598 496294 531654 496350
rect 531722 496294 531778 496350
rect 531846 496294 531902 496350
rect 531474 496170 531530 496226
rect 531598 496170 531654 496226
rect 531722 496170 531778 496226
rect 531846 496170 531902 496226
rect 531474 496046 531530 496102
rect 531598 496046 531654 496102
rect 531722 496046 531778 496102
rect 531846 496046 531902 496102
rect 531474 495922 531530 495978
rect 531598 495922 531654 495978
rect 531722 495922 531778 495978
rect 531846 495922 531902 495978
rect 527754 472294 527810 472350
rect 527878 472294 527934 472350
rect 528002 472294 528058 472350
rect 528126 472294 528182 472350
rect 527754 472170 527810 472226
rect 527878 472170 527934 472226
rect 528002 472170 528058 472226
rect 528126 472170 528182 472226
rect 527754 472046 527810 472102
rect 527878 472046 527934 472102
rect 528002 472046 528058 472102
rect 528126 472046 528182 472102
rect 527754 471922 527810 471978
rect 527878 471922 527934 471978
rect 528002 471922 528058 471978
rect 528126 471922 528182 471978
rect 500754 460294 500810 460350
rect 500878 460294 500934 460350
rect 501002 460294 501058 460350
rect 501126 460294 501182 460350
rect 500754 460170 500810 460226
rect 500878 460170 500934 460226
rect 501002 460170 501058 460226
rect 501126 460170 501182 460226
rect 500754 460046 500810 460102
rect 500878 460046 500934 460102
rect 501002 460046 501058 460102
rect 501126 460046 501182 460102
rect 500754 459922 500810 459978
rect 500878 459922 500934 459978
rect 501002 459922 501058 459978
rect 501126 459922 501182 459978
rect 517078 460294 517134 460350
rect 517202 460294 517258 460350
rect 517078 460170 517134 460226
rect 517202 460170 517258 460226
rect 517078 460046 517134 460102
rect 517202 460046 517258 460102
rect 517078 459922 517134 459978
rect 517202 459922 517258 459978
rect 501718 454294 501774 454350
rect 501842 454294 501898 454350
rect 501718 454170 501774 454226
rect 501842 454170 501898 454226
rect 501718 454046 501774 454102
rect 501842 454046 501898 454102
rect 501718 453922 501774 453978
rect 501842 453922 501898 453978
rect 527754 454294 527810 454350
rect 527878 454294 527934 454350
rect 528002 454294 528058 454350
rect 528126 454294 528182 454350
rect 527754 454170 527810 454226
rect 527878 454170 527934 454226
rect 528002 454170 528058 454226
rect 528126 454170 528182 454226
rect 527754 454046 527810 454102
rect 527878 454046 527934 454102
rect 528002 454046 528058 454102
rect 528126 454046 528182 454102
rect 527754 453922 527810 453978
rect 527878 453922 527934 453978
rect 528002 453922 528058 453978
rect 528126 453922 528182 453978
rect 500754 442294 500810 442350
rect 500878 442294 500934 442350
rect 501002 442294 501058 442350
rect 501126 442294 501182 442350
rect 500754 442170 500810 442226
rect 500878 442170 500934 442226
rect 501002 442170 501058 442226
rect 501126 442170 501182 442226
rect 500754 442046 500810 442102
rect 500878 442046 500934 442102
rect 501002 442046 501058 442102
rect 501126 442046 501182 442102
rect 500754 441922 500810 441978
rect 500878 441922 500934 441978
rect 501002 441922 501058 441978
rect 501126 441922 501182 441978
rect 517078 442294 517134 442350
rect 517202 442294 517258 442350
rect 517078 442170 517134 442226
rect 517202 442170 517258 442226
rect 517078 442046 517134 442102
rect 517202 442046 517258 442102
rect 517078 441922 517134 441978
rect 517202 441922 517258 441978
rect 501718 436294 501774 436350
rect 501842 436294 501898 436350
rect 501718 436170 501774 436226
rect 501842 436170 501898 436226
rect 501718 436046 501774 436102
rect 501842 436046 501898 436102
rect 501718 435922 501774 435978
rect 501842 435922 501898 435978
rect 527754 436294 527810 436350
rect 527878 436294 527934 436350
rect 528002 436294 528058 436350
rect 528126 436294 528182 436350
rect 527754 436170 527810 436226
rect 527878 436170 527934 436226
rect 528002 436170 528058 436226
rect 528126 436170 528182 436226
rect 527754 436046 527810 436102
rect 527878 436046 527934 436102
rect 528002 436046 528058 436102
rect 528126 436046 528182 436102
rect 527754 435922 527810 435978
rect 527878 435922 527934 435978
rect 528002 435922 528058 435978
rect 528126 435922 528182 435978
rect 500754 424294 500810 424350
rect 500878 424294 500934 424350
rect 501002 424294 501058 424350
rect 501126 424294 501182 424350
rect 500754 424170 500810 424226
rect 500878 424170 500934 424226
rect 501002 424170 501058 424226
rect 501126 424170 501182 424226
rect 500754 424046 500810 424102
rect 500878 424046 500934 424102
rect 501002 424046 501058 424102
rect 501126 424046 501182 424102
rect 500754 423922 500810 423978
rect 500878 423922 500934 423978
rect 501002 423922 501058 423978
rect 501126 423922 501182 423978
rect 499324 410282 499380 410338
rect 517078 424294 517134 424350
rect 517202 424294 517258 424350
rect 517078 424170 517134 424226
rect 517202 424170 517258 424226
rect 517078 424046 517134 424102
rect 517202 424046 517258 424102
rect 517078 423922 517134 423978
rect 517202 423922 517258 423978
rect 501718 418294 501774 418350
rect 501842 418294 501898 418350
rect 501718 418170 501774 418226
rect 501842 418170 501898 418226
rect 501718 418046 501774 418102
rect 501842 418046 501898 418102
rect 501718 417922 501774 417978
rect 501842 417922 501898 417978
rect 527754 418294 527810 418350
rect 527878 418294 527934 418350
rect 528002 418294 528058 418350
rect 528126 418294 528182 418350
rect 527754 418170 527810 418226
rect 527878 418170 527934 418226
rect 528002 418170 528058 418226
rect 528126 418170 528182 418226
rect 527754 418046 527810 418102
rect 527878 418046 527934 418102
rect 528002 418046 528058 418102
rect 528126 418046 528182 418102
rect 527754 417922 527810 417978
rect 527878 417922 527934 417978
rect 528002 417922 528058 417978
rect 528126 417922 528182 417978
rect 514108 408302 514164 408358
rect 500754 406294 500810 406350
rect 500878 406294 500934 406350
rect 501002 406294 501058 406350
rect 501126 406294 501182 406350
rect 500754 406170 500810 406226
rect 500878 406170 500934 406226
rect 501002 406170 501058 406226
rect 501126 406170 501182 406226
rect 500754 406046 500810 406102
rect 500878 406046 500934 406102
rect 501002 406046 501058 406102
rect 501126 406046 501182 406102
rect 500754 405922 500810 405978
rect 500878 405922 500934 405978
rect 501002 405922 501058 405978
rect 501126 405922 501182 405978
rect 511868 402542 511924 402598
rect 522172 404162 522228 404218
rect 517020 402362 517076 402418
rect 531474 478294 531530 478350
rect 531598 478294 531654 478350
rect 531722 478294 531778 478350
rect 531846 478294 531902 478350
rect 531474 478170 531530 478226
rect 531598 478170 531654 478226
rect 531722 478170 531778 478226
rect 531846 478170 531902 478226
rect 531474 478046 531530 478102
rect 531598 478046 531654 478102
rect 531722 478046 531778 478102
rect 531846 478046 531902 478102
rect 531474 477922 531530 477978
rect 531598 477922 531654 477978
rect 531722 477922 531778 477978
rect 531846 477922 531902 477978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 531474 460294 531530 460350
rect 531598 460294 531654 460350
rect 531722 460294 531778 460350
rect 531846 460294 531902 460350
rect 531474 460170 531530 460226
rect 531598 460170 531654 460226
rect 531722 460170 531778 460226
rect 531846 460170 531902 460226
rect 531474 460046 531530 460102
rect 531598 460046 531654 460102
rect 531722 460046 531778 460102
rect 531846 460046 531902 460102
rect 531474 459922 531530 459978
rect 531598 459922 531654 459978
rect 531722 459922 531778 459978
rect 531846 459922 531902 459978
rect 531474 442294 531530 442350
rect 531598 442294 531654 442350
rect 531722 442294 531778 442350
rect 531846 442294 531902 442350
rect 531474 442170 531530 442226
rect 531598 442170 531654 442226
rect 531722 442170 531778 442226
rect 531846 442170 531902 442226
rect 531474 442046 531530 442102
rect 531598 442046 531654 442102
rect 531722 442046 531778 442102
rect 531846 442046 531902 442102
rect 531474 441922 531530 441978
rect 531598 441922 531654 441978
rect 531722 441922 531778 441978
rect 531846 441922 531902 441978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 531474 424294 531530 424350
rect 531598 424294 531654 424350
rect 531722 424294 531778 424350
rect 531846 424294 531902 424350
rect 531474 424170 531530 424226
rect 531598 424170 531654 424226
rect 531722 424170 531778 424226
rect 531846 424170 531902 424226
rect 531474 424046 531530 424102
rect 531598 424046 531654 424102
rect 531722 424046 531778 424102
rect 531846 424046 531902 424102
rect 531474 423922 531530 423978
rect 531598 423922 531654 423978
rect 531722 423922 531778 423978
rect 531846 423922 531902 423978
rect 528892 407222 528948 407278
rect 532588 409022 532644 409078
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 558236 408122 558292 408178
rect 543676 407042 543732 407098
rect 551068 406862 551124 406918
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 590492 573722 590548 573778
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 590604 571202 590660 571258
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 590492 569762 590548 569818
rect 590828 569582 590884 569638
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 580636 407582 580692 407638
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 565852 403082 565908 403138
rect 582092 403982 582148 404038
rect 367836 401462 367892 401518
rect 346108 401102 346164 401158
rect 341516 400562 341572 400618
rect 344518 400294 344574 400350
rect 344642 400294 344698 400350
rect 344518 400170 344574 400226
rect 344642 400170 344698 400226
rect 344518 400046 344574 400102
rect 344642 400046 344698 400102
rect 344518 399922 344574 399978
rect 344642 399922 344698 399978
rect 375238 400294 375294 400350
rect 375362 400294 375418 400350
rect 375238 400170 375294 400226
rect 375362 400170 375418 400226
rect 375238 400046 375294 400102
rect 375362 400046 375418 400102
rect 375238 399922 375294 399978
rect 375362 399922 375418 399978
rect 405958 400294 406014 400350
rect 406082 400294 406138 400350
rect 405958 400170 406014 400226
rect 406082 400170 406138 400226
rect 405958 400046 406014 400102
rect 406082 400046 406138 400102
rect 405958 399922 406014 399978
rect 406082 399922 406138 399978
rect 436678 400294 436734 400350
rect 436802 400294 436858 400350
rect 436678 400170 436734 400226
rect 436802 400170 436858 400226
rect 436678 400046 436734 400102
rect 436802 400046 436858 400102
rect 436678 399922 436734 399978
rect 436802 399922 436858 399978
rect 467398 400294 467454 400350
rect 467522 400294 467578 400350
rect 467398 400170 467454 400226
rect 467522 400170 467578 400226
rect 467398 400046 467454 400102
rect 467522 400046 467578 400102
rect 467398 399922 467454 399978
rect 467522 399922 467578 399978
rect 498118 400294 498174 400350
rect 498242 400294 498298 400350
rect 498118 400170 498174 400226
rect 498242 400170 498298 400226
rect 498118 400046 498174 400102
rect 498242 400046 498298 400102
rect 498118 399922 498174 399978
rect 498242 399922 498298 399978
rect 528838 400294 528894 400350
rect 528962 400294 529018 400350
rect 528838 400170 528894 400226
rect 528962 400170 529018 400226
rect 528838 400046 528894 400102
rect 528962 400046 529018 400102
rect 528838 399922 528894 399978
rect 528962 399922 529018 399978
rect 559558 400294 559614 400350
rect 559682 400294 559738 400350
rect 559558 400170 559614 400226
rect 559682 400170 559738 400226
rect 559558 400046 559614 400102
rect 559682 400046 559738 400102
rect 559558 399922 559614 399978
rect 559682 399922 559738 399978
rect 341180 399662 341236 399718
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 582092 391382 582148 391438
rect 587132 391382 587188 391438
rect 359878 388294 359934 388350
rect 360002 388294 360058 388350
rect 359878 388170 359934 388226
rect 360002 388170 360058 388226
rect 359878 388046 359934 388102
rect 360002 388046 360058 388102
rect 359878 387922 359934 387978
rect 360002 387922 360058 387978
rect 390598 388294 390654 388350
rect 390722 388294 390778 388350
rect 390598 388170 390654 388226
rect 390722 388170 390778 388226
rect 390598 388046 390654 388102
rect 390722 388046 390778 388102
rect 390598 387922 390654 387978
rect 390722 387922 390778 387978
rect 421318 388294 421374 388350
rect 421442 388294 421498 388350
rect 421318 388170 421374 388226
rect 421442 388170 421498 388226
rect 421318 388046 421374 388102
rect 421442 388046 421498 388102
rect 421318 387922 421374 387978
rect 421442 387922 421498 387978
rect 452038 388294 452094 388350
rect 452162 388294 452218 388350
rect 452038 388170 452094 388226
rect 452162 388170 452218 388226
rect 452038 388046 452094 388102
rect 452162 388046 452218 388102
rect 452038 387922 452094 387978
rect 452162 387922 452218 387978
rect 482758 388294 482814 388350
rect 482882 388294 482938 388350
rect 482758 388170 482814 388226
rect 482882 388170 482938 388226
rect 482758 388046 482814 388102
rect 482882 388046 482938 388102
rect 482758 387922 482814 387978
rect 482882 387922 482938 387978
rect 513478 388294 513534 388350
rect 513602 388294 513658 388350
rect 513478 388170 513534 388226
rect 513602 388170 513658 388226
rect 513478 388046 513534 388102
rect 513602 388046 513658 388102
rect 513478 387922 513534 387978
rect 513602 387922 513658 387978
rect 544198 388294 544254 388350
rect 544322 388294 544378 388350
rect 544198 388170 544254 388226
rect 544322 388170 544378 388226
rect 544198 388046 544254 388102
rect 544322 388046 544378 388102
rect 544198 387922 544254 387978
rect 544322 387922 544378 387978
rect 574918 388294 574974 388350
rect 575042 388294 575098 388350
rect 574918 388170 574974 388226
rect 575042 388170 575098 388226
rect 574918 388046 574974 388102
rect 575042 388046 575098 388102
rect 574918 387922 574974 387978
rect 575042 387922 575098 387978
rect 338044 311642 338100 311698
rect 338380 240902 338436 240958
rect 338828 249362 338884 249418
rect 338716 145322 338772 145378
rect 338604 142442 338660 142498
rect 337708 132182 337764 132238
rect 337148 127502 337204 127558
rect 334236 33542 334292 33598
rect 330764 31742 330820 31798
rect 344518 382294 344574 382350
rect 344642 382294 344698 382350
rect 344518 382170 344574 382226
rect 344642 382170 344698 382226
rect 344518 382046 344574 382102
rect 344642 382046 344698 382102
rect 344518 381922 344574 381978
rect 344642 381922 344698 381978
rect 375238 382294 375294 382350
rect 375362 382294 375418 382350
rect 375238 382170 375294 382226
rect 375362 382170 375418 382226
rect 375238 382046 375294 382102
rect 375362 382046 375418 382102
rect 375238 381922 375294 381978
rect 375362 381922 375418 381978
rect 405958 382294 406014 382350
rect 406082 382294 406138 382350
rect 405958 382170 406014 382226
rect 406082 382170 406138 382226
rect 405958 382046 406014 382102
rect 406082 382046 406138 382102
rect 405958 381922 406014 381978
rect 406082 381922 406138 381978
rect 436678 382294 436734 382350
rect 436802 382294 436858 382350
rect 436678 382170 436734 382226
rect 436802 382170 436858 382226
rect 436678 382046 436734 382102
rect 436802 382046 436858 382102
rect 436678 381922 436734 381978
rect 436802 381922 436858 381978
rect 467398 382294 467454 382350
rect 467522 382294 467578 382350
rect 467398 382170 467454 382226
rect 467522 382170 467578 382226
rect 467398 382046 467454 382102
rect 467522 382046 467578 382102
rect 467398 381922 467454 381978
rect 467522 381922 467578 381978
rect 498118 382294 498174 382350
rect 498242 382294 498298 382350
rect 498118 382170 498174 382226
rect 498242 382170 498298 382226
rect 498118 382046 498174 382102
rect 498242 382046 498298 382102
rect 498118 381922 498174 381978
rect 498242 381922 498298 381978
rect 528838 382294 528894 382350
rect 528962 382294 529018 382350
rect 528838 382170 528894 382226
rect 528962 382170 529018 382226
rect 528838 382046 528894 382102
rect 528962 382046 529018 382102
rect 528838 381922 528894 381978
rect 528962 381922 529018 381978
rect 559558 382294 559614 382350
rect 559682 382294 559738 382350
rect 559558 382170 559614 382226
rect 559682 382170 559738 382226
rect 559558 382046 559614 382102
rect 559682 382046 559738 382102
rect 559558 381922 559614 381978
rect 559682 381922 559738 381978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 340060 160802 340116 160858
rect 339276 30122 339332 30178
rect 340396 294542 340452 294598
rect 340396 283742 340452 283798
rect 359878 370294 359934 370350
rect 360002 370294 360058 370350
rect 359878 370170 359934 370226
rect 360002 370170 360058 370226
rect 359878 370046 359934 370102
rect 360002 370046 360058 370102
rect 359878 369922 359934 369978
rect 360002 369922 360058 369978
rect 390598 370294 390654 370350
rect 390722 370294 390778 370350
rect 390598 370170 390654 370226
rect 390722 370170 390778 370226
rect 390598 370046 390654 370102
rect 390722 370046 390778 370102
rect 390598 369922 390654 369978
rect 390722 369922 390778 369978
rect 421318 370294 421374 370350
rect 421442 370294 421498 370350
rect 421318 370170 421374 370226
rect 421442 370170 421498 370226
rect 421318 370046 421374 370102
rect 421442 370046 421498 370102
rect 421318 369922 421374 369978
rect 421442 369922 421498 369978
rect 452038 370294 452094 370350
rect 452162 370294 452218 370350
rect 452038 370170 452094 370226
rect 452162 370170 452218 370226
rect 452038 370046 452094 370102
rect 452162 370046 452218 370102
rect 452038 369922 452094 369978
rect 452162 369922 452218 369978
rect 482758 370294 482814 370350
rect 482882 370294 482938 370350
rect 482758 370170 482814 370226
rect 482882 370170 482938 370226
rect 482758 370046 482814 370102
rect 482882 370046 482938 370102
rect 482758 369922 482814 369978
rect 482882 369922 482938 369978
rect 513478 370294 513534 370350
rect 513602 370294 513658 370350
rect 513478 370170 513534 370226
rect 513602 370170 513658 370226
rect 513478 370046 513534 370102
rect 513602 370046 513658 370102
rect 513478 369922 513534 369978
rect 513602 369922 513658 369978
rect 544198 370294 544254 370350
rect 544322 370294 544378 370350
rect 544198 370170 544254 370226
rect 544322 370170 544378 370226
rect 544198 370046 544254 370102
rect 544322 370046 544378 370102
rect 544198 369922 544254 369978
rect 544322 369922 544378 369978
rect 574918 370294 574974 370350
rect 575042 370294 575098 370350
rect 574918 370170 574974 370226
rect 575042 370170 575098 370226
rect 574918 370046 574974 370102
rect 575042 370046 575098 370102
rect 574918 369922 574974 369978
rect 575042 369922 575098 369978
rect 344518 364294 344574 364350
rect 344642 364294 344698 364350
rect 344518 364170 344574 364226
rect 344642 364170 344698 364226
rect 344518 364046 344574 364102
rect 344642 364046 344698 364102
rect 344518 363922 344574 363978
rect 344642 363922 344698 363978
rect 375238 364294 375294 364350
rect 375362 364294 375418 364350
rect 375238 364170 375294 364226
rect 375362 364170 375418 364226
rect 375238 364046 375294 364102
rect 375362 364046 375418 364102
rect 375238 363922 375294 363978
rect 375362 363922 375418 363978
rect 405958 364294 406014 364350
rect 406082 364294 406138 364350
rect 405958 364170 406014 364226
rect 406082 364170 406138 364226
rect 405958 364046 406014 364102
rect 406082 364046 406138 364102
rect 405958 363922 406014 363978
rect 406082 363922 406138 363978
rect 436678 364294 436734 364350
rect 436802 364294 436858 364350
rect 436678 364170 436734 364226
rect 436802 364170 436858 364226
rect 436678 364046 436734 364102
rect 436802 364046 436858 364102
rect 436678 363922 436734 363978
rect 436802 363922 436858 363978
rect 467398 364294 467454 364350
rect 467522 364294 467578 364350
rect 467398 364170 467454 364226
rect 467522 364170 467578 364226
rect 467398 364046 467454 364102
rect 467522 364046 467578 364102
rect 467398 363922 467454 363978
rect 467522 363922 467578 363978
rect 498118 364294 498174 364350
rect 498242 364294 498298 364350
rect 498118 364170 498174 364226
rect 498242 364170 498298 364226
rect 498118 364046 498174 364102
rect 498242 364046 498298 364102
rect 498118 363922 498174 363978
rect 498242 363922 498298 363978
rect 528838 364294 528894 364350
rect 528962 364294 529018 364350
rect 528838 364170 528894 364226
rect 528962 364170 529018 364226
rect 528838 364046 528894 364102
rect 528962 364046 529018 364102
rect 528838 363922 528894 363978
rect 528962 363922 529018 363978
rect 559558 364294 559614 364350
rect 559682 364294 559738 364350
rect 559558 364170 559614 364226
rect 559682 364170 559738 364226
rect 559558 364046 559614 364102
rect 559682 364046 559738 364102
rect 559558 363922 559614 363978
rect 559682 363922 559738 363978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 340508 157562 340564 157618
rect 359878 352294 359934 352350
rect 360002 352294 360058 352350
rect 359878 352170 359934 352226
rect 360002 352170 360058 352226
rect 359878 352046 359934 352102
rect 360002 352046 360058 352102
rect 359878 351922 359934 351978
rect 360002 351922 360058 351978
rect 390598 352294 390654 352350
rect 390722 352294 390778 352350
rect 390598 352170 390654 352226
rect 390722 352170 390778 352226
rect 390598 352046 390654 352102
rect 390722 352046 390778 352102
rect 390598 351922 390654 351978
rect 390722 351922 390778 351978
rect 421318 352294 421374 352350
rect 421442 352294 421498 352350
rect 421318 352170 421374 352226
rect 421442 352170 421498 352226
rect 421318 352046 421374 352102
rect 421442 352046 421498 352102
rect 421318 351922 421374 351978
rect 421442 351922 421498 351978
rect 452038 352294 452094 352350
rect 452162 352294 452218 352350
rect 452038 352170 452094 352226
rect 452162 352170 452218 352226
rect 452038 352046 452094 352102
rect 452162 352046 452218 352102
rect 452038 351922 452094 351978
rect 452162 351922 452218 351978
rect 482758 352294 482814 352350
rect 482882 352294 482938 352350
rect 482758 352170 482814 352226
rect 482882 352170 482938 352226
rect 482758 352046 482814 352102
rect 482882 352046 482938 352102
rect 482758 351922 482814 351978
rect 482882 351922 482938 351978
rect 513478 352294 513534 352350
rect 513602 352294 513658 352350
rect 513478 352170 513534 352226
rect 513602 352170 513658 352226
rect 513478 352046 513534 352102
rect 513602 352046 513658 352102
rect 513478 351922 513534 351978
rect 513602 351922 513658 351978
rect 544198 352294 544254 352350
rect 544322 352294 544378 352350
rect 544198 352170 544254 352226
rect 544322 352170 544378 352226
rect 544198 352046 544254 352102
rect 544322 352046 544378 352102
rect 544198 351922 544254 351978
rect 544322 351922 544378 351978
rect 574918 352294 574974 352350
rect 575042 352294 575098 352350
rect 574918 352170 574974 352226
rect 575042 352170 575098 352226
rect 574918 352046 574974 352102
rect 575042 352046 575098 352102
rect 574918 351922 574974 351978
rect 575042 351922 575098 351978
rect 344518 346294 344574 346350
rect 344642 346294 344698 346350
rect 344518 346170 344574 346226
rect 344642 346170 344698 346226
rect 344518 346046 344574 346102
rect 344642 346046 344698 346102
rect 344518 345922 344574 345978
rect 344642 345922 344698 345978
rect 375238 346294 375294 346350
rect 375362 346294 375418 346350
rect 375238 346170 375294 346226
rect 375362 346170 375418 346226
rect 375238 346046 375294 346102
rect 375362 346046 375418 346102
rect 375238 345922 375294 345978
rect 375362 345922 375418 345978
rect 405958 346294 406014 346350
rect 406082 346294 406138 346350
rect 405958 346170 406014 346226
rect 406082 346170 406138 346226
rect 405958 346046 406014 346102
rect 406082 346046 406138 346102
rect 405958 345922 406014 345978
rect 406082 345922 406138 345978
rect 436678 346294 436734 346350
rect 436802 346294 436858 346350
rect 436678 346170 436734 346226
rect 436802 346170 436858 346226
rect 436678 346046 436734 346102
rect 436802 346046 436858 346102
rect 436678 345922 436734 345978
rect 436802 345922 436858 345978
rect 467398 346294 467454 346350
rect 467522 346294 467578 346350
rect 467398 346170 467454 346226
rect 467522 346170 467578 346226
rect 467398 346046 467454 346102
rect 467522 346046 467578 346102
rect 467398 345922 467454 345978
rect 467522 345922 467578 345978
rect 498118 346294 498174 346350
rect 498242 346294 498298 346350
rect 498118 346170 498174 346226
rect 498242 346170 498298 346226
rect 498118 346046 498174 346102
rect 498242 346046 498298 346102
rect 498118 345922 498174 345978
rect 498242 345922 498298 345978
rect 528838 346294 528894 346350
rect 528962 346294 529018 346350
rect 528838 346170 528894 346226
rect 528962 346170 529018 346226
rect 528838 346046 528894 346102
rect 528962 346046 529018 346102
rect 528838 345922 528894 345978
rect 528962 345922 529018 345978
rect 559558 346294 559614 346350
rect 559682 346294 559738 346350
rect 559558 346170 559614 346226
rect 559682 346170 559738 346226
rect 559558 346046 559614 346102
rect 559682 346046 559738 346102
rect 559558 345922 559614 345978
rect 559682 345922 559738 345978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 359878 334294 359934 334350
rect 360002 334294 360058 334350
rect 359878 334170 359934 334226
rect 360002 334170 360058 334226
rect 359878 334046 359934 334102
rect 360002 334046 360058 334102
rect 359878 333922 359934 333978
rect 360002 333922 360058 333978
rect 390598 334294 390654 334350
rect 390722 334294 390778 334350
rect 390598 334170 390654 334226
rect 390722 334170 390778 334226
rect 390598 334046 390654 334102
rect 390722 334046 390778 334102
rect 390598 333922 390654 333978
rect 390722 333922 390778 333978
rect 421318 334294 421374 334350
rect 421442 334294 421498 334350
rect 421318 334170 421374 334226
rect 421442 334170 421498 334226
rect 421318 334046 421374 334102
rect 421442 334046 421498 334102
rect 421318 333922 421374 333978
rect 421442 333922 421498 333978
rect 452038 334294 452094 334350
rect 452162 334294 452218 334350
rect 452038 334170 452094 334226
rect 452162 334170 452218 334226
rect 452038 334046 452094 334102
rect 452162 334046 452218 334102
rect 452038 333922 452094 333978
rect 452162 333922 452218 333978
rect 482758 334294 482814 334350
rect 482882 334294 482938 334350
rect 482758 334170 482814 334226
rect 482882 334170 482938 334226
rect 482758 334046 482814 334102
rect 482882 334046 482938 334102
rect 482758 333922 482814 333978
rect 482882 333922 482938 333978
rect 513478 334294 513534 334350
rect 513602 334294 513658 334350
rect 513478 334170 513534 334226
rect 513602 334170 513658 334226
rect 513478 334046 513534 334102
rect 513602 334046 513658 334102
rect 513478 333922 513534 333978
rect 513602 333922 513658 333978
rect 544198 334294 544254 334350
rect 544322 334294 544378 334350
rect 544198 334170 544254 334226
rect 544322 334170 544378 334226
rect 544198 334046 544254 334102
rect 544322 334046 544378 334102
rect 544198 333922 544254 333978
rect 544322 333922 544378 333978
rect 574918 334294 574974 334350
rect 575042 334294 575098 334350
rect 574918 334170 574974 334226
rect 575042 334170 575098 334226
rect 574918 334046 574974 334102
rect 575042 334046 575098 334102
rect 574918 333922 574974 333978
rect 575042 333922 575098 333978
rect 344518 328294 344574 328350
rect 344642 328294 344698 328350
rect 344518 328170 344574 328226
rect 344642 328170 344698 328226
rect 344518 328046 344574 328102
rect 344642 328046 344698 328102
rect 344518 327922 344574 327978
rect 344642 327922 344698 327978
rect 375238 328294 375294 328350
rect 375362 328294 375418 328350
rect 375238 328170 375294 328226
rect 375362 328170 375418 328226
rect 375238 328046 375294 328102
rect 375362 328046 375418 328102
rect 375238 327922 375294 327978
rect 375362 327922 375418 327978
rect 405958 328294 406014 328350
rect 406082 328294 406138 328350
rect 405958 328170 406014 328226
rect 406082 328170 406138 328226
rect 405958 328046 406014 328102
rect 406082 328046 406138 328102
rect 405958 327922 406014 327978
rect 406082 327922 406138 327978
rect 436678 328294 436734 328350
rect 436802 328294 436858 328350
rect 436678 328170 436734 328226
rect 436802 328170 436858 328226
rect 436678 328046 436734 328102
rect 436802 328046 436858 328102
rect 436678 327922 436734 327978
rect 436802 327922 436858 327978
rect 467398 328294 467454 328350
rect 467522 328294 467578 328350
rect 467398 328170 467454 328226
rect 467522 328170 467578 328226
rect 467398 328046 467454 328102
rect 467522 328046 467578 328102
rect 467398 327922 467454 327978
rect 467522 327922 467578 327978
rect 498118 328294 498174 328350
rect 498242 328294 498298 328350
rect 498118 328170 498174 328226
rect 498242 328170 498298 328226
rect 498118 328046 498174 328102
rect 498242 328046 498298 328102
rect 498118 327922 498174 327978
rect 498242 327922 498298 327978
rect 528838 328294 528894 328350
rect 528962 328294 529018 328350
rect 528838 328170 528894 328226
rect 528962 328170 529018 328226
rect 528838 328046 528894 328102
rect 528962 328046 529018 328102
rect 528838 327922 528894 327978
rect 528962 327922 529018 327978
rect 559558 328294 559614 328350
rect 559682 328294 559738 328350
rect 559558 328170 559614 328226
rect 559682 328170 559738 328226
rect 559558 328046 559614 328102
rect 559682 328046 559738 328102
rect 559558 327922 559614 327978
rect 559682 327922 559738 327978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 359878 316294 359934 316350
rect 360002 316294 360058 316350
rect 359878 316170 359934 316226
rect 360002 316170 360058 316226
rect 359878 316046 359934 316102
rect 360002 316046 360058 316102
rect 359878 315922 359934 315978
rect 360002 315922 360058 315978
rect 390598 316294 390654 316350
rect 390722 316294 390778 316350
rect 390598 316170 390654 316226
rect 390722 316170 390778 316226
rect 390598 316046 390654 316102
rect 390722 316046 390778 316102
rect 390598 315922 390654 315978
rect 390722 315922 390778 315978
rect 421318 316294 421374 316350
rect 421442 316294 421498 316350
rect 421318 316170 421374 316226
rect 421442 316170 421498 316226
rect 421318 316046 421374 316102
rect 421442 316046 421498 316102
rect 421318 315922 421374 315978
rect 421442 315922 421498 315978
rect 452038 316294 452094 316350
rect 452162 316294 452218 316350
rect 452038 316170 452094 316226
rect 452162 316170 452218 316226
rect 452038 316046 452094 316102
rect 452162 316046 452218 316102
rect 452038 315922 452094 315978
rect 452162 315922 452218 315978
rect 482758 316294 482814 316350
rect 482882 316294 482938 316350
rect 482758 316170 482814 316226
rect 482882 316170 482938 316226
rect 482758 316046 482814 316102
rect 482882 316046 482938 316102
rect 482758 315922 482814 315978
rect 482882 315922 482938 315978
rect 513478 316294 513534 316350
rect 513602 316294 513658 316350
rect 513478 316170 513534 316226
rect 513602 316170 513658 316226
rect 513478 316046 513534 316102
rect 513602 316046 513658 316102
rect 513478 315922 513534 315978
rect 513602 315922 513658 315978
rect 544198 316294 544254 316350
rect 544322 316294 544378 316350
rect 544198 316170 544254 316226
rect 544322 316170 544378 316226
rect 544198 316046 544254 316102
rect 544322 316046 544378 316102
rect 544198 315922 544254 315978
rect 544322 315922 544378 315978
rect 574918 316294 574974 316350
rect 575042 316294 575098 316350
rect 574918 316170 574974 316226
rect 575042 316170 575098 316226
rect 574918 316046 574974 316102
rect 575042 316046 575098 316102
rect 574918 315922 574974 315978
rect 575042 315922 575098 315978
rect 344518 310294 344574 310350
rect 344642 310294 344698 310350
rect 344518 310170 344574 310226
rect 344642 310170 344698 310226
rect 344518 310046 344574 310102
rect 344642 310046 344698 310102
rect 344518 309922 344574 309978
rect 344642 309922 344698 309978
rect 375238 310294 375294 310350
rect 375362 310294 375418 310350
rect 375238 310170 375294 310226
rect 375362 310170 375418 310226
rect 375238 310046 375294 310102
rect 375362 310046 375418 310102
rect 375238 309922 375294 309978
rect 375362 309922 375418 309978
rect 405958 310294 406014 310350
rect 406082 310294 406138 310350
rect 405958 310170 406014 310226
rect 406082 310170 406138 310226
rect 405958 310046 406014 310102
rect 406082 310046 406138 310102
rect 405958 309922 406014 309978
rect 406082 309922 406138 309978
rect 436678 310294 436734 310350
rect 436802 310294 436858 310350
rect 436678 310170 436734 310226
rect 436802 310170 436858 310226
rect 436678 310046 436734 310102
rect 436802 310046 436858 310102
rect 436678 309922 436734 309978
rect 436802 309922 436858 309978
rect 467398 310294 467454 310350
rect 467522 310294 467578 310350
rect 467398 310170 467454 310226
rect 467522 310170 467578 310226
rect 467398 310046 467454 310102
rect 467522 310046 467578 310102
rect 467398 309922 467454 309978
rect 467522 309922 467578 309978
rect 498118 310294 498174 310350
rect 498242 310294 498298 310350
rect 498118 310170 498174 310226
rect 498242 310170 498298 310226
rect 498118 310046 498174 310102
rect 498242 310046 498298 310102
rect 498118 309922 498174 309978
rect 498242 309922 498298 309978
rect 528838 310294 528894 310350
rect 528962 310294 529018 310350
rect 528838 310170 528894 310226
rect 528962 310170 529018 310226
rect 528838 310046 528894 310102
rect 528962 310046 529018 310102
rect 528838 309922 528894 309978
rect 528962 309922 529018 309978
rect 559558 310294 559614 310350
rect 559682 310294 559738 310350
rect 559558 310170 559614 310226
rect 559682 310170 559738 310226
rect 559558 310046 559614 310102
rect 559682 310046 559738 310102
rect 559558 309922 559614 309978
rect 559682 309922 559738 309978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 341068 301562 341124 301618
rect 340844 157382 340900 157438
rect 340956 294542 341012 294598
rect 359878 298294 359934 298350
rect 360002 298294 360058 298350
rect 359878 298170 359934 298226
rect 360002 298170 360058 298226
rect 359878 298046 359934 298102
rect 360002 298046 360058 298102
rect 359878 297922 359934 297978
rect 360002 297922 360058 297978
rect 390598 298294 390654 298350
rect 390722 298294 390778 298350
rect 390598 298170 390654 298226
rect 390722 298170 390778 298226
rect 390598 298046 390654 298102
rect 390722 298046 390778 298102
rect 390598 297922 390654 297978
rect 390722 297922 390778 297978
rect 421318 298294 421374 298350
rect 421442 298294 421498 298350
rect 421318 298170 421374 298226
rect 421442 298170 421498 298226
rect 421318 298046 421374 298102
rect 421442 298046 421498 298102
rect 421318 297922 421374 297978
rect 421442 297922 421498 297978
rect 452038 298294 452094 298350
rect 452162 298294 452218 298350
rect 452038 298170 452094 298226
rect 452162 298170 452218 298226
rect 452038 298046 452094 298102
rect 452162 298046 452218 298102
rect 452038 297922 452094 297978
rect 452162 297922 452218 297978
rect 482758 298294 482814 298350
rect 482882 298294 482938 298350
rect 482758 298170 482814 298226
rect 482882 298170 482938 298226
rect 482758 298046 482814 298102
rect 482882 298046 482938 298102
rect 482758 297922 482814 297978
rect 482882 297922 482938 297978
rect 513478 298294 513534 298350
rect 513602 298294 513658 298350
rect 513478 298170 513534 298226
rect 513602 298170 513658 298226
rect 513478 298046 513534 298102
rect 513602 298046 513658 298102
rect 513478 297922 513534 297978
rect 513602 297922 513658 297978
rect 544198 298294 544254 298350
rect 544322 298294 544378 298350
rect 544198 298170 544254 298226
rect 544322 298170 544378 298226
rect 544198 298046 544254 298102
rect 544322 298046 544378 298102
rect 544198 297922 544254 297978
rect 544322 297922 544378 297978
rect 574918 298294 574974 298350
rect 575042 298294 575098 298350
rect 574918 298170 574974 298226
rect 575042 298170 575098 298226
rect 574918 298046 574974 298102
rect 575042 298046 575098 298102
rect 574918 297922 574974 297978
rect 575042 297922 575098 297978
rect 344518 292294 344574 292350
rect 344642 292294 344698 292350
rect 344518 292170 344574 292226
rect 344642 292170 344698 292226
rect 344518 292046 344574 292102
rect 344642 292046 344698 292102
rect 344518 291922 344574 291978
rect 344642 291922 344698 291978
rect 375238 292294 375294 292350
rect 375362 292294 375418 292350
rect 375238 292170 375294 292226
rect 375362 292170 375418 292226
rect 375238 292046 375294 292102
rect 375362 292046 375418 292102
rect 375238 291922 375294 291978
rect 375362 291922 375418 291978
rect 405958 292294 406014 292350
rect 406082 292294 406138 292350
rect 405958 292170 406014 292226
rect 406082 292170 406138 292226
rect 405958 292046 406014 292102
rect 406082 292046 406138 292102
rect 405958 291922 406014 291978
rect 406082 291922 406138 291978
rect 436678 292294 436734 292350
rect 436802 292294 436858 292350
rect 436678 292170 436734 292226
rect 436802 292170 436858 292226
rect 436678 292046 436734 292102
rect 436802 292046 436858 292102
rect 436678 291922 436734 291978
rect 436802 291922 436858 291978
rect 467398 292294 467454 292350
rect 467522 292294 467578 292350
rect 467398 292170 467454 292226
rect 467522 292170 467578 292226
rect 467398 292046 467454 292102
rect 467522 292046 467578 292102
rect 467398 291922 467454 291978
rect 467522 291922 467578 291978
rect 498118 292294 498174 292350
rect 498242 292294 498298 292350
rect 498118 292170 498174 292226
rect 498242 292170 498298 292226
rect 498118 292046 498174 292102
rect 498242 292046 498298 292102
rect 498118 291922 498174 291978
rect 498242 291922 498298 291978
rect 528838 292294 528894 292350
rect 528962 292294 529018 292350
rect 528838 292170 528894 292226
rect 528962 292170 529018 292226
rect 528838 292046 528894 292102
rect 528962 292046 529018 292102
rect 528838 291922 528894 291978
rect 528962 291922 529018 291978
rect 559558 292294 559614 292350
rect 559682 292294 559738 292350
rect 559558 292170 559614 292226
rect 559682 292170 559738 292226
rect 559558 292046 559614 292102
rect 559682 292046 559738 292102
rect 559558 291922 559614 291978
rect 559682 291922 559738 291978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 341068 283742 341124 283798
rect 341292 283922 341348 283978
rect 341068 243422 341124 243478
rect 359878 280294 359934 280350
rect 360002 280294 360058 280350
rect 359878 280170 359934 280226
rect 360002 280170 360058 280226
rect 359878 280046 359934 280102
rect 360002 280046 360058 280102
rect 359878 279922 359934 279978
rect 360002 279922 360058 279978
rect 390598 280294 390654 280350
rect 390722 280294 390778 280350
rect 390598 280170 390654 280226
rect 390722 280170 390778 280226
rect 390598 280046 390654 280102
rect 390722 280046 390778 280102
rect 390598 279922 390654 279978
rect 390722 279922 390778 279978
rect 421318 280294 421374 280350
rect 421442 280294 421498 280350
rect 421318 280170 421374 280226
rect 421442 280170 421498 280226
rect 421318 280046 421374 280102
rect 421442 280046 421498 280102
rect 421318 279922 421374 279978
rect 421442 279922 421498 279978
rect 452038 280294 452094 280350
rect 452162 280294 452218 280350
rect 452038 280170 452094 280226
rect 452162 280170 452218 280226
rect 452038 280046 452094 280102
rect 452162 280046 452218 280102
rect 452038 279922 452094 279978
rect 452162 279922 452218 279978
rect 482758 280294 482814 280350
rect 482882 280294 482938 280350
rect 482758 280170 482814 280226
rect 482882 280170 482938 280226
rect 482758 280046 482814 280102
rect 482882 280046 482938 280102
rect 482758 279922 482814 279978
rect 482882 279922 482938 279978
rect 513478 280294 513534 280350
rect 513602 280294 513658 280350
rect 513478 280170 513534 280226
rect 513602 280170 513658 280226
rect 513478 280046 513534 280102
rect 513602 280046 513658 280102
rect 513478 279922 513534 279978
rect 513602 279922 513658 279978
rect 544198 280294 544254 280350
rect 544322 280294 544378 280350
rect 544198 280170 544254 280226
rect 544322 280170 544378 280226
rect 544198 280046 544254 280102
rect 544322 280046 544378 280102
rect 544198 279922 544254 279978
rect 544322 279922 544378 279978
rect 574918 280294 574974 280350
rect 575042 280294 575098 280350
rect 574918 280170 574974 280226
rect 575042 280170 575098 280226
rect 574918 280046 574974 280102
rect 575042 280046 575098 280102
rect 574918 279922 574974 279978
rect 575042 279922 575098 279978
rect 344518 274294 344574 274350
rect 344642 274294 344698 274350
rect 344518 274170 344574 274226
rect 344642 274170 344698 274226
rect 344518 274046 344574 274102
rect 344642 274046 344698 274102
rect 344518 273922 344574 273978
rect 344642 273922 344698 273978
rect 375238 274294 375294 274350
rect 375362 274294 375418 274350
rect 375238 274170 375294 274226
rect 375362 274170 375418 274226
rect 375238 274046 375294 274102
rect 375362 274046 375418 274102
rect 375238 273922 375294 273978
rect 375362 273922 375418 273978
rect 405958 274294 406014 274350
rect 406082 274294 406138 274350
rect 405958 274170 406014 274226
rect 406082 274170 406138 274226
rect 405958 274046 406014 274102
rect 406082 274046 406138 274102
rect 405958 273922 406014 273978
rect 406082 273922 406138 273978
rect 436678 274294 436734 274350
rect 436802 274294 436858 274350
rect 436678 274170 436734 274226
rect 436802 274170 436858 274226
rect 436678 274046 436734 274102
rect 436802 274046 436858 274102
rect 436678 273922 436734 273978
rect 436802 273922 436858 273978
rect 467398 274294 467454 274350
rect 467522 274294 467578 274350
rect 467398 274170 467454 274226
rect 467522 274170 467578 274226
rect 467398 274046 467454 274102
rect 467522 274046 467578 274102
rect 467398 273922 467454 273978
rect 467522 273922 467578 273978
rect 498118 274294 498174 274350
rect 498242 274294 498298 274350
rect 498118 274170 498174 274226
rect 498242 274170 498298 274226
rect 498118 274046 498174 274102
rect 498242 274046 498298 274102
rect 498118 273922 498174 273978
rect 498242 273922 498298 273978
rect 528838 274294 528894 274350
rect 528962 274294 529018 274350
rect 528838 274170 528894 274226
rect 528962 274170 529018 274226
rect 528838 274046 528894 274102
rect 528962 274046 529018 274102
rect 528838 273922 528894 273978
rect 528962 273922 529018 273978
rect 559558 274294 559614 274350
rect 559682 274294 559738 274350
rect 559558 274170 559614 274226
rect 559682 274170 559738 274226
rect 559558 274046 559614 274102
rect 559682 274046 559738 274102
rect 559558 273922 559614 273978
rect 559682 273922 559738 273978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 359878 262294 359934 262350
rect 360002 262294 360058 262350
rect 359878 262170 359934 262226
rect 360002 262170 360058 262226
rect 359878 262046 359934 262102
rect 360002 262046 360058 262102
rect 359878 261922 359934 261978
rect 360002 261922 360058 261978
rect 390598 262294 390654 262350
rect 390722 262294 390778 262350
rect 390598 262170 390654 262226
rect 390722 262170 390778 262226
rect 390598 262046 390654 262102
rect 390722 262046 390778 262102
rect 390598 261922 390654 261978
rect 390722 261922 390778 261978
rect 421318 262294 421374 262350
rect 421442 262294 421498 262350
rect 421318 262170 421374 262226
rect 421442 262170 421498 262226
rect 421318 262046 421374 262102
rect 421442 262046 421498 262102
rect 421318 261922 421374 261978
rect 421442 261922 421498 261978
rect 452038 262294 452094 262350
rect 452162 262294 452218 262350
rect 452038 262170 452094 262226
rect 452162 262170 452218 262226
rect 452038 262046 452094 262102
rect 452162 262046 452218 262102
rect 452038 261922 452094 261978
rect 452162 261922 452218 261978
rect 482758 262294 482814 262350
rect 482882 262294 482938 262350
rect 482758 262170 482814 262226
rect 482882 262170 482938 262226
rect 482758 262046 482814 262102
rect 482882 262046 482938 262102
rect 482758 261922 482814 261978
rect 482882 261922 482938 261978
rect 513478 262294 513534 262350
rect 513602 262294 513658 262350
rect 513478 262170 513534 262226
rect 513602 262170 513658 262226
rect 513478 262046 513534 262102
rect 513602 262046 513658 262102
rect 513478 261922 513534 261978
rect 513602 261922 513658 261978
rect 544198 262294 544254 262350
rect 544322 262294 544378 262350
rect 544198 262170 544254 262226
rect 544322 262170 544378 262226
rect 544198 262046 544254 262102
rect 544322 262046 544378 262102
rect 544198 261922 544254 261978
rect 544322 261922 544378 261978
rect 574918 262294 574974 262350
rect 575042 262294 575098 262350
rect 574918 262170 574974 262226
rect 575042 262170 575098 262226
rect 574918 262046 574974 262102
rect 575042 262046 575098 262102
rect 574918 261922 574974 261978
rect 575042 261922 575098 261978
rect 344518 256294 344574 256350
rect 344642 256294 344698 256350
rect 344518 256170 344574 256226
rect 344642 256170 344698 256226
rect 344518 256046 344574 256102
rect 344642 256046 344698 256102
rect 344518 255922 344574 255978
rect 344642 255922 344698 255978
rect 375238 256294 375294 256350
rect 375362 256294 375418 256350
rect 375238 256170 375294 256226
rect 375362 256170 375418 256226
rect 375238 256046 375294 256102
rect 375362 256046 375418 256102
rect 375238 255922 375294 255978
rect 375362 255922 375418 255978
rect 405958 256294 406014 256350
rect 406082 256294 406138 256350
rect 405958 256170 406014 256226
rect 406082 256170 406138 256226
rect 405958 256046 406014 256102
rect 406082 256046 406138 256102
rect 405958 255922 406014 255978
rect 406082 255922 406138 255978
rect 436678 256294 436734 256350
rect 436802 256294 436858 256350
rect 436678 256170 436734 256226
rect 436802 256170 436858 256226
rect 436678 256046 436734 256102
rect 436802 256046 436858 256102
rect 436678 255922 436734 255978
rect 436802 255922 436858 255978
rect 467398 256294 467454 256350
rect 467522 256294 467578 256350
rect 467398 256170 467454 256226
rect 467522 256170 467578 256226
rect 467398 256046 467454 256102
rect 467522 256046 467578 256102
rect 467398 255922 467454 255978
rect 467522 255922 467578 255978
rect 498118 256294 498174 256350
rect 498242 256294 498298 256350
rect 498118 256170 498174 256226
rect 498242 256170 498298 256226
rect 498118 256046 498174 256102
rect 498242 256046 498298 256102
rect 498118 255922 498174 255978
rect 498242 255922 498298 255978
rect 528838 256294 528894 256350
rect 528962 256294 529018 256350
rect 528838 256170 528894 256226
rect 528962 256170 529018 256226
rect 528838 256046 528894 256102
rect 528962 256046 529018 256102
rect 528838 255922 528894 255978
rect 528962 255922 529018 255978
rect 559558 256294 559614 256350
rect 559682 256294 559738 256350
rect 559558 256170 559614 256226
rect 559682 256170 559738 256226
rect 559558 256046 559614 256102
rect 559682 256046 559738 256102
rect 559558 255922 559614 255978
rect 559682 255922 559738 255978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 359878 244294 359934 244350
rect 360002 244294 360058 244350
rect 359878 244170 359934 244226
rect 360002 244170 360058 244226
rect 359878 244046 359934 244102
rect 360002 244046 360058 244102
rect 359878 243922 359934 243978
rect 360002 243922 360058 243978
rect 390598 244294 390654 244350
rect 390722 244294 390778 244350
rect 390598 244170 390654 244226
rect 390722 244170 390778 244226
rect 390598 244046 390654 244102
rect 390722 244046 390778 244102
rect 390598 243922 390654 243978
rect 390722 243922 390778 243978
rect 421318 244294 421374 244350
rect 421442 244294 421498 244350
rect 421318 244170 421374 244226
rect 421442 244170 421498 244226
rect 421318 244046 421374 244102
rect 421442 244046 421498 244102
rect 421318 243922 421374 243978
rect 421442 243922 421498 243978
rect 452038 244294 452094 244350
rect 452162 244294 452218 244350
rect 452038 244170 452094 244226
rect 452162 244170 452218 244226
rect 452038 244046 452094 244102
rect 452162 244046 452218 244102
rect 452038 243922 452094 243978
rect 452162 243922 452218 243978
rect 482758 244294 482814 244350
rect 482882 244294 482938 244350
rect 482758 244170 482814 244226
rect 482882 244170 482938 244226
rect 482758 244046 482814 244102
rect 482882 244046 482938 244102
rect 482758 243922 482814 243978
rect 482882 243922 482938 243978
rect 513478 244294 513534 244350
rect 513602 244294 513658 244350
rect 513478 244170 513534 244226
rect 513602 244170 513658 244226
rect 513478 244046 513534 244102
rect 513602 244046 513658 244102
rect 513478 243922 513534 243978
rect 513602 243922 513658 243978
rect 544198 244294 544254 244350
rect 544322 244294 544378 244350
rect 544198 244170 544254 244226
rect 544322 244170 544378 244226
rect 544198 244046 544254 244102
rect 544322 244046 544378 244102
rect 544198 243922 544254 243978
rect 544322 243922 544378 243978
rect 574918 244294 574974 244350
rect 575042 244294 575098 244350
rect 574918 244170 574974 244226
rect 575042 244170 575098 244226
rect 574918 244046 574974 244102
rect 575042 244046 575098 244102
rect 574918 243922 574974 243978
rect 575042 243922 575098 243978
rect 341292 239282 341348 239338
rect 344518 238294 344574 238350
rect 344642 238294 344698 238350
rect 344518 238170 344574 238226
rect 344642 238170 344698 238226
rect 344518 238046 344574 238102
rect 344642 238046 344698 238102
rect 344518 237922 344574 237978
rect 344642 237922 344698 237978
rect 375238 238294 375294 238350
rect 375362 238294 375418 238350
rect 375238 238170 375294 238226
rect 375362 238170 375418 238226
rect 375238 238046 375294 238102
rect 375362 238046 375418 238102
rect 375238 237922 375294 237978
rect 375362 237922 375418 237978
rect 405958 238294 406014 238350
rect 406082 238294 406138 238350
rect 405958 238170 406014 238226
rect 406082 238170 406138 238226
rect 405958 238046 406014 238102
rect 406082 238046 406138 238102
rect 405958 237922 406014 237978
rect 406082 237922 406138 237978
rect 436678 238294 436734 238350
rect 436802 238294 436858 238350
rect 436678 238170 436734 238226
rect 436802 238170 436858 238226
rect 436678 238046 436734 238102
rect 436802 238046 436858 238102
rect 436678 237922 436734 237978
rect 436802 237922 436858 237978
rect 467398 238294 467454 238350
rect 467522 238294 467578 238350
rect 467398 238170 467454 238226
rect 467522 238170 467578 238226
rect 467398 238046 467454 238102
rect 467522 238046 467578 238102
rect 467398 237922 467454 237978
rect 467522 237922 467578 237978
rect 498118 238294 498174 238350
rect 498242 238294 498298 238350
rect 498118 238170 498174 238226
rect 498242 238170 498298 238226
rect 498118 238046 498174 238102
rect 498242 238046 498298 238102
rect 498118 237922 498174 237978
rect 498242 237922 498298 237978
rect 528838 238294 528894 238350
rect 528962 238294 529018 238350
rect 528838 238170 528894 238226
rect 528962 238170 529018 238226
rect 528838 238046 528894 238102
rect 528962 238046 529018 238102
rect 528838 237922 528894 237978
rect 528962 237922 529018 237978
rect 559558 238294 559614 238350
rect 559682 238294 559738 238350
rect 559558 238170 559614 238226
rect 559682 238170 559738 238226
rect 559558 238046 559614 238102
rect 559682 238046 559738 238102
rect 559558 237922 559614 237978
rect 559682 237922 559738 237978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 341068 236042 341124 236098
rect 359878 226294 359934 226350
rect 360002 226294 360058 226350
rect 359878 226170 359934 226226
rect 360002 226170 360058 226226
rect 359878 226046 359934 226102
rect 360002 226046 360058 226102
rect 359878 225922 359934 225978
rect 360002 225922 360058 225978
rect 390598 226294 390654 226350
rect 390722 226294 390778 226350
rect 390598 226170 390654 226226
rect 390722 226170 390778 226226
rect 390598 226046 390654 226102
rect 390722 226046 390778 226102
rect 390598 225922 390654 225978
rect 390722 225922 390778 225978
rect 421318 226294 421374 226350
rect 421442 226294 421498 226350
rect 421318 226170 421374 226226
rect 421442 226170 421498 226226
rect 421318 226046 421374 226102
rect 421442 226046 421498 226102
rect 421318 225922 421374 225978
rect 421442 225922 421498 225978
rect 452038 226294 452094 226350
rect 452162 226294 452218 226350
rect 452038 226170 452094 226226
rect 452162 226170 452218 226226
rect 452038 226046 452094 226102
rect 452162 226046 452218 226102
rect 452038 225922 452094 225978
rect 452162 225922 452218 225978
rect 482758 226294 482814 226350
rect 482882 226294 482938 226350
rect 482758 226170 482814 226226
rect 482882 226170 482938 226226
rect 482758 226046 482814 226102
rect 482882 226046 482938 226102
rect 482758 225922 482814 225978
rect 482882 225922 482938 225978
rect 513478 226294 513534 226350
rect 513602 226294 513658 226350
rect 513478 226170 513534 226226
rect 513602 226170 513658 226226
rect 513478 226046 513534 226102
rect 513602 226046 513658 226102
rect 513478 225922 513534 225978
rect 513602 225922 513658 225978
rect 544198 226294 544254 226350
rect 544322 226294 544378 226350
rect 544198 226170 544254 226226
rect 544322 226170 544378 226226
rect 544198 226046 544254 226102
rect 544322 226046 544378 226102
rect 544198 225922 544254 225978
rect 544322 225922 544378 225978
rect 574918 226294 574974 226350
rect 575042 226294 575098 226350
rect 574918 226170 574974 226226
rect 575042 226170 575098 226226
rect 574918 226046 574974 226102
rect 575042 226046 575098 226102
rect 574918 225922 574974 225978
rect 575042 225922 575098 225978
rect 344518 220294 344574 220350
rect 344642 220294 344698 220350
rect 344518 220170 344574 220226
rect 344642 220170 344698 220226
rect 344518 220046 344574 220102
rect 344642 220046 344698 220102
rect 344518 219922 344574 219978
rect 344642 219922 344698 219978
rect 375238 220294 375294 220350
rect 375362 220294 375418 220350
rect 375238 220170 375294 220226
rect 375362 220170 375418 220226
rect 375238 220046 375294 220102
rect 375362 220046 375418 220102
rect 375238 219922 375294 219978
rect 375362 219922 375418 219978
rect 405958 220294 406014 220350
rect 406082 220294 406138 220350
rect 405958 220170 406014 220226
rect 406082 220170 406138 220226
rect 405958 220046 406014 220102
rect 406082 220046 406138 220102
rect 405958 219922 406014 219978
rect 406082 219922 406138 219978
rect 436678 220294 436734 220350
rect 436802 220294 436858 220350
rect 436678 220170 436734 220226
rect 436802 220170 436858 220226
rect 436678 220046 436734 220102
rect 436802 220046 436858 220102
rect 436678 219922 436734 219978
rect 436802 219922 436858 219978
rect 467398 220294 467454 220350
rect 467522 220294 467578 220350
rect 467398 220170 467454 220226
rect 467522 220170 467578 220226
rect 467398 220046 467454 220102
rect 467522 220046 467578 220102
rect 467398 219922 467454 219978
rect 467522 219922 467578 219978
rect 498118 220294 498174 220350
rect 498242 220294 498298 220350
rect 498118 220170 498174 220226
rect 498242 220170 498298 220226
rect 498118 220046 498174 220102
rect 498242 220046 498298 220102
rect 498118 219922 498174 219978
rect 498242 219922 498298 219978
rect 528838 220294 528894 220350
rect 528962 220294 529018 220350
rect 528838 220170 528894 220226
rect 528962 220170 529018 220226
rect 528838 220046 528894 220102
rect 528962 220046 529018 220102
rect 528838 219922 528894 219978
rect 528962 219922 529018 219978
rect 559558 220294 559614 220350
rect 559682 220294 559738 220350
rect 559558 220170 559614 220226
rect 559682 220170 559738 220226
rect 559558 220046 559614 220102
rect 559682 220046 559738 220102
rect 559558 219922 559614 219978
rect 559682 219922 559738 219978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 359878 208294 359934 208350
rect 360002 208294 360058 208350
rect 359878 208170 359934 208226
rect 360002 208170 360058 208226
rect 359878 208046 359934 208102
rect 360002 208046 360058 208102
rect 359878 207922 359934 207978
rect 360002 207922 360058 207978
rect 390598 208294 390654 208350
rect 390722 208294 390778 208350
rect 390598 208170 390654 208226
rect 390722 208170 390778 208226
rect 390598 208046 390654 208102
rect 390722 208046 390778 208102
rect 390598 207922 390654 207978
rect 390722 207922 390778 207978
rect 421318 208294 421374 208350
rect 421442 208294 421498 208350
rect 421318 208170 421374 208226
rect 421442 208170 421498 208226
rect 421318 208046 421374 208102
rect 421442 208046 421498 208102
rect 421318 207922 421374 207978
rect 421442 207922 421498 207978
rect 452038 208294 452094 208350
rect 452162 208294 452218 208350
rect 452038 208170 452094 208226
rect 452162 208170 452218 208226
rect 452038 208046 452094 208102
rect 452162 208046 452218 208102
rect 452038 207922 452094 207978
rect 452162 207922 452218 207978
rect 482758 208294 482814 208350
rect 482882 208294 482938 208350
rect 482758 208170 482814 208226
rect 482882 208170 482938 208226
rect 482758 208046 482814 208102
rect 482882 208046 482938 208102
rect 482758 207922 482814 207978
rect 482882 207922 482938 207978
rect 513478 208294 513534 208350
rect 513602 208294 513658 208350
rect 513478 208170 513534 208226
rect 513602 208170 513658 208226
rect 513478 208046 513534 208102
rect 513602 208046 513658 208102
rect 513478 207922 513534 207978
rect 513602 207922 513658 207978
rect 544198 208294 544254 208350
rect 544322 208294 544378 208350
rect 544198 208170 544254 208226
rect 544322 208170 544378 208226
rect 544198 208046 544254 208102
rect 544322 208046 544378 208102
rect 544198 207922 544254 207978
rect 544322 207922 544378 207978
rect 574918 208294 574974 208350
rect 575042 208294 575098 208350
rect 574918 208170 574974 208226
rect 575042 208170 575098 208226
rect 574918 208046 574974 208102
rect 575042 208046 575098 208102
rect 574918 207922 574974 207978
rect 575042 207922 575098 207978
rect 344518 202294 344574 202350
rect 344642 202294 344698 202350
rect 344518 202170 344574 202226
rect 344642 202170 344698 202226
rect 344518 202046 344574 202102
rect 344642 202046 344698 202102
rect 344518 201922 344574 201978
rect 344642 201922 344698 201978
rect 375238 202294 375294 202350
rect 375362 202294 375418 202350
rect 375238 202170 375294 202226
rect 375362 202170 375418 202226
rect 375238 202046 375294 202102
rect 375362 202046 375418 202102
rect 375238 201922 375294 201978
rect 375362 201922 375418 201978
rect 405958 202294 406014 202350
rect 406082 202294 406138 202350
rect 405958 202170 406014 202226
rect 406082 202170 406138 202226
rect 405958 202046 406014 202102
rect 406082 202046 406138 202102
rect 405958 201922 406014 201978
rect 406082 201922 406138 201978
rect 436678 202294 436734 202350
rect 436802 202294 436858 202350
rect 436678 202170 436734 202226
rect 436802 202170 436858 202226
rect 436678 202046 436734 202102
rect 436802 202046 436858 202102
rect 436678 201922 436734 201978
rect 436802 201922 436858 201978
rect 467398 202294 467454 202350
rect 467522 202294 467578 202350
rect 467398 202170 467454 202226
rect 467522 202170 467578 202226
rect 467398 202046 467454 202102
rect 467522 202046 467578 202102
rect 467398 201922 467454 201978
rect 467522 201922 467578 201978
rect 498118 202294 498174 202350
rect 498242 202294 498298 202350
rect 498118 202170 498174 202226
rect 498242 202170 498298 202226
rect 498118 202046 498174 202102
rect 498242 202046 498298 202102
rect 498118 201922 498174 201978
rect 498242 201922 498298 201978
rect 528838 202294 528894 202350
rect 528962 202294 529018 202350
rect 528838 202170 528894 202226
rect 528962 202170 529018 202226
rect 528838 202046 528894 202102
rect 528962 202046 529018 202102
rect 528838 201922 528894 201978
rect 528962 201922 529018 201978
rect 559558 202294 559614 202350
rect 559682 202294 559738 202350
rect 559558 202170 559614 202226
rect 559682 202170 559738 202226
rect 559558 202046 559614 202102
rect 559682 202046 559738 202102
rect 559558 201922 559614 201978
rect 559682 201922 559738 201978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 359878 190294 359934 190350
rect 360002 190294 360058 190350
rect 359878 190170 359934 190226
rect 360002 190170 360058 190226
rect 359878 190046 359934 190102
rect 360002 190046 360058 190102
rect 359878 189922 359934 189978
rect 360002 189922 360058 189978
rect 390598 190294 390654 190350
rect 390722 190294 390778 190350
rect 390598 190170 390654 190226
rect 390722 190170 390778 190226
rect 390598 190046 390654 190102
rect 390722 190046 390778 190102
rect 390598 189922 390654 189978
rect 390722 189922 390778 189978
rect 421318 190294 421374 190350
rect 421442 190294 421498 190350
rect 421318 190170 421374 190226
rect 421442 190170 421498 190226
rect 421318 190046 421374 190102
rect 421442 190046 421498 190102
rect 421318 189922 421374 189978
rect 421442 189922 421498 189978
rect 452038 190294 452094 190350
rect 452162 190294 452218 190350
rect 452038 190170 452094 190226
rect 452162 190170 452218 190226
rect 452038 190046 452094 190102
rect 452162 190046 452218 190102
rect 452038 189922 452094 189978
rect 452162 189922 452218 189978
rect 482758 190294 482814 190350
rect 482882 190294 482938 190350
rect 482758 190170 482814 190226
rect 482882 190170 482938 190226
rect 482758 190046 482814 190102
rect 482882 190046 482938 190102
rect 482758 189922 482814 189978
rect 482882 189922 482938 189978
rect 513478 190294 513534 190350
rect 513602 190294 513658 190350
rect 513478 190170 513534 190226
rect 513602 190170 513658 190226
rect 513478 190046 513534 190102
rect 513602 190046 513658 190102
rect 513478 189922 513534 189978
rect 513602 189922 513658 189978
rect 544198 190294 544254 190350
rect 544322 190294 544378 190350
rect 544198 190170 544254 190226
rect 544322 190170 544378 190226
rect 544198 190046 544254 190102
rect 544322 190046 544378 190102
rect 544198 189922 544254 189978
rect 544322 189922 544378 189978
rect 574918 190294 574974 190350
rect 575042 190294 575098 190350
rect 574918 190170 574974 190226
rect 575042 190170 575098 190226
rect 574918 190046 574974 190102
rect 575042 190046 575098 190102
rect 574918 189922 574974 189978
rect 575042 189922 575098 189978
rect 344518 184294 344574 184350
rect 344642 184294 344698 184350
rect 344518 184170 344574 184226
rect 344642 184170 344698 184226
rect 344518 184046 344574 184102
rect 344642 184046 344698 184102
rect 344518 183922 344574 183978
rect 344642 183922 344698 183978
rect 375238 184294 375294 184350
rect 375362 184294 375418 184350
rect 375238 184170 375294 184226
rect 375362 184170 375418 184226
rect 375238 184046 375294 184102
rect 375362 184046 375418 184102
rect 375238 183922 375294 183978
rect 375362 183922 375418 183978
rect 405958 184294 406014 184350
rect 406082 184294 406138 184350
rect 405958 184170 406014 184226
rect 406082 184170 406138 184226
rect 405958 184046 406014 184102
rect 406082 184046 406138 184102
rect 405958 183922 406014 183978
rect 406082 183922 406138 183978
rect 436678 184294 436734 184350
rect 436802 184294 436858 184350
rect 436678 184170 436734 184226
rect 436802 184170 436858 184226
rect 436678 184046 436734 184102
rect 436802 184046 436858 184102
rect 436678 183922 436734 183978
rect 436802 183922 436858 183978
rect 467398 184294 467454 184350
rect 467522 184294 467578 184350
rect 467398 184170 467454 184226
rect 467522 184170 467578 184226
rect 467398 184046 467454 184102
rect 467522 184046 467578 184102
rect 467398 183922 467454 183978
rect 467522 183922 467578 183978
rect 498118 184294 498174 184350
rect 498242 184294 498298 184350
rect 498118 184170 498174 184226
rect 498242 184170 498298 184226
rect 498118 184046 498174 184102
rect 498242 184046 498298 184102
rect 498118 183922 498174 183978
rect 498242 183922 498298 183978
rect 528838 184294 528894 184350
rect 528962 184294 529018 184350
rect 528838 184170 528894 184226
rect 528962 184170 529018 184226
rect 528838 184046 528894 184102
rect 528962 184046 529018 184102
rect 528838 183922 528894 183978
rect 528962 183922 529018 183978
rect 559558 184294 559614 184350
rect 559682 184294 559738 184350
rect 559558 184170 559614 184226
rect 559682 184170 559738 184226
rect 559558 184046 559614 184102
rect 559682 184046 559738 184102
rect 559558 183922 559614 183978
rect 559682 183922 559738 183978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 341404 173042 341460 173098
rect 341292 168002 341348 168058
rect 341180 162242 341236 162298
rect 359878 172294 359934 172350
rect 360002 172294 360058 172350
rect 359878 172170 359934 172226
rect 360002 172170 360058 172226
rect 359878 172046 359934 172102
rect 360002 172046 360058 172102
rect 359878 171922 359934 171978
rect 360002 171922 360058 171978
rect 390598 172294 390654 172350
rect 390722 172294 390778 172350
rect 390598 172170 390654 172226
rect 390722 172170 390778 172226
rect 390598 172046 390654 172102
rect 390722 172046 390778 172102
rect 390598 171922 390654 171978
rect 390722 171922 390778 171978
rect 421318 172294 421374 172350
rect 421442 172294 421498 172350
rect 421318 172170 421374 172226
rect 421442 172170 421498 172226
rect 421318 172046 421374 172102
rect 421442 172046 421498 172102
rect 421318 171922 421374 171978
rect 421442 171922 421498 171978
rect 452038 172294 452094 172350
rect 452162 172294 452218 172350
rect 452038 172170 452094 172226
rect 452162 172170 452218 172226
rect 452038 172046 452094 172102
rect 452162 172046 452218 172102
rect 452038 171922 452094 171978
rect 452162 171922 452218 171978
rect 482758 172294 482814 172350
rect 482882 172294 482938 172350
rect 482758 172170 482814 172226
rect 482882 172170 482938 172226
rect 482758 172046 482814 172102
rect 482882 172046 482938 172102
rect 482758 171922 482814 171978
rect 482882 171922 482938 171978
rect 513478 172294 513534 172350
rect 513602 172294 513658 172350
rect 513478 172170 513534 172226
rect 513602 172170 513658 172226
rect 513478 172046 513534 172102
rect 513602 172046 513658 172102
rect 513478 171922 513534 171978
rect 513602 171922 513658 171978
rect 544198 172294 544254 172350
rect 544322 172294 544378 172350
rect 544198 172170 544254 172226
rect 544322 172170 544378 172226
rect 544198 172046 544254 172102
rect 544322 172046 544378 172102
rect 544198 171922 544254 171978
rect 544322 171922 544378 171978
rect 574918 172294 574974 172350
rect 575042 172294 575098 172350
rect 574918 172170 574974 172226
rect 575042 172170 575098 172226
rect 574918 172046 574974 172102
rect 575042 172046 575098 172102
rect 574918 171922 574974 171978
rect 575042 171922 575098 171978
rect 344518 166294 344574 166350
rect 344642 166294 344698 166350
rect 344518 166170 344574 166226
rect 344642 166170 344698 166226
rect 344518 166046 344574 166102
rect 344642 166046 344698 166102
rect 344518 165922 344574 165978
rect 344642 165922 344698 165978
rect 375238 166294 375294 166350
rect 375362 166294 375418 166350
rect 375238 166170 375294 166226
rect 375362 166170 375418 166226
rect 375238 166046 375294 166102
rect 375362 166046 375418 166102
rect 375238 165922 375294 165978
rect 375362 165922 375418 165978
rect 405958 166294 406014 166350
rect 406082 166294 406138 166350
rect 405958 166170 406014 166226
rect 406082 166170 406138 166226
rect 405958 166046 406014 166102
rect 406082 166046 406138 166102
rect 405958 165922 406014 165978
rect 406082 165922 406138 165978
rect 436678 166294 436734 166350
rect 436802 166294 436858 166350
rect 436678 166170 436734 166226
rect 436802 166170 436858 166226
rect 436678 166046 436734 166102
rect 436802 166046 436858 166102
rect 436678 165922 436734 165978
rect 436802 165922 436858 165978
rect 467398 166294 467454 166350
rect 467522 166294 467578 166350
rect 467398 166170 467454 166226
rect 467522 166170 467578 166226
rect 467398 166046 467454 166102
rect 467522 166046 467578 166102
rect 467398 165922 467454 165978
rect 467522 165922 467578 165978
rect 498118 166294 498174 166350
rect 498242 166294 498298 166350
rect 498118 166170 498174 166226
rect 498242 166170 498298 166226
rect 498118 166046 498174 166102
rect 498242 166046 498298 166102
rect 498118 165922 498174 165978
rect 498242 165922 498298 165978
rect 528838 166294 528894 166350
rect 528962 166294 529018 166350
rect 528838 166170 528894 166226
rect 528962 166170 529018 166226
rect 528838 166046 528894 166102
rect 528962 166046 529018 166102
rect 528838 165922 528894 165978
rect 528962 165922 529018 165978
rect 559558 166294 559614 166350
rect 559682 166294 559738 166350
rect 559558 166170 559614 166226
rect 559682 166170 559738 166226
rect 559558 166046 559614 166102
rect 559682 166046 559738 166102
rect 559558 165922 559614 165978
rect 559682 165922 559738 165978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 341516 162062 341572 162118
rect 357868 159542 357924 159598
rect 340956 138482 341012 138538
rect 343434 148294 343490 148350
rect 343558 148294 343614 148350
rect 343682 148294 343738 148350
rect 343806 148294 343862 148350
rect 343434 148170 343490 148226
rect 343558 148170 343614 148226
rect 343682 148170 343738 148226
rect 343806 148170 343862 148226
rect 343434 148046 343490 148102
rect 343558 148046 343614 148102
rect 343682 148046 343738 148102
rect 343806 148046 343862 148102
rect 343434 147922 343490 147978
rect 343558 147922 343614 147978
rect 343682 147922 343738 147978
rect 343806 147922 343862 147978
rect 343434 130294 343490 130350
rect 343558 130294 343614 130350
rect 343682 130294 343738 130350
rect 343806 130294 343862 130350
rect 343434 130170 343490 130226
rect 343558 130170 343614 130226
rect 343682 130170 343738 130226
rect 343806 130170 343862 130226
rect 343434 130046 343490 130102
rect 343558 130046 343614 130102
rect 343682 130046 343738 130102
rect 343806 130046 343862 130102
rect 343434 129922 343490 129978
rect 343558 129922 343614 129978
rect 343682 129922 343738 129978
rect 343806 129922 343862 129978
rect 343434 112294 343490 112350
rect 343558 112294 343614 112350
rect 343682 112294 343738 112350
rect 343806 112294 343862 112350
rect 343434 112170 343490 112226
rect 343558 112170 343614 112226
rect 343682 112170 343738 112226
rect 343806 112170 343862 112226
rect 343434 112046 343490 112102
rect 343558 112046 343614 112102
rect 343682 112046 343738 112102
rect 343806 112046 343862 112102
rect 343434 111922 343490 111978
rect 343558 111922 343614 111978
rect 343682 111922 343738 111978
rect 343806 111922 343862 111978
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 343434 76294 343490 76350
rect 343558 76294 343614 76350
rect 343682 76294 343738 76350
rect 343806 76294 343862 76350
rect 343434 76170 343490 76226
rect 343558 76170 343614 76226
rect 343682 76170 343738 76226
rect 343806 76170 343862 76226
rect 343434 76046 343490 76102
rect 343558 76046 343614 76102
rect 343682 76046 343738 76102
rect 343806 76046 343862 76102
rect 343434 75922 343490 75978
rect 343558 75922 343614 75978
rect 343682 75922 343738 75978
rect 343806 75922 343862 75978
rect 343434 58294 343490 58350
rect 343558 58294 343614 58350
rect 343682 58294 343738 58350
rect 343806 58294 343862 58350
rect 343434 58170 343490 58226
rect 343558 58170 343614 58226
rect 343682 58170 343738 58226
rect 343806 58170 343862 58226
rect 343434 58046 343490 58102
rect 343558 58046 343614 58102
rect 343682 58046 343738 58102
rect 343806 58046 343862 58102
rect 343434 57922 343490 57978
rect 343558 57922 343614 57978
rect 343682 57922 343738 57978
rect 343806 57922 343862 57978
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 347154 154294 347210 154350
rect 347278 154294 347334 154350
rect 347402 154294 347458 154350
rect 347526 154294 347582 154350
rect 347154 154170 347210 154226
rect 347278 154170 347334 154226
rect 347402 154170 347458 154226
rect 347526 154170 347582 154226
rect 347154 154046 347210 154102
rect 347278 154046 347334 154102
rect 347402 154046 347458 154102
rect 347526 154046 347582 154102
rect 347154 153922 347210 153978
rect 347278 153922 347334 153978
rect 347402 153922 347458 153978
rect 347526 153922 347582 153978
rect 347154 136294 347210 136350
rect 347278 136294 347334 136350
rect 347402 136294 347458 136350
rect 347526 136294 347582 136350
rect 347154 136170 347210 136226
rect 347278 136170 347334 136226
rect 347402 136170 347458 136226
rect 347526 136170 347582 136226
rect 347154 136046 347210 136102
rect 347278 136046 347334 136102
rect 347402 136046 347458 136102
rect 347526 136046 347582 136102
rect 347154 135922 347210 135978
rect 347278 135922 347334 135978
rect 347402 135922 347458 135978
rect 347526 135922 347582 135978
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 347154 118294 347210 118350
rect 347278 118294 347334 118350
rect 347402 118294 347458 118350
rect 347526 118294 347582 118350
rect 347154 118170 347210 118226
rect 347278 118170 347334 118226
rect 347402 118170 347458 118226
rect 347526 118170 347582 118226
rect 347154 118046 347210 118102
rect 347278 118046 347334 118102
rect 347402 118046 347458 118102
rect 347526 118046 347582 118102
rect 347154 117922 347210 117978
rect 347278 117922 347334 117978
rect 347402 117922 347458 117978
rect 347526 117922 347582 117978
rect 347154 100294 347210 100350
rect 347278 100294 347334 100350
rect 347402 100294 347458 100350
rect 347526 100294 347582 100350
rect 347154 100170 347210 100226
rect 347278 100170 347334 100226
rect 347402 100170 347458 100226
rect 347526 100170 347582 100226
rect 347154 100046 347210 100102
rect 347278 100046 347334 100102
rect 347402 100046 347458 100102
rect 347526 100046 347582 100102
rect 347154 99922 347210 99978
rect 347278 99922 347334 99978
rect 347402 99922 347458 99978
rect 347526 99922 347582 99978
rect 367052 135422 367108 135478
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 374154 112294 374210 112350
rect 374278 112294 374334 112350
rect 374402 112294 374458 112350
rect 374526 112294 374582 112350
rect 374154 112170 374210 112226
rect 374278 112170 374334 112226
rect 374402 112170 374458 112226
rect 374526 112170 374582 112226
rect 374154 112046 374210 112102
rect 374278 112046 374334 112102
rect 374402 112046 374458 112102
rect 374526 112046 374582 112102
rect 374154 111922 374210 111978
rect 374278 111922 374334 111978
rect 374402 111922 374458 111978
rect 374526 111922 374582 111978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 404874 148294 404930 148350
rect 404998 148294 405054 148350
rect 405122 148294 405178 148350
rect 405246 148294 405302 148350
rect 404874 148170 404930 148226
rect 404998 148170 405054 148226
rect 405122 148170 405178 148226
rect 405246 148170 405302 148226
rect 404874 148046 404930 148102
rect 404998 148046 405054 148102
rect 405122 148046 405178 148102
rect 405246 148046 405302 148102
rect 404874 147922 404930 147978
rect 404998 147922 405054 147978
rect 405122 147922 405178 147978
rect 405246 147922 405302 147978
rect 404874 130294 404930 130350
rect 404998 130294 405054 130350
rect 405122 130294 405178 130350
rect 405246 130294 405302 130350
rect 404874 130170 404930 130226
rect 404998 130170 405054 130226
rect 405122 130170 405178 130226
rect 405246 130170 405302 130226
rect 404874 130046 404930 130102
rect 404998 130046 405054 130102
rect 405122 130046 405178 130102
rect 405246 130046 405302 130102
rect 404874 129922 404930 129978
rect 404998 129922 405054 129978
rect 405122 129922 405178 129978
rect 405246 129922 405302 129978
rect 404874 112294 404930 112350
rect 404998 112294 405054 112350
rect 405122 112294 405178 112350
rect 405246 112294 405302 112350
rect 404874 112170 404930 112226
rect 404998 112170 405054 112226
rect 405122 112170 405178 112226
rect 405246 112170 405302 112226
rect 404874 112046 404930 112102
rect 404998 112046 405054 112102
rect 405122 112046 405178 112102
rect 405246 112046 405302 112102
rect 404874 111922 404930 111978
rect 404998 111922 405054 111978
rect 405122 111922 405178 111978
rect 405246 111922 405302 111978
rect 403228 103922 403284 103978
rect 377874 100294 377930 100350
rect 377998 100294 378054 100350
rect 378122 100294 378178 100350
rect 378246 100294 378302 100350
rect 377874 100170 377930 100226
rect 377998 100170 378054 100226
rect 378122 100170 378178 100226
rect 378246 100170 378302 100226
rect 377874 100046 377930 100102
rect 377998 100046 378054 100102
rect 378122 100046 378178 100102
rect 378246 100046 378302 100102
rect 377874 99922 377930 99978
rect 377998 99922 378054 99978
rect 378122 99922 378178 99978
rect 378246 99922 378302 99978
rect 408594 154294 408650 154350
rect 408718 154294 408774 154350
rect 408842 154294 408898 154350
rect 408966 154294 409022 154350
rect 408594 154170 408650 154226
rect 408718 154170 408774 154226
rect 408842 154170 408898 154226
rect 408966 154170 409022 154226
rect 408594 154046 408650 154102
rect 408718 154046 408774 154102
rect 408842 154046 408898 154102
rect 408966 154046 409022 154102
rect 408594 153922 408650 153978
rect 408718 153922 408774 153978
rect 408842 153922 408898 153978
rect 408966 153922 409022 153978
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 423276 122462 423332 122518
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 406700 104102 406756 104158
rect 413308 115262 413364 115318
rect 414988 115082 415044 115138
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 408594 100294 408650 100350
rect 408718 100294 408774 100350
rect 408842 100294 408898 100350
rect 408966 100294 409022 100350
rect 408594 100170 408650 100226
rect 408718 100170 408774 100226
rect 408842 100170 408898 100226
rect 408966 100170 409022 100226
rect 408594 100046 408650 100102
rect 408718 100046 408774 100102
rect 408842 100046 408898 100102
rect 408966 100046 409022 100102
rect 408594 99922 408650 99978
rect 408718 99922 408774 99978
rect 408842 99922 408898 99978
rect 408966 99922 409022 99978
rect 374518 94294 374574 94350
rect 374642 94294 374698 94350
rect 374518 94170 374574 94226
rect 374642 94170 374698 94226
rect 374518 94046 374574 94102
rect 374642 94046 374698 94102
rect 374518 93922 374574 93978
rect 374642 93922 374698 93978
rect 405238 94294 405294 94350
rect 405362 94294 405418 94350
rect 405238 94170 405294 94226
rect 405362 94170 405418 94226
rect 405238 94046 405294 94102
rect 405362 94046 405418 94102
rect 405238 93922 405294 93978
rect 405362 93922 405418 93978
rect 347154 82294 347210 82350
rect 347278 82294 347334 82350
rect 347402 82294 347458 82350
rect 347526 82294 347582 82350
rect 347154 82170 347210 82226
rect 347278 82170 347334 82226
rect 347402 82170 347458 82226
rect 347526 82170 347582 82226
rect 347154 82046 347210 82102
rect 347278 82046 347334 82102
rect 347402 82046 347458 82102
rect 347526 82046 347582 82102
rect 347154 81922 347210 81978
rect 347278 81922 347334 81978
rect 347402 81922 347458 81978
rect 347526 81922 347582 81978
rect 389878 82294 389934 82350
rect 390002 82294 390058 82350
rect 389878 82170 389934 82226
rect 390002 82170 390058 82226
rect 389878 82046 389934 82102
rect 390002 82046 390058 82102
rect 389878 81922 389934 81978
rect 390002 81922 390058 81978
rect 374518 76294 374574 76350
rect 374642 76294 374698 76350
rect 374518 76170 374574 76226
rect 374642 76170 374698 76226
rect 374518 76046 374574 76102
rect 374642 76046 374698 76102
rect 374518 75922 374574 75978
rect 374642 75922 374698 75978
rect 405238 76294 405294 76350
rect 405362 76294 405418 76350
rect 405238 76170 405294 76226
rect 405362 76170 405418 76226
rect 405238 76046 405294 76102
rect 405362 76046 405418 76102
rect 405238 75922 405294 75978
rect 405362 75922 405418 75978
rect 347154 64294 347210 64350
rect 347278 64294 347334 64350
rect 347402 64294 347458 64350
rect 347526 64294 347582 64350
rect 347154 64170 347210 64226
rect 347278 64170 347334 64226
rect 347402 64170 347458 64226
rect 347526 64170 347582 64226
rect 347154 64046 347210 64102
rect 347278 64046 347334 64102
rect 347402 64046 347458 64102
rect 347526 64046 347582 64102
rect 347154 63922 347210 63978
rect 347278 63922 347334 63978
rect 347402 63922 347458 63978
rect 347526 63922 347582 63978
rect 389878 64294 389934 64350
rect 390002 64294 390058 64350
rect 389878 64170 389934 64226
rect 390002 64170 390058 64226
rect 389878 64046 389934 64102
rect 390002 64046 390058 64102
rect 389878 63922 389934 63978
rect 390002 63922 390058 63978
rect 374518 58294 374574 58350
rect 374642 58294 374698 58350
rect 374518 58170 374574 58226
rect 374642 58170 374698 58226
rect 374518 58046 374574 58102
rect 374642 58046 374698 58102
rect 374518 57922 374574 57978
rect 374642 57922 374698 57978
rect 405238 58294 405294 58350
rect 405362 58294 405418 58350
rect 405238 58170 405294 58226
rect 405362 58170 405418 58226
rect 405238 58046 405294 58102
rect 405362 58046 405418 58102
rect 405238 57922 405294 57978
rect 405362 57922 405418 57978
rect 347154 46294 347210 46350
rect 347278 46294 347334 46350
rect 347402 46294 347458 46350
rect 347526 46294 347582 46350
rect 347154 46170 347210 46226
rect 347278 46170 347334 46226
rect 347402 46170 347458 46226
rect 347526 46170 347582 46226
rect 347154 46046 347210 46102
rect 347278 46046 347334 46102
rect 347402 46046 347458 46102
rect 347526 46046 347582 46102
rect 347154 45922 347210 45978
rect 347278 45922 347334 45978
rect 347402 45922 347458 45978
rect 347526 45922 347582 45978
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 408594 46294 408650 46350
rect 408718 46294 408774 46350
rect 408842 46294 408898 46350
rect 408966 46294 409022 46350
rect 408594 46170 408650 46226
rect 408718 46170 408774 46226
rect 408842 46170 408898 46226
rect 408966 46170 409022 46226
rect 408594 46046 408650 46102
rect 408718 46046 408774 46102
rect 408842 46046 408898 46102
rect 408966 46046 409022 46102
rect 408594 45922 408650 45978
rect 408718 45922 408774 45978
rect 408842 45922 408898 45978
rect 408966 45922 409022 45978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 408594 28294 408650 28350
rect 408718 28294 408774 28350
rect 408842 28294 408898 28350
rect 408966 28294 409022 28350
rect 408594 28170 408650 28226
rect 408718 28170 408774 28226
rect 408842 28170 408898 28226
rect 408966 28170 409022 28226
rect 408594 28046 408650 28102
rect 408718 28046 408774 28102
rect 408842 28046 408898 28102
rect 408966 28046 409022 28102
rect 408594 27922 408650 27978
rect 408718 27922 408774 27978
rect 408842 27922 408898 27978
rect 408966 27922 409022 27978
rect 408594 10294 408650 10350
rect 408718 10294 408774 10350
rect 408842 10294 408898 10350
rect 408966 10294 409022 10350
rect 408594 10170 408650 10226
rect 408718 10170 408774 10226
rect 408842 10170 408898 10226
rect 408966 10170 409022 10226
rect 408594 10046 408650 10102
rect 408718 10046 408774 10102
rect 408842 10046 408898 10102
rect 408966 10046 409022 10102
rect 408594 9922 408650 9978
rect 408718 9922 408774 9978
rect 408842 9922 408898 9978
rect 408966 9922 409022 9978
rect 408594 -1176 408650 -1120
rect 408718 -1176 408774 -1120
rect 408842 -1176 408898 -1120
rect 408966 -1176 409022 -1120
rect 408594 -1300 408650 -1244
rect 408718 -1300 408774 -1244
rect 408842 -1300 408898 -1244
rect 408966 -1300 409022 -1244
rect 408594 -1424 408650 -1368
rect 408718 -1424 408774 -1368
rect 408842 -1424 408898 -1368
rect 408966 -1424 409022 -1368
rect 408594 -1548 408650 -1492
rect 408718 -1548 408774 -1492
rect 408842 -1548 408898 -1492
rect 408966 -1548 409022 -1492
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 576268 158642 576324 158698
rect 558460 157612 558516 157618
rect 558460 157562 558516 157612
rect 514108 157382 514164 157438
rect 574812 155582 574868 155638
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 457996 149642 458052 149698
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 463148 144602 463204 144658
rect 462924 137402 462980 137458
rect 463148 135602 463204 135658
rect 463260 141182 463316 141238
rect 465388 139742 465444 139798
rect 465388 135242 465444 135298
rect 465500 139562 465556 139618
rect 463260 134342 463316 134398
rect 463036 132542 463092 132598
rect 462812 132362 462868 132418
rect 465500 132182 465556 132238
rect 464518 130294 464574 130350
rect 464642 130294 464698 130350
rect 464518 130170 464574 130226
rect 464642 130170 464698 130226
rect 464518 130046 464574 130102
rect 464642 130046 464698 130102
rect 464518 129922 464574 129978
rect 464642 129922 464698 129978
rect 466732 144782 466788 144838
rect 466396 135422 466452 135478
rect 490028 144782 490084 144838
rect 497868 144602 497924 144658
rect 505708 144422 505764 144478
rect 513548 143882 513604 143938
rect 507276 143702 507332 143758
rect 508844 143522 508900 143578
rect 511980 142828 512036 142858
rect 511980 142802 512036 142828
rect 472892 142622 472948 142678
rect 468636 142442 468692 142498
rect 480620 139748 480676 139798
rect 480620 139742 480676 139748
rect 482188 139580 482244 139618
rect 482188 139562 482244 139580
rect 466732 137582 466788 137638
rect 574252 138482 574308 138538
rect 479878 136294 479934 136350
rect 480002 136294 480058 136350
rect 479878 136170 479934 136226
rect 480002 136170 480058 136226
rect 479878 136046 479934 136102
rect 480002 136046 480058 136102
rect 479878 135922 479934 135978
rect 480002 135922 480058 135978
rect 510598 136294 510654 136350
rect 510722 136294 510778 136350
rect 510598 136170 510654 136226
rect 510722 136170 510778 136226
rect 510598 136046 510654 136102
rect 510722 136046 510778 136102
rect 510598 135922 510654 135978
rect 510722 135922 510778 135978
rect 541318 136294 541374 136350
rect 541442 136294 541498 136350
rect 541318 136170 541374 136226
rect 541442 136170 541498 136226
rect 541318 136046 541374 136102
rect 541442 136046 541498 136102
rect 541318 135922 541374 135978
rect 541442 135922 541498 135978
rect 572038 136294 572094 136350
rect 572162 136294 572218 136350
rect 572038 136170 572094 136226
rect 572162 136170 572218 136226
rect 572038 136046 572094 136102
rect 572162 136046 572218 136102
rect 572038 135922 572094 135978
rect 572162 135922 572218 135978
rect 467068 134162 467124 134218
rect 466620 133982 466676 134038
rect 495238 130294 495294 130350
rect 495362 130294 495418 130350
rect 495238 130170 495294 130226
rect 495362 130170 495418 130226
rect 495238 130046 495294 130102
rect 495362 130046 495418 130102
rect 495238 129922 495294 129978
rect 495362 129922 495418 129978
rect 525958 130294 526014 130350
rect 526082 130294 526138 130350
rect 525958 130170 526014 130226
rect 526082 130170 526138 130226
rect 525958 130046 526014 130102
rect 526082 130046 526138 130102
rect 525958 129922 526014 129978
rect 526082 129922 526138 129978
rect 556678 130294 556734 130350
rect 556802 130294 556858 130350
rect 556678 130170 556734 130226
rect 556802 130170 556858 130226
rect 556678 130046 556734 130102
rect 556802 130046 556858 130102
rect 556678 129922 556734 129978
rect 556802 129922 556858 129978
rect 466284 127502 466340 127558
rect 466172 122462 466228 122518
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 479878 118294 479934 118350
rect 480002 118294 480058 118350
rect 479878 118170 479934 118226
rect 480002 118170 480058 118226
rect 479878 118046 479934 118102
rect 480002 118046 480058 118102
rect 479878 117922 479934 117978
rect 480002 117922 480058 117978
rect 510598 118294 510654 118350
rect 510722 118294 510778 118350
rect 510598 118170 510654 118226
rect 510722 118170 510778 118226
rect 510598 118046 510654 118102
rect 510722 118046 510778 118102
rect 510598 117922 510654 117978
rect 510722 117922 510778 117978
rect 541318 118294 541374 118350
rect 541442 118294 541498 118350
rect 541318 118170 541374 118226
rect 541442 118170 541498 118226
rect 541318 118046 541374 118102
rect 541442 118046 541498 118102
rect 541318 117922 541374 117978
rect 541442 117922 541498 117978
rect 572038 118294 572094 118350
rect 572162 118294 572218 118350
rect 572038 118170 572094 118226
rect 572162 118170 572218 118226
rect 572038 118046 572094 118102
rect 572162 118046 572218 118102
rect 572038 117922 572094 117978
rect 572162 117922 572218 117978
rect 574140 113822 574196 113878
rect 464518 112294 464574 112350
rect 464642 112294 464698 112350
rect 464518 112170 464574 112226
rect 464642 112170 464698 112226
rect 464518 112046 464574 112102
rect 464642 112046 464698 112102
rect 464518 111922 464574 111978
rect 464642 111922 464698 111978
rect 495238 112294 495294 112350
rect 495362 112294 495418 112350
rect 495238 112170 495294 112226
rect 495362 112170 495418 112226
rect 495238 112046 495294 112102
rect 495362 112046 495418 112102
rect 495238 111922 495294 111978
rect 495362 111922 495418 111978
rect 525958 112294 526014 112350
rect 526082 112294 526138 112350
rect 525958 112170 526014 112226
rect 526082 112170 526138 112226
rect 525958 112046 526014 112102
rect 526082 112046 526138 112102
rect 525958 111922 526014 111978
rect 526082 111922 526138 111978
rect 556678 112294 556734 112350
rect 556802 112294 556858 112350
rect 556678 112170 556734 112226
rect 556802 112170 556858 112226
rect 556678 112046 556734 112102
rect 556802 112046 556858 112102
rect 556678 111922 556734 111978
rect 556802 111922 556858 111978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 479878 100294 479934 100350
rect 480002 100294 480058 100350
rect 479878 100170 479934 100226
rect 480002 100170 480058 100226
rect 479878 100046 479934 100102
rect 480002 100046 480058 100102
rect 479878 99922 479934 99978
rect 480002 99922 480058 99978
rect 510598 100294 510654 100350
rect 510722 100294 510778 100350
rect 510598 100170 510654 100226
rect 510722 100170 510778 100226
rect 510598 100046 510654 100102
rect 510722 100046 510778 100102
rect 510598 99922 510654 99978
rect 510722 99922 510778 99978
rect 541318 100294 541374 100350
rect 541442 100294 541498 100350
rect 541318 100170 541374 100226
rect 541442 100170 541498 100226
rect 541318 100046 541374 100102
rect 541442 100046 541498 100102
rect 541318 99922 541374 99978
rect 541442 99922 541498 99978
rect 572038 100294 572094 100350
rect 572162 100294 572218 100350
rect 572038 100170 572094 100226
rect 572162 100170 572218 100226
rect 572038 100046 572094 100102
rect 572162 100046 572218 100102
rect 572038 99922 572094 99978
rect 572162 99922 572218 99978
rect 464518 94294 464574 94350
rect 464642 94294 464698 94350
rect 464518 94170 464574 94226
rect 464642 94170 464698 94226
rect 464518 94046 464574 94102
rect 464642 94046 464698 94102
rect 464518 93922 464574 93978
rect 464642 93922 464698 93978
rect 495238 94294 495294 94350
rect 495362 94294 495418 94350
rect 495238 94170 495294 94226
rect 495362 94170 495418 94226
rect 495238 94046 495294 94102
rect 495362 94046 495418 94102
rect 495238 93922 495294 93978
rect 495362 93922 495418 93978
rect 525958 94294 526014 94350
rect 526082 94294 526138 94350
rect 525958 94170 526014 94226
rect 526082 94170 526138 94226
rect 525958 94046 526014 94102
rect 526082 94046 526138 94102
rect 525958 93922 526014 93978
rect 526082 93922 526138 93978
rect 556678 94294 556734 94350
rect 556802 94294 556858 94350
rect 556678 94170 556734 94226
rect 556802 94170 556858 94226
rect 556678 94046 556734 94102
rect 556802 94046 556858 94102
rect 556678 93922 556734 93978
rect 556802 93922 556858 93978
rect 479878 82294 479934 82350
rect 480002 82294 480058 82350
rect 479878 82170 479934 82226
rect 480002 82170 480058 82226
rect 479878 82046 479934 82102
rect 480002 82046 480058 82102
rect 479878 81922 479934 81978
rect 480002 81922 480058 81978
rect 510598 82294 510654 82350
rect 510722 82294 510778 82350
rect 510598 82170 510654 82226
rect 510722 82170 510778 82226
rect 510598 82046 510654 82102
rect 510722 82046 510778 82102
rect 510598 81922 510654 81978
rect 510722 81922 510778 81978
rect 541318 82294 541374 82350
rect 541442 82294 541498 82350
rect 541318 82170 541374 82226
rect 541442 82170 541498 82226
rect 541318 82046 541374 82102
rect 541442 82046 541498 82102
rect 541318 81922 541374 81978
rect 541442 81922 541498 81978
rect 572038 82294 572094 82350
rect 572162 82294 572218 82350
rect 572038 82170 572094 82226
rect 572162 82170 572218 82226
rect 572038 82046 572094 82102
rect 572162 82046 572218 82102
rect 572038 81922 572094 81978
rect 572162 81922 572218 81978
rect 464518 76294 464574 76350
rect 464642 76294 464698 76350
rect 464518 76170 464574 76226
rect 464642 76170 464698 76226
rect 464518 76046 464574 76102
rect 464642 76046 464698 76102
rect 464518 75922 464574 75978
rect 464642 75922 464698 75978
rect 495238 76294 495294 76350
rect 495362 76294 495418 76350
rect 495238 76170 495294 76226
rect 495362 76170 495418 76226
rect 495238 76046 495294 76102
rect 495362 76046 495418 76102
rect 495238 75922 495294 75978
rect 495362 75922 495418 75978
rect 525958 76294 526014 76350
rect 526082 76294 526138 76350
rect 525958 76170 526014 76226
rect 526082 76170 526138 76226
rect 525958 76046 526014 76102
rect 526082 76046 526138 76102
rect 525958 75922 526014 75978
rect 526082 75922 526138 75978
rect 556678 76294 556734 76350
rect 556802 76294 556858 76350
rect 556678 76170 556734 76226
rect 556802 76170 556858 76226
rect 556678 76046 556734 76102
rect 556802 76046 556858 76102
rect 556678 75922 556734 75978
rect 556802 75922 556858 75978
rect 479878 64294 479934 64350
rect 480002 64294 480058 64350
rect 479878 64170 479934 64226
rect 480002 64170 480058 64226
rect 479878 64046 479934 64102
rect 480002 64046 480058 64102
rect 479878 63922 479934 63978
rect 480002 63922 480058 63978
rect 510598 64294 510654 64350
rect 510722 64294 510778 64350
rect 510598 64170 510654 64226
rect 510722 64170 510778 64226
rect 510598 64046 510654 64102
rect 510722 64046 510778 64102
rect 510598 63922 510654 63978
rect 510722 63922 510778 63978
rect 541318 64294 541374 64350
rect 541442 64294 541498 64350
rect 541318 64170 541374 64226
rect 541442 64170 541498 64226
rect 541318 64046 541374 64102
rect 541442 64046 541498 64102
rect 541318 63922 541374 63978
rect 541442 63922 541498 63978
rect 572038 64294 572094 64350
rect 572162 64294 572218 64350
rect 572038 64170 572094 64226
rect 572162 64170 572218 64226
rect 572038 64046 572094 64102
rect 572162 64046 572218 64102
rect 572038 63922 572094 63978
rect 572162 63922 572218 63978
rect 574588 145322 574644 145378
rect 574924 146942 574980 146998
rect 575148 113876 575204 113878
rect 575148 113822 575204 113876
rect 464518 58294 464574 58350
rect 464642 58294 464698 58350
rect 464518 58170 464574 58226
rect 464642 58170 464698 58226
rect 464518 58046 464574 58102
rect 464642 58046 464698 58102
rect 464518 57922 464574 57978
rect 464642 57922 464698 57978
rect 495238 58294 495294 58350
rect 495362 58294 495418 58350
rect 495238 58170 495294 58226
rect 495362 58170 495418 58226
rect 495238 58046 495294 58102
rect 495362 58046 495418 58102
rect 495238 57922 495294 57978
rect 495362 57922 495418 57978
rect 525958 58294 526014 58350
rect 526082 58294 526138 58350
rect 525958 58170 526014 58226
rect 526082 58170 526138 58226
rect 525958 58046 526014 58102
rect 526082 58046 526138 58102
rect 525958 57922 526014 57978
rect 526082 57922 526138 57978
rect 556678 58294 556734 58350
rect 556802 58294 556858 58350
rect 556678 58170 556734 58226
rect 556802 58170 556858 58226
rect 556678 58046 556734 58102
rect 556802 58046 556858 58102
rect 556678 57922 556734 57978
rect 556802 57922 556858 57978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 479878 46294 479934 46350
rect 480002 46294 480058 46350
rect 479878 46170 479934 46226
rect 480002 46170 480058 46226
rect 479878 46046 479934 46102
rect 480002 46046 480058 46102
rect 479878 45922 479934 45978
rect 480002 45922 480058 45978
rect 510598 46294 510654 46350
rect 510722 46294 510778 46350
rect 510598 46170 510654 46226
rect 510722 46170 510778 46226
rect 510598 46046 510654 46102
rect 510722 46046 510778 46102
rect 510598 45922 510654 45978
rect 510722 45922 510778 45978
rect 541318 46294 541374 46350
rect 541442 46294 541498 46350
rect 541318 46170 541374 46226
rect 541442 46170 541498 46226
rect 541318 46046 541374 46102
rect 541442 46046 541498 46102
rect 541318 45922 541374 45978
rect 541442 45922 541498 45978
rect 572038 46294 572094 46350
rect 572162 46294 572218 46350
rect 572038 46170 572094 46226
rect 572162 46170 572218 46226
rect 572038 46046 572094 46102
rect 572162 46046 572218 46102
rect 572038 45922 572094 45978
rect 572162 45922 572218 45978
rect 578060 155402 578116 155458
rect 576380 149642 576436 149698
rect 577948 141902 578004 141958
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 590492 160982 590548 161038
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 590828 160802 590884 160858
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 591276 161162 591332 161218
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 591052 157742 591108 157798
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 590044 152740 590100 152758
rect 590044 152702 590100 152740
rect 590604 151982 590660 152038
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 578844 140282 578900 140338
rect 590492 150362 590548 150418
rect 590156 139412 590212 139438
rect 590156 139382 590212 139412
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 590716 141182 590772 141238
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 464518 40294 464574 40350
rect 464642 40294 464698 40350
rect 464518 40170 464574 40226
rect 464642 40170 464698 40226
rect 464518 40046 464574 40102
rect 464642 40046 464698 40102
rect 464518 39922 464574 39978
rect 464642 39922 464698 39978
rect 495238 40294 495294 40350
rect 495362 40294 495418 40350
rect 495238 40170 495294 40226
rect 495362 40170 495418 40226
rect 495238 40046 495294 40102
rect 495362 40046 495418 40102
rect 495238 39922 495294 39978
rect 495362 39922 495418 39978
rect 525958 40294 526014 40350
rect 526082 40294 526138 40350
rect 525958 40170 526014 40226
rect 526082 40170 526138 40226
rect 525958 40046 526014 40102
rect 526082 40046 526138 40102
rect 525958 39922 526014 39978
rect 526082 39922 526138 39978
rect 556678 40294 556734 40350
rect 556802 40294 556858 40350
rect 556678 40170 556734 40226
rect 556802 40170 556858 40226
rect 556678 40046 556734 40102
rect 556802 40046 556858 40102
rect 556678 39922 556734 39978
rect 556802 39922 556858 39978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 479878 28294 479934 28350
rect 480002 28294 480058 28350
rect 479878 28170 479934 28226
rect 480002 28170 480058 28226
rect 479878 28046 479934 28102
rect 480002 28046 480058 28102
rect 479878 27922 479934 27978
rect 480002 27922 480058 27978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 510598 28294 510654 28350
rect 510722 28294 510778 28350
rect 510598 28170 510654 28226
rect 510722 28170 510778 28226
rect 510598 28046 510654 28102
rect 510722 28046 510778 28102
rect 510598 27922 510654 27978
rect 510722 27922 510778 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 541318 28294 541374 28350
rect 541442 28294 541498 28350
rect 541318 28170 541374 28226
rect 541442 28170 541498 28226
rect 541318 28046 541374 28102
rect 541442 28046 541498 28102
rect 541318 27922 541374 27978
rect 541442 27922 541498 27978
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 577948 31742 578004 31798
rect 574588 30122 574644 30178
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 572038 28294 572094 28350
rect 572162 28294 572218 28350
rect 572038 28170 572094 28226
rect 572162 28170 572218 28226
rect 572038 28046 572094 28102
rect 572162 28046 572218 28102
rect 572038 27922 572094 27978
rect 572162 27922 572218 27978
rect 578172 33542 578228 33598
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 589932 35162 589988 35218
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580063 159114 580102
rect 98102 580046 130346 580063
rect -1916 580007 130346 580046
rect 130402 580007 130470 580063
rect 130526 580007 130594 580063
rect 130650 580007 130718 580063
rect 130774 580046 159114 580063
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect 130774 580007 597980 580046
rect -1916 579978 597980 580007
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579939 159114 579978
rect 98102 579922 130346 579939
rect -1916 579883 130346 579922
rect 130402 579883 130470 579939
rect 130526 579883 130594 579939
rect 130650 579883 130718 579939
rect 130774 579922 159114 579939
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect 130774 579883 597980 579922
rect -1916 579826 597980 579883
rect 174620 573778 590564 573794
rect 174620 573722 174636 573778
rect 174692 573722 590492 573778
rect 590548 573722 590564 573778
rect 174620 573706 590564 573722
rect 179660 571978 341140 571994
rect 179660 571922 179676 571978
rect 179732 571922 341068 571978
rect 341124 571922 341140 571978
rect 179660 571906 341140 571922
rect 199708 571258 590676 571274
rect 199708 571202 199724 571258
rect 199780 571202 590604 571258
rect 590660 571202 590676 571258
rect 199708 571186 590676 571202
rect 202396 570358 253780 570374
rect 202396 570302 202412 570358
rect 202468 570302 253708 570358
rect 253764 570302 253780 570358
rect 202396 570286 253780 570302
rect 179996 569818 590564 569834
rect 179996 569762 180012 569818
rect 180068 569762 590492 569818
rect 590548 569762 590564 569818
rect 179996 569746 590564 569762
rect 176300 569638 590900 569654
rect 176300 569582 176316 569638
rect 176372 569582 590828 569638
rect 590884 569582 590900 569638
rect 176300 569566 590900 569582
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect 197580 566218 533220 566234
rect 197580 566162 197596 566218
rect 197652 566162 533148 566218
rect 533204 566162 533220 566218
rect 197580 566146 533220 566162
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562272 597980 562294
rect -1916 562226 116228 562272
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562216 116228 562226
rect 116284 562216 116352 562272
rect 116408 562216 116476 562272
rect 116532 562216 116600 562272
rect 116656 562216 116724 562272
rect 116780 562216 116848 562272
rect 116904 562216 116972 562272
rect 117028 562216 117096 562272
rect 117152 562216 117220 562272
rect 117276 562216 117344 562272
rect 117400 562216 117468 562272
rect 117524 562216 117592 562272
rect 117648 562216 117716 562272
rect 117772 562216 117840 562272
rect 117896 562216 117964 562272
rect 118020 562216 118088 562272
rect 118144 562216 118212 562272
rect 118268 562216 118336 562272
rect 118392 562216 118460 562272
rect 118516 562216 118584 562272
rect 118640 562216 118708 562272
rect 118764 562216 118832 562272
rect 118888 562216 118956 562272
rect 119012 562216 119080 562272
rect 119136 562216 119204 562272
rect 119260 562216 119328 562272
rect 119384 562216 119452 562272
rect 119508 562216 119576 562272
rect 119632 562216 119700 562272
rect 119756 562216 119824 562272
rect 119880 562216 119948 562272
rect 120004 562216 120072 562272
rect 120128 562216 120196 562272
rect 120252 562216 120320 562272
rect 120376 562216 120444 562272
rect 120500 562216 120568 562272
rect 120624 562216 120692 562272
rect 120748 562216 120816 562272
rect 120872 562216 120940 562272
rect 120996 562216 121064 562272
rect 121120 562216 121188 562272
rect 121244 562216 121312 562272
rect 121368 562216 121436 562272
rect 121492 562216 121560 562272
rect 121616 562216 121684 562272
rect 121740 562216 121808 562272
rect 121864 562216 121932 562272
rect 121988 562216 122056 562272
rect 122112 562216 122180 562272
rect 122236 562216 122304 562272
rect 122360 562216 122428 562272
rect 122484 562216 122552 562272
rect 122608 562216 122676 562272
rect 122732 562216 122800 562272
rect 122856 562216 122924 562272
rect 122980 562216 123048 562272
rect 123104 562216 123172 562272
rect 123228 562216 123296 562272
rect 123352 562216 123420 562272
rect 123476 562216 123544 562272
rect 123600 562216 123668 562272
rect 123724 562216 123792 562272
rect 123848 562216 123916 562272
rect 123972 562216 124040 562272
rect 124096 562216 124164 562272
rect 124220 562216 124288 562272
rect 124344 562216 124412 562272
rect 124468 562216 124536 562272
rect 124592 562216 124660 562272
rect 124716 562216 124784 562272
rect 124840 562216 124908 562272
rect 124964 562216 125032 562272
rect 125088 562216 125156 562272
rect 125212 562216 125280 562272
rect 125336 562216 125404 562272
rect 125460 562216 125528 562272
rect 125584 562216 125652 562272
rect 125708 562216 125776 562272
rect 125832 562216 125900 562272
rect 125956 562216 126024 562272
rect 126080 562216 126148 562272
rect 126204 562216 126272 562272
rect 126328 562216 126396 562272
rect 126452 562216 126520 562272
rect 126576 562216 126644 562272
rect 126700 562216 126768 562272
rect 126824 562216 126892 562272
rect 126948 562216 127016 562272
rect 127072 562216 127140 562272
rect 127196 562216 127264 562272
rect 127320 562216 127388 562272
rect 127444 562216 127512 562272
rect 127568 562216 127636 562272
rect 127692 562216 127760 562272
rect 127816 562216 127884 562272
rect 127940 562216 128008 562272
rect 128064 562216 128132 562272
rect 128188 562216 128256 562272
rect 128312 562216 128380 562272
rect 128436 562216 128504 562272
rect 128560 562216 128628 562272
rect 128684 562216 128752 562272
rect 128808 562216 128876 562272
rect 128932 562216 129000 562272
rect 129056 562216 129124 562272
rect 129180 562216 129248 562272
rect 129304 562216 129372 562272
rect 129428 562216 129496 562272
rect 129552 562216 129620 562272
rect 129676 562216 129744 562272
rect 129800 562216 129868 562272
rect 129924 562216 129992 562272
rect 130048 562216 130116 562272
rect 130172 562216 130240 562272
rect 130296 562216 130364 562272
rect 130420 562216 130488 562272
rect 130544 562216 130612 562272
rect 130668 562216 130736 562272
rect 130792 562216 130860 562272
rect 130916 562216 130984 562272
rect 131040 562216 131108 562272
rect 131164 562216 131232 562272
rect 131288 562216 131356 562272
rect 131412 562216 131480 562272
rect 131536 562216 131604 562272
rect 131660 562216 131728 562272
rect 131784 562216 131852 562272
rect 131908 562216 131976 562272
rect 132032 562216 132100 562272
rect 132156 562216 132224 562272
rect 132280 562216 132348 562272
rect 132404 562216 132472 562272
rect 132528 562216 132596 562272
rect 132652 562226 597980 562272
rect 132652 562216 159114 562226
rect 98102 562170 159114 562216
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562148 597980 562170
rect -1916 562102 116228 562148
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562092 116228 562102
rect 116284 562092 116352 562148
rect 116408 562092 116476 562148
rect 116532 562092 116600 562148
rect 116656 562092 116724 562148
rect 116780 562092 116848 562148
rect 116904 562092 116972 562148
rect 117028 562092 117096 562148
rect 117152 562092 117220 562148
rect 117276 562092 117344 562148
rect 117400 562092 117468 562148
rect 117524 562092 117592 562148
rect 117648 562092 117716 562148
rect 117772 562092 117840 562148
rect 117896 562092 117964 562148
rect 118020 562092 118088 562148
rect 118144 562092 118212 562148
rect 118268 562092 118336 562148
rect 118392 562092 118460 562148
rect 118516 562092 118584 562148
rect 118640 562092 118708 562148
rect 118764 562092 118832 562148
rect 118888 562092 118956 562148
rect 119012 562092 119080 562148
rect 119136 562092 119204 562148
rect 119260 562092 119328 562148
rect 119384 562092 119452 562148
rect 119508 562092 119576 562148
rect 119632 562092 119700 562148
rect 119756 562092 119824 562148
rect 119880 562092 119948 562148
rect 120004 562092 120072 562148
rect 120128 562092 120196 562148
rect 120252 562092 120320 562148
rect 120376 562092 120444 562148
rect 120500 562092 120568 562148
rect 120624 562092 120692 562148
rect 120748 562092 120816 562148
rect 120872 562092 120940 562148
rect 120996 562092 121064 562148
rect 121120 562092 121188 562148
rect 121244 562092 121312 562148
rect 121368 562092 121436 562148
rect 121492 562092 121560 562148
rect 121616 562092 121684 562148
rect 121740 562092 121808 562148
rect 121864 562092 121932 562148
rect 121988 562092 122056 562148
rect 122112 562092 122180 562148
rect 122236 562092 122304 562148
rect 122360 562092 122428 562148
rect 122484 562092 122552 562148
rect 122608 562092 122676 562148
rect 122732 562092 122800 562148
rect 122856 562092 122924 562148
rect 122980 562092 123048 562148
rect 123104 562092 123172 562148
rect 123228 562092 123296 562148
rect 123352 562092 123420 562148
rect 123476 562092 123544 562148
rect 123600 562092 123668 562148
rect 123724 562092 123792 562148
rect 123848 562092 123916 562148
rect 123972 562092 124040 562148
rect 124096 562092 124164 562148
rect 124220 562092 124288 562148
rect 124344 562092 124412 562148
rect 124468 562092 124536 562148
rect 124592 562092 124660 562148
rect 124716 562092 124784 562148
rect 124840 562092 124908 562148
rect 124964 562092 125032 562148
rect 125088 562092 125156 562148
rect 125212 562092 125280 562148
rect 125336 562092 125404 562148
rect 125460 562092 125528 562148
rect 125584 562092 125652 562148
rect 125708 562092 125776 562148
rect 125832 562092 125900 562148
rect 125956 562092 126024 562148
rect 126080 562092 126148 562148
rect 126204 562092 126272 562148
rect 126328 562092 126396 562148
rect 126452 562092 126520 562148
rect 126576 562092 126644 562148
rect 126700 562092 126768 562148
rect 126824 562092 126892 562148
rect 126948 562092 127016 562148
rect 127072 562092 127140 562148
rect 127196 562092 127264 562148
rect 127320 562092 127388 562148
rect 127444 562092 127512 562148
rect 127568 562092 127636 562148
rect 127692 562092 127760 562148
rect 127816 562092 127884 562148
rect 127940 562092 128008 562148
rect 128064 562092 128132 562148
rect 128188 562092 128256 562148
rect 128312 562092 128380 562148
rect 128436 562092 128504 562148
rect 128560 562092 128628 562148
rect 128684 562092 128752 562148
rect 128808 562092 128876 562148
rect 128932 562092 129000 562148
rect 129056 562092 129124 562148
rect 129180 562092 129248 562148
rect 129304 562092 129372 562148
rect 129428 562092 129496 562148
rect 129552 562092 129620 562148
rect 129676 562092 129744 562148
rect 129800 562092 129868 562148
rect 129924 562092 129992 562148
rect 130048 562092 130116 562148
rect 130172 562092 130240 562148
rect 130296 562092 130364 562148
rect 130420 562092 130488 562148
rect 130544 562092 130612 562148
rect 130668 562092 130736 562148
rect 130792 562092 130860 562148
rect 130916 562092 130984 562148
rect 131040 562092 131108 562148
rect 131164 562092 131232 562148
rect 131288 562092 131356 562148
rect 131412 562092 131480 562148
rect 131536 562092 131604 562148
rect 131660 562092 131728 562148
rect 131784 562092 131852 562148
rect 131908 562092 131976 562148
rect 132032 562092 132100 562148
rect 132156 562092 132224 562148
rect 132280 562092 132348 562148
rect 132404 562092 132472 562148
rect 132528 562092 132596 562148
rect 132652 562102 597980 562148
rect 132652 562092 159114 562102
rect 98102 562046 159114 562092
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 562024 597980 562046
rect -1916 561978 116228 562024
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561968 116228 561978
rect 116284 561968 116352 562024
rect 116408 561968 116476 562024
rect 116532 561968 116600 562024
rect 116656 561968 116724 562024
rect 116780 561968 116848 562024
rect 116904 561968 116972 562024
rect 117028 561968 117096 562024
rect 117152 561968 117220 562024
rect 117276 561968 117344 562024
rect 117400 561968 117468 562024
rect 117524 561968 117592 562024
rect 117648 561968 117716 562024
rect 117772 561968 117840 562024
rect 117896 561968 117964 562024
rect 118020 561968 118088 562024
rect 118144 561968 118212 562024
rect 118268 561968 118336 562024
rect 118392 561968 118460 562024
rect 118516 561968 118584 562024
rect 118640 561968 118708 562024
rect 118764 561968 118832 562024
rect 118888 561968 118956 562024
rect 119012 561968 119080 562024
rect 119136 561968 119204 562024
rect 119260 561968 119328 562024
rect 119384 561968 119452 562024
rect 119508 561968 119576 562024
rect 119632 561968 119700 562024
rect 119756 561968 119824 562024
rect 119880 561968 119948 562024
rect 120004 561968 120072 562024
rect 120128 561968 120196 562024
rect 120252 561968 120320 562024
rect 120376 561968 120444 562024
rect 120500 561968 120568 562024
rect 120624 561968 120692 562024
rect 120748 561968 120816 562024
rect 120872 561968 120940 562024
rect 120996 561968 121064 562024
rect 121120 561968 121188 562024
rect 121244 561968 121312 562024
rect 121368 561968 121436 562024
rect 121492 561968 121560 562024
rect 121616 561968 121684 562024
rect 121740 561968 121808 562024
rect 121864 561968 121932 562024
rect 121988 561968 122056 562024
rect 122112 561968 122180 562024
rect 122236 561968 122304 562024
rect 122360 561968 122428 562024
rect 122484 561968 122552 562024
rect 122608 561968 122676 562024
rect 122732 561968 122800 562024
rect 122856 561968 122924 562024
rect 122980 561968 123048 562024
rect 123104 561968 123172 562024
rect 123228 561968 123296 562024
rect 123352 561968 123420 562024
rect 123476 561968 123544 562024
rect 123600 561968 123668 562024
rect 123724 561968 123792 562024
rect 123848 561968 123916 562024
rect 123972 561968 124040 562024
rect 124096 561968 124164 562024
rect 124220 561968 124288 562024
rect 124344 561968 124412 562024
rect 124468 561968 124536 562024
rect 124592 561968 124660 562024
rect 124716 561968 124784 562024
rect 124840 561968 124908 562024
rect 124964 561968 125032 562024
rect 125088 561968 125156 562024
rect 125212 561968 125280 562024
rect 125336 561968 125404 562024
rect 125460 561968 125528 562024
rect 125584 561968 125652 562024
rect 125708 561968 125776 562024
rect 125832 561968 125900 562024
rect 125956 561968 126024 562024
rect 126080 561968 126148 562024
rect 126204 561968 126272 562024
rect 126328 561968 126396 562024
rect 126452 561968 126520 562024
rect 126576 561968 126644 562024
rect 126700 561968 126768 562024
rect 126824 561968 126892 562024
rect 126948 561968 127016 562024
rect 127072 561968 127140 562024
rect 127196 561968 127264 562024
rect 127320 561968 127388 562024
rect 127444 561968 127512 562024
rect 127568 561968 127636 562024
rect 127692 561968 127760 562024
rect 127816 561968 127884 562024
rect 127940 561968 128008 562024
rect 128064 561968 128132 562024
rect 128188 561968 128256 562024
rect 128312 561968 128380 562024
rect 128436 561968 128504 562024
rect 128560 561968 128628 562024
rect 128684 561968 128752 562024
rect 128808 561968 128876 562024
rect 128932 561968 129000 562024
rect 129056 561968 129124 562024
rect 129180 561968 129248 562024
rect 129304 561968 129372 562024
rect 129428 561968 129496 562024
rect 129552 561968 129620 562024
rect 129676 561968 129744 562024
rect 129800 561968 129868 562024
rect 129924 561968 129992 562024
rect 130048 561968 130116 562024
rect 130172 561968 130240 562024
rect 130296 561968 130364 562024
rect 130420 561968 130488 562024
rect 130544 561968 130612 562024
rect 130668 561968 130736 562024
rect 130792 561968 130860 562024
rect 130916 561968 130984 562024
rect 131040 561968 131108 562024
rect 131164 561968 131232 562024
rect 131288 561968 131356 562024
rect 131412 561968 131480 562024
rect 131536 561968 131604 562024
rect 131660 561968 131728 562024
rect 131784 561968 131852 562024
rect 131908 561968 131976 562024
rect 132032 561968 132100 562024
rect 132156 561968 132224 562024
rect 132280 561968 132348 562024
rect 132404 561968 132472 562024
rect 132528 561968 132596 562024
rect 132652 561978 597980 562024
rect 132652 561968 159114 561978
rect 98102 561922 159114 561968
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544058 159114 544102
rect 67382 544046 104348 544058
rect -1916 544002 104348 544046
rect 104404 544002 104472 544058
rect 104528 544002 104596 544058
rect 104652 544002 104720 544058
rect 104776 544002 104844 544058
rect 104900 544002 104968 544058
rect 105024 544002 105092 544058
rect 105148 544002 105216 544058
rect 105272 544002 105340 544058
rect 105396 544002 105464 544058
rect 105520 544002 105588 544058
rect 105644 544002 105712 544058
rect 105768 544002 105836 544058
rect 105892 544002 105960 544058
rect 106016 544002 106084 544058
rect 106140 544002 106208 544058
rect 106264 544002 106332 544058
rect 106388 544002 106456 544058
rect 106512 544002 106580 544058
rect 106636 544002 106704 544058
rect 106760 544002 106828 544058
rect 106884 544002 106952 544058
rect 107008 544002 107076 544058
rect 107132 544002 107200 544058
rect 107256 544002 107324 544058
rect 107380 544002 107448 544058
rect 107504 544002 107572 544058
rect 107628 544002 107696 544058
rect 107752 544002 107820 544058
rect 107876 544002 107944 544058
rect 108000 544002 108068 544058
rect 108124 544002 108192 544058
rect 108248 544002 108316 544058
rect 108372 544002 108440 544058
rect 108496 544002 108564 544058
rect 108620 544002 108688 544058
rect 108744 544002 108812 544058
rect 108868 544002 108936 544058
rect 108992 544002 109060 544058
rect 109116 544002 109184 544058
rect 109240 544002 109308 544058
rect 109364 544002 109432 544058
rect 109488 544002 109556 544058
rect 109612 544002 109680 544058
rect 109736 544002 109804 544058
rect 109860 544002 109928 544058
rect 109984 544002 110052 544058
rect 110108 544002 110176 544058
rect 110232 544002 110300 544058
rect 110356 544002 110424 544058
rect 110480 544002 110548 544058
rect 110604 544002 110672 544058
rect 110728 544002 110796 544058
rect 110852 544002 110920 544058
rect 110976 544002 111044 544058
rect 111100 544002 111168 544058
rect 111224 544002 111292 544058
rect 111348 544002 111416 544058
rect 111472 544002 111540 544058
rect 111596 544002 111664 544058
rect 111720 544002 111788 544058
rect 111844 544002 111912 544058
rect 111968 544002 112036 544058
rect 112092 544002 112160 544058
rect 112216 544002 112284 544058
rect 112340 544002 112408 544058
rect 112464 544002 112532 544058
rect 112588 544002 112656 544058
rect 112712 544002 112780 544058
rect 112836 544002 112904 544058
rect 112960 544002 113028 544058
rect 113084 544002 113152 544058
rect 113208 544002 113276 544058
rect 113332 544002 113400 544058
rect 113456 544002 113524 544058
rect 113580 544002 113648 544058
rect 113704 544002 113772 544058
rect 113828 544002 113896 544058
rect 113952 544002 114020 544058
rect 114076 544002 114144 544058
rect 114200 544002 114268 544058
rect 114324 544002 114392 544058
rect 114448 544002 114516 544058
rect 114572 544002 114640 544058
rect 114696 544002 114764 544058
rect 114820 544002 114888 544058
rect 114944 544002 115012 544058
rect 115068 544002 115136 544058
rect 115192 544002 115260 544058
rect 115316 544002 115384 544058
rect 115440 544002 115508 544058
rect 115564 544002 115632 544058
rect 115688 544002 115756 544058
rect 115812 544002 115880 544058
rect 115936 544002 116004 544058
rect 116060 544002 116128 544058
rect 116184 544002 116252 544058
rect 116308 544002 116376 544058
rect 116432 544002 116500 544058
rect 116556 544002 116624 544058
rect 116680 544002 116748 544058
rect 116804 544002 116872 544058
rect 116928 544002 116996 544058
rect 117052 544002 117120 544058
rect 117176 544002 117244 544058
rect 117300 544002 117368 544058
rect 117424 544002 117492 544058
rect 117548 544002 117616 544058
rect 117672 544002 117740 544058
rect 117796 544002 117864 544058
rect 117920 544002 117988 544058
rect 118044 544002 118112 544058
rect 118168 544002 118236 544058
rect 118292 544002 118360 544058
rect 118416 544002 118484 544058
rect 118540 544002 118608 544058
rect 118664 544002 118732 544058
rect 118788 544002 118856 544058
rect 118912 544002 118980 544058
rect 119036 544002 119104 544058
rect 119160 544002 119228 544058
rect 119284 544002 119352 544058
rect 119408 544002 119476 544058
rect 119532 544002 119600 544058
rect 119656 544002 119724 544058
rect 119780 544002 119848 544058
rect 119904 544002 119972 544058
rect 120028 544002 120096 544058
rect 120152 544002 120220 544058
rect 120276 544002 120344 544058
rect 120400 544002 120468 544058
rect 120524 544002 120592 544058
rect 120648 544002 120716 544058
rect 120772 544002 120840 544058
rect 120896 544002 120964 544058
rect 121020 544002 121088 544058
rect 121144 544002 121212 544058
rect 121268 544002 121336 544058
rect 121392 544002 121460 544058
rect 121516 544002 121584 544058
rect 121640 544002 121708 544058
rect 121764 544002 121832 544058
rect 121888 544002 121956 544058
rect 122012 544002 122080 544058
rect 122136 544002 122204 544058
rect 122260 544002 122328 544058
rect 122384 544002 122452 544058
rect 122508 544002 122576 544058
rect 122632 544002 122700 544058
rect 122756 544002 122824 544058
rect 122880 544002 122948 544058
rect 123004 544002 123072 544058
rect 123128 544002 123196 544058
rect 123252 544002 123320 544058
rect 123376 544002 123444 544058
rect 123500 544002 123568 544058
rect 123624 544002 123692 544058
rect 123748 544002 123816 544058
rect 123872 544002 123940 544058
rect 123996 544002 124064 544058
rect 124120 544002 124188 544058
rect 124244 544002 124312 544058
rect 124368 544002 124436 544058
rect 124492 544002 124560 544058
rect 124616 544002 124684 544058
rect 124740 544002 124808 544058
rect 124864 544002 124932 544058
rect 124988 544002 125056 544058
rect 125112 544002 125180 544058
rect 125236 544002 125304 544058
rect 125360 544002 125428 544058
rect 125484 544002 125552 544058
rect 125608 544002 125676 544058
rect 125732 544002 125800 544058
rect 125856 544002 125924 544058
rect 125980 544002 126048 544058
rect 126104 544002 126172 544058
rect 126228 544002 126296 544058
rect 126352 544046 159114 544058
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect 126352 544002 597980 544046
rect -1916 543978 597980 544002
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532358 597980 532446
rect -1916 532350 66714 532358
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532302 66714 532350
rect 66770 532302 66838 532358
rect 66894 532302 66962 532358
rect 67018 532302 67086 532358
rect 67142 532302 67210 532358
rect 67266 532302 67334 532358
rect 67390 532302 67458 532358
rect 67514 532302 67582 532358
rect 67638 532302 67706 532358
rect 67762 532302 67830 532358
rect 67886 532302 67954 532358
rect 68010 532302 68078 532358
rect 68134 532302 68202 532358
rect 68258 532302 68326 532358
rect 68382 532302 68450 532358
rect 68506 532302 68574 532358
rect 68630 532302 68698 532358
rect 68754 532302 68822 532358
rect 68878 532302 68946 532358
rect 69002 532302 69070 532358
rect 69126 532302 69194 532358
rect 69250 532302 69318 532358
rect 69374 532302 69442 532358
rect 69498 532302 69566 532358
rect 69622 532302 69690 532358
rect 69746 532302 69814 532358
rect 69870 532302 69938 532358
rect 69994 532302 70062 532358
rect 70118 532302 70186 532358
rect 70242 532302 70310 532358
rect 70366 532302 70434 532358
rect 70490 532302 70558 532358
rect 70614 532302 70682 532358
rect 70738 532302 70806 532358
rect 70862 532302 70930 532358
rect 70986 532302 71054 532358
rect 71110 532302 71178 532358
rect 71234 532302 71302 532358
rect 71358 532302 71426 532358
rect 71482 532302 71550 532358
rect 71606 532302 71674 532358
rect 71730 532302 71798 532358
rect 71854 532302 71922 532358
rect 71978 532302 72046 532358
rect 72102 532302 72170 532358
rect 72226 532302 72294 532358
rect 72350 532302 72418 532358
rect 72474 532302 72542 532358
rect 72598 532302 72666 532358
rect 72722 532302 72790 532358
rect 72846 532302 72914 532358
rect 72970 532302 73038 532358
rect 73094 532302 73162 532358
rect 73218 532302 73286 532358
rect 73342 532302 73410 532358
rect 73466 532302 73534 532358
rect 73590 532302 73658 532358
rect 73714 532302 73782 532358
rect 73838 532302 73906 532358
rect 73962 532302 74030 532358
rect 74086 532302 74154 532358
rect 74210 532302 74278 532358
rect 74334 532302 74402 532358
rect 74458 532302 74526 532358
rect 74582 532302 74650 532358
rect 74706 532350 597980 532358
rect 74706 532302 162834 532350
rect 40382 532294 162834 532302
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531998 597980 532046
rect -1916 531978 66506 531998
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531942 66506 531978
rect 66562 531942 66630 531998
rect 66686 531942 66754 531998
rect 66810 531942 66878 531998
rect 66934 531942 67002 531998
rect 67058 531942 67126 531998
rect 67182 531942 67250 531998
rect 67306 531942 67374 531998
rect 67430 531942 67498 531998
rect 67554 531942 67622 531998
rect 67678 531942 67746 531998
rect 67802 531942 67870 531998
rect 67926 531942 67994 531998
rect 68050 531942 68118 531998
rect 68174 531942 68242 531998
rect 68298 531942 68366 531998
rect 68422 531942 68490 531998
rect 68546 531942 68614 531998
rect 68670 531942 68738 531998
rect 68794 531942 68862 531998
rect 68918 531942 68986 531998
rect 69042 531942 69110 531998
rect 69166 531942 69234 531998
rect 69290 531942 69358 531998
rect 69414 531942 69482 531998
rect 69538 531942 69606 531998
rect 69662 531942 69730 531998
rect 69786 531942 69854 531998
rect 69910 531942 69978 531998
rect 70034 531942 70102 531998
rect 70158 531942 70226 531998
rect 70282 531942 70350 531998
rect 70406 531942 70474 531998
rect 70530 531942 70598 531998
rect 70654 531942 70722 531998
rect 70778 531942 70846 531998
rect 70902 531942 70970 531998
rect 71026 531942 71094 531998
rect 71150 531942 71218 531998
rect 71274 531942 71342 531998
rect 71398 531942 71466 531998
rect 71522 531942 71590 531998
rect 71646 531942 71714 531998
rect 71770 531942 71838 531998
rect 71894 531942 71962 531998
rect 72018 531942 72086 531998
rect 72142 531942 72210 531998
rect 72266 531942 72334 531998
rect 72390 531942 72458 531998
rect 72514 531942 72582 531998
rect 72638 531942 72706 531998
rect 72762 531942 72830 531998
rect 72886 531942 72954 531998
rect 73010 531942 73078 531998
rect 73134 531942 73202 531998
rect 73258 531942 73326 531998
rect 73382 531942 73450 531998
rect 73506 531942 73574 531998
rect 73630 531942 73698 531998
rect 73754 531942 73822 531998
rect 73878 531942 73946 531998
rect 74002 531942 74070 531998
rect 74126 531942 74194 531998
rect 74250 531942 74318 531998
rect 74374 531978 597980 531998
rect 74374 531942 162834 531978
rect 40382 531922 162834 531942
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526058 159114 526102
rect 36662 526046 95846 526058
rect -1916 526002 95846 526046
rect 95902 526002 95970 526058
rect 96026 526002 96094 526058
rect 96150 526002 96218 526058
rect 96274 526002 96342 526058
rect 96398 526002 96466 526058
rect 96522 526002 96590 526058
rect 96646 526002 96714 526058
rect 96770 526002 96838 526058
rect 96894 526002 96962 526058
rect 97018 526002 97086 526058
rect 97142 526002 97210 526058
rect 97266 526002 97334 526058
rect 97390 526002 97458 526058
rect 97514 526002 97582 526058
rect 97638 526002 97706 526058
rect 97762 526002 97830 526058
rect 97886 526002 97954 526058
rect 98010 526002 98078 526058
rect 98134 526002 98202 526058
rect 98258 526002 98326 526058
rect 98382 526002 98450 526058
rect 98506 526002 98574 526058
rect 98630 526002 98698 526058
rect 98754 526002 98822 526058
rect 98878 526002 98946 526058
rect 99002 526002 99070 526058
rect 99126 526002 99194 526058
rect 99250 526002 99318 526058
rect 99374 526002 99442 526058
rect 99498 526002 99566 526058
rect 99622 526002 99690 526058
rect 99746 526002 99814 526058
rect 99870 526002 99938 526058
rect 99994 526002 100062 526058
rect 100118 526002 100186 526058
rect 100242 526002 100310 526058
rect 100366 526002 100434 526058
rect 100490 526002 100558 526058
rect 100614 526002 100682 526058
rect 100738 526002 100806 526058
rect 100862 526002 100930 526058
rect 100986 526002 101054 526058
rect 101110 526002 101178 526058
rect 101234 526002 101302 526058
rect 101358 526002 101426 526058
rect 101482 526002 101550 526058
rect 101606 526002 101674 526058
rect 101730 526002 101798 526058
rect 101854 526002 101922 526058
rect 101978 526002 102046 526058
rect 102102 526002 102170 526058
rect 102226 526002 102294 526058
rect 102350 526002 102418 526058
rect 102474 526002 102542 526058
rect 102598 526002 102666 526058
rect 102722 526002 102790 526058
rect 102846 526002 102914 526058
rect 102970 526002 103038 526058
rect 103094 526002 103162 526058
rect 103218 526002 103286 526058
rect 103342 526002 103410 526058
rect 103466 526002 103534 526058
rect 103590 526002 103658 526058
rect 103714 526002 103782 526058
rect 103838 526002 103906 526058
rect 103962 526002 104030 526058
rect 104086 526002 104154 526058
rect 104210 526002 104278 526058
rect 104334 526002 104402 526058
rect 104458 526002 104526 526058
rect 104582 526002 104650 526058
rect 104706 526002 104774 526058
rect 104830 526002 104898 526058
rect 104954 526002 105022 526058
rect 105078 526002 105146 526058
rect 105202 526002 105270 526058
rect 105326 526002 105394 526058
rect 105450 526002 105518 526058
rect 105574 526002 105642 526058
rect 105698 526002 105766 526058
rect 105822 526002 105890 526058
rect 105946 526002 106014 526058
rect 106070 526002 106138 526058
rect 106194 526002 106262 526058
rect 106318 526002 106386 526058
rect 106442 526002 106510 526058
rect 106566 526002 106634 526058
rect 106690 526002 106758 526058
rect 106814 526002 106882 526058
rect 106938 526002 107006 526058
rect 107062 526002 107130 526058
rect 107186 526002 107254 526058
rect 107310 526002 107378 526058
rect 107434 526002 107502 526058
rect 107558 526002 107626 526058
rect 107682 526002 107750 526058
rect 107806 526002 107874 526058
rect 107930 526002 107998 526058
rect 108054 526002 108122 526058
rect 108178 526002 108246 526058
rect 108302 526002 108370 526058
rect 108426 526002 108494 526058
rect 108550 526002 108618 526058
rect 108674 526002 108742 526058
rect 108798 526002 108866 526058
rect 108922 526002 108990 526058
rect 109046 526002 109114 526058
rect 109170 526002 109238 526058
rect 109294 526002 109362 526058
rect 109418 526002 109486 526058
rect 109542 526002 109610 526058
rect 109666 526002 109734 526058
rect 109790 526002 109858 526058
rect 109914 526002 109982 526058
rect 110038 526002 110106 526058
rect 110162 526002 110230 526058
rect 110286 526002 110354 526058
rect 110410 526002 110478 526058
rect 110534 526002 110602 526058
rect 110658 526002 110726 526058
rect 110782 526002 110850 526058
rect 110906 526002 110974 526058
rect 111030 526002 111098 526058
rect 111154 526002 111222 526058
rect 111278 526002 111346 526058
rect 111402 526002 111470 526058
rect 111526 526002 111594 526058
rect 111650 526002 111718 526058
rect 111774 526002 111842 526058
rect 111898 526002 111966 526058
rect 112022 526002 112090 526058
rect 112146 526002 112214 526058
rect 112270 526002 112338 526058
rect 112394 526002 112462 526058
rect 112518 526002 112586 526058
rect 112642 526002 112710 526058
rect 112766 526002 112834 526058
rect 112890 526002 112958 526058
rect 113014 526002 113082 526058
rect 113138 526002 113206 526058
rect 113262 526002 113330 526058
rect 113386 526002 113454 526058
rect 113510 526002 113578 526058
rect 113634 526002 113702 526058
rect 113758 526002 113826 526058
rect 113882 526002 113950 526058
rect 114006 526002 114074 526058
rect 114130 526002 114198 526058
rect 114254 526002 114322 526058
rect 114378 526002 114446 526058
rect 114502 526002 114570 526058
rect 114626 526002 114694 526058
rect 114750 526002 114818 526058
rect 114874 526046 159114 526058
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect 114874 526002 597980 526046
rect -1916 525978 597980 526002
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514412 597980 514446
rect -1916 514356 60202 514412
rect 60258 514356 60326 514412
rect 60382 514356 60450 514412
rect 60506 514356 60574 514412
rect 60630 514356 60698 514412
rect 60754 514356 60822 514412
rect 60878 514356 60946 514412
rect 61002 514356 61070 514412
rect 61126 514356 61194 514412
rect 61250 514356 61318 514412
rect 61374 514356 61442 514412
rect 61498 514356 61566 514412
rect 61622 514356 61690 514412
rect 61746 514356 61814 514412
rect 61870 514356 61938 514412
rect 61994 514356 62062 514412
rect 62118 514356 62186 514412
rect 62242 514356 62310 514412
rect 62366 514356 62434 514412
rect 62490 514356 62558 514412
rect 62614 514356 62682 514412
rect 62738 514356 62806 514412
rect 62862 514356 62930 514412
rect 62986 514356 63054 514412
rect 63110 514356 63178 514412
rect 63234 514356 63302 514412
rect 63358 514356 63426 514412
rect 63482 514356 63550 514412
rect 63606 514356 63674 514412
rect 63730 514356 63798 514412
rect 63854 514356 63922 514412
rect 63978 514356 64046 514412
rect 64102 514356 64170 514412
rect 64226 514356 64294 514412
rect 64350 514356 64418 514412
rect 64474 514356 64542 514412
rect 64598 514356 64666 514412
rect 64722 514356 64790 514412
rect 64846 514356 64914 514412
rect 64970 514356 65038 514412
rect 65094 514356 65162 514412
rect 65218 514356 65286 514412
rect 65342 514356 65410 514412
rect 65466 514356 65534 514412
rect 65590 514356 65658 514412
rect 65714 514356 65782 514412
rect 65838 514356 65906 514412
rect 65962 514356 66030 514412
rect 66086 514356 66154 514412
rect 66210 514356 66278 514412
rect 66334 514356 66402 514412
rect 66458 514356 597980 514412
rect -1916 514350 597980 514356
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514288 597980 514294
rect -1916 514232 60202 514288
rect 60258 514232 60326 514288
rect 60382 514232 60450 514288
rect 60506 514232 60574 514288
rect 60630 514232 60698 514288
rect 60754 514232 60822 514288
rect 60878 514232 60946 514288
rect 61002 514232 61070 514288
rect 61126 514232 61194 514288
rect 61250 514232 61318 514288
rect 61374 514232 61442 514288
rect 61498 514232 61566 514288
rect 61622 514232 61690 514288
rect 61746 514232 61814 514288
rect 61870 514232 61938 514288
rect 61994 514232 62062 514288
rect 62118 514232 62186 514288
rect 62242 514232 62310 514288
rect 62366 514232 62434 514288
rect 62490 514232 62558 514288
rect 62614 514232 62682 514288
rect 62738 514232 62806 514288
rect 62862 514232 62930 514288
rect 62986 514232 63054 514288
rect 63110 514232 63178 514288
rect 63234 514232 63302 514288
rect 63358 514232 63426 514288
rect 63482 514232 63550 514288
rect 63606 514232 63674 514288
rect 63730 514232 63798 514288
rect 63854 514232 63922 514288
rect 63978 514232 64046 514288
rect 64102 514232 64170 514288
rect 64226 514232 64294 514288
rect 64350 514232 64418 514288
rect 64474 514232 64542 514288
rect 64598 514232 64666 514288
rect 64722 514232 64790 514288
rect 64846 514232 64914 514288
rect 64970 514232 65038 514288
rect 65094 514232 65162 514288
rect 65218 514232 65286 514288
rect 65342 514232 65410 514288
rect 65466 514232 65534 514288
rect 65590 514232 65658 514288
rect 65714 514232 65782 514288
rect 65838 514232 65906 514288
rect 65962 514232 66030 514288
rect 66086 514232 66154 514288
rect 66210 514232 66278 514288
rect 66334 514232 66402 514288
rect 66458 514232 597980 514288
rect -1916 514226 597980 514232
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514164 597980 514170
rect -1916 514108 60202 514164
rect 60258 514108 60326 514164
rect 60382 514108 60450 514164
rect 60506 514108 60574 514164
rect 60630 514108 60698 514164
rect 60754 514108 60822 514164
rect 60878 514108 60946 514164
rect 61002 514108 61070 514164
rect 61126 514108 61194 514164
rect 61250 514108 61318 514164
rect 61374 514108 61442 514164
rect 61498 514108 61566 514164
rect 61622 514108 61690 514164
rect 61746 514108 61814 514164
rect 61870 514108 61938 514164
rect 61994 514108 62062 514164
rect 62118 514108 62186 514164
rect 62242 514108 62310 514164
rect 62366 514108 62434 514164
rect 62490 514108 62558 514164
rect 62614 514108 62682 514164
rect 62738 514108 62806 514164
rect 62862 514108 62930 514164
rect 62986 514108 63054 514164
rect 63110 514108 63178 514164
rect 63234 514108 63302 514164
rect 63358 514108 63426 514164
rect 63482 514108 63550 514164
rect 63606 514108 63674 514164
rect 63730 514108 63798 514164
rect 63854 514108 63922 514164
rect 63978 514108 64046 514164
rect 64102 514108 64170 514164
rect 64226 514108 64294 514164
rect 64350 514108 64418 514164
rect 64474 514108 64542 514164
rect 64598 514108 64666 514164
rect 64722 514108 64790 514164
rect 64846 514108 64914 514164
rect 64970 514108 65038 514164
rect 65094 514108 65162 514164
rect 65218 514108 65286 514164
rect 65342 514108 65410 514164
rect 65466 514108 65534 514164
rect 65590 514108 65658 514164
rect 65714 514108 65782 514164
rect 65838 514108 65906 514164
rect 65962 514108 66030 514164
rect 66086 514108 66154 514164
rect 66210 514108 66278 514164
rect 66334 514108 66402 514164
rect 66458 514108 597980 514164
rect -1916 514102 597980 514108
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 514040 597980 514046
rect -1916 513984 60202 514040
rect 60258 513984 60326 514040
rect 60382 513984 60450 514040
rect 60506 513984 60574 514040
rect 60630 513984 60698 514040
rect 60754 513984 60822 514040
rect 60878 513984 60946 514040
rect 61002 513984 61070 514040
rect 61126 513984 61194 514040
rect 61250 513984 61318 514040
rect 61374 513984 61442 514040
rect 61498 513984 61566 514040
rect 61622 513984 61690 514040
rect 61746 513984 61814 514040
rect 61870 513984 61938 514040
rect 61994 513984 62062 514040
rect 62118 513984 62186 514040
rect 62242 513984 62310 514040
rect 62366 513984 62434 514040
rect 62490 513984 62558 514040
rect 62614 513984 62682 514040
rect 62738 513984 62806 514040
rect 62862 513984 62930 514040
rect 62986 513984 63054 514040
rect 63110 513984 63178 514040
rect 63234 513984 63302 514040
rect 63358 513984 63426 514040
rect 63482 513984 63550 514040
rect 63606 513984 63674 514040
rect 63730 513984 63798 514040
rect 63854 513984 63922 514040
rect 63978 513984 64046 514040
rect 64102 513984 64170 514040
rect 64226 513984 64294 514040
rect 64350 513984 64418 514040
rect 64474 513984 64542 514040
rect 64598 513984 64666 514040
rect 64722 513984 64790 514040
rect 64846 513984 64914 514040
rect 64970 513984 65038 514040
rect 65094 513984 65162 514040
rect 65218 513984 65286 514040
rect 65342 513984 65410 514040
rect 65466 513984 65534 514040
rect 65590 513984 65658 514040
rect 65714 513984 65782 514040
rect 65838 513984 65906 514040
rect 65962 513984 66030 514040
rect 66086 513984 66154 514040
rect 66210 513984 66278 514040
rect 66334 513984 66402 514040
rect 66458 513984 597980 514040
rect -1916 513978 597980 513984
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513916 597980 513922
rect -1916 513860 60202 513916
rect 60258 513860 60326 513916
rect 60382 513860 60450 513916
rect 60506 513860 60574 513916
rect 60630 513860 60698 513916
rect 60754 513860 60822 513916
rect 60878 513860 60946 513916
rect 61002 513860 61070 513916
rect 61126 513860 61194 513916
rect 61250 513860 61318 513916
rect 61374 513860 61442 513916
rect 61498 513860 61566 513916
rect 61622 513860 61690 513916
rect 61746 513860 61814 513916
rect 61870 513860 61938 513916
rect 61994 513860 62062 513916
rect 62118 513860 62186 513916
rect 62242 513860 62310 513916
rect 62366 513860 62434 513916
rect 62490 513860 62558 513916
rect 62614 513860 62682 513916
rect 62738 513860 62806 513916
rect 62862 513860 62930 513916
rect 62986 513860 63054 513916
rect 63110 513860 63178 513916
rect 63234 513860 63302 513916
rect 63358 513860 63426 513916
rect 63482 513860 63550 513916
rect 63606 513860 63674 513916
rect 63730 513860 63798 513916
rect 63854 513860 63922 513916
rect 63978 513860 64046 513916
rect 64102 513860 64170 513916
rect 64226 513860 64294 513916
rect 64350 513860 64418 513916
rect 64474 513860 64542 513916
rect 64598 513860 64666 513916
rect 64722 513860 64790 513916
rect 64846 513860 64914 513916
rect 64970 513860 65038 513916
rect 65094 513860 65162 513916
rect 65218 513860 65286 513916
rect 65342 513860 65410 513916
rect 65466 513860 65534 513916
rect 65590 513860 65658 513916
rect 65714 513860 65782 513916
rect 65838 513860 65906 513916
rect 65962 513860 66030 513916
rect 66086 513860 66154 513916
rect 66210 513860 66278 513916
rect 66334 513860 66402 513916
rect 66458 513860 597980 513916
rect -1916 513826 597980 513860
rect -1916 508435 597980 508446
rect -1916 508379 90112 508435
rect 90168 508379 90236 508435
rect 90292 508379 90360 508435
rect 90416 508379 90484 508435
rect 90540 508379 90608 508435
rect 90664 508379 90732 508435
rect 90788 508379 90856 508435
rect 90912 508379 90980 508435
rect 91036 508379 91104 508435
rect 91160 508379 91228 508435
rect 91284 508379 91352 508435
rect 91408 508379 91476 508435
rect 91532 508379 91600 508435
rect 91656 508379 91724 508435
rect 91780 508379 91848 508435
rect 91904 508379 91972 508435
rect 92028 508379 92096 508435
rect 92152 508379 92220 508435
rect 92276 508379 92344 508435
rect 92400 508379 92468 508435
rect 92524 508379 92592 508435
rect 92648 508379 92716 508435
rect 92772 508379 92840 508435
rect 92896 508379 92964 508435
rect 93020 508379 93088 508435
rect 93144 508379 93212 508435
rect 93268 508379 93336 508435
rect 93392 508379 93460 508435
rect 93516 508379 93584 508435
rect 93640 508379 93708 508435
rect 93764 508379 93832 508435
rect 93888 508379 93956 508435
rect 94012 508379 94080 508435
rect 94136 508379 94204 508435
rect 94260 508379 94328 508435
rect 94384 508379 94452 508435
rect 94508 508379 94576 508435
rect 94632 508379 94700 508435
rect 94756 508379 94824 508435
rect 94880 508379 94948 508435
rect 95004 508379 95072 508435
rect 95128 508379 95196 508435
rect 95252 508379 95320 508435
rect 95376 508379 95444 508435
rect 95500 508379 95568 508435
rect 95624 508379 95692 508435
rect 95748 508379 95816 508435
rect 95872 508379 95940 508435
rect 95996 508379 96064 508435
rect 96120 508379 96188 508435
rect 96244 508379 96312 508435
rect 96368 508379 96436 508435
rect 96492 508379 96560 508435
rect 96616 508379 96684 508435
rect 96740 508379 96808 508435
rect 96864 508379 96932 508435
rect 96988 508379 97056 508435
rect 97112 508379 97180 508435
rect 97236 508379 97304 508435
rect 97360 508379 97428 508435
rect 97484 508379 97552 508435
rect 97608 508379 97676 508435
rect 97732 508379 97800 508435
rect 97856 508379 97924 508435
rect 97980 508379 98048 508435
rect 98104 508379 98172 508435
rect 98228 508379 98296 508435
rect 98352 508379 98420 508435
rect 98476 508379 98544 508435
rect 98600 508379 98668 508435
rect 98724 508379 98792 508435
rect 98848 508379 98916 508435
rect 98972 508379 99040 508435
rect 99096 508379 99164 508435
rect 99220 508379 99288 508435
rect 99344 508379 99412 508435
rect 99468 508379 99536 508435
rect 99592 508379 99660 508435
rect 99716 508379 99784 508435
rect 99840 508379 99908 508435
rect 99964 508379 100032 508435
rect 100088 508379 597980 508435
rect -1916 508350 597980 508379
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508311 159114 508350
rect 36662 508294 90112 508311
rect -1916 508255 90112 508294
rect 90168 508255 90236 508311
rect 90292 508255 90360 508311
rect 90416 508255 90484 508311
rect 90540 508255 90608 508311
rect 90664 508255 90732 508311
rect 90788 508255 90856 508311
rect 90912 508255 90980 508311
rect 91036 508255 91104 508311
rect 91160 508255 91228 508311
rect 91284 508255 91352 508311
rect 91408 508255 91476 508311
rect 91532 508255 91600 508311
rect 91656 508255 91724 508311
rect 91780 508255 91848 508311
rect 91904 508255 91972 508311
rect 92028 508255 92096 508311
rect 92152 508255 92220 508311
rect 92276 508255 92344 508311
rect 92400 508255 92468 508311
rect 92524 508255 92592 508311
rect 92648 508255 92716 508311
rect 92772 508255 92840 508311
rect 92896 508255 92964 508311
rect 93020 508255 93088 508311
rect 93144 508255 93212 508311
rect 93268 508255 93336 508311
rect 93392 508255 93460 508311
rect 93516 508255 93584 508311
rect 93640 508255 93708 508311
rect 93764 508255 93832 508311
rect 93888 508255 93956 508311
rect 94012 508255 94080 508311
rect 94136 508255 94204 508311
rect 94260 508255 94328 508311
rect 94384 508255 94452 508311
rect 94508 508255 94576 508311
rect 94632 508255 94700 508311
rect 94756 508255 94824 508311
rect 94880 508255 94948 508311
rect 95004 508255 95072 508311
rect 95128 508255 95196 508311
rect 95252 508255 95320 508311
rect 95376 508255 95444 508311
rect 95500 508255 95568 508311
rect 95624 508255 95692 508311
rect 95748 508255 95816 508311
rect 95872 508255 95940 508311
rect 95996 508255 96064 508311
rect 96120 508255 96188 508311
rect 96244 508255 96312 508311
rect 96368 508255 96436 508311
rect 96492 508255 96560 508311
rect 96616 508255 96684 508311
rect 96740 508255 96808 508311
rect 96864 508255 96932 508311
rect 96988 508255 97056 508311
rect 97112 508255 97180 508311
rect 97236 508255 97304 508311
rect 97360 508255 97428 508311
rect 97484 508255 97552 508311
rect 97608 508255 97676 508311
rect 97732 508255 97800 508311
rect 97856 508255 97924 508311
rect 97980 508255 98048 508311
rect 98104 508255 98172 508311
rect 98228 508255 98296 508311
rect 98352 508255 98420 508311
rect 98476 508255 98544 508311
rect 98600 508255 98668 508311
rect 98724 508255 98792 508311
rect 98848 508255 98916 508311
rect 98972 508255 99040 508311
rect 99096 508255 99164 508311
rect 99220 508255 99288 508311
rect 99344 508255 99412 508311
rect 99468 508255 99536 508311
rect 99592 508255 99660 508311
rect 99716 508255 99784 508311
rect 99840 508255 99908 508311
rect 99964 508255 100032 508311
rect 100088 508294 159114 508311
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect 100088 508255 597980 508294
rect -1916 508226 597980 508255
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508187 159114 508226
rect 36662 508170 90112 508187
rect -1916 508131 90112 508170
rect 90168 508131 90236 508187
rect 90292 508131 90360 508187
rect 90416 508131 90484 508187
rect 90540 508131 90608 508187
rect 90664 508131 90732 508187
rect 90788 508131 90856 508187
rect 90912 508131 90980 508187
rect 91036 508131 91104 508187
rect 91160 508131 91228 508187
rect 91284 508131 91352 508187
rect 91408 508131 91476 508187
rect 91532 508131 91600 508187
rect 91656 508131 91724 508187
rect 91780 508131 91848 508187
rect 91904 508131 91972 508187
rect 92028 508131 92096 508187
rect 92152 508131 92220 508187
rect 92276 508131 92344 508187
rect 92400 508131 92468 508187
rect 92524 508131 92592 508187
rect 92648 508131 92716 508187
rect 92772 508131 92840 508187
rect 92896 508131 92964 508187
rect 93020 508131 93088 508187
rect 93144 508131 93212 508187
rect 93268 508131 93336 508187
rect 93392 508131 93460 508187
rect 93516 508131 93584 508187
rect 93640 508131 93708 508187
rect 93764 508131 93832 508187
rect 93888 508131 93956 508187
rect 94012 508131 94080 508187
rect 94136 508131 94204 508187
rect 94260 508131 94328 508187
rect 94384 508131 94452 508187
rect 94508 508131 94576 508187
rect 94632 508131 94700 508187
rect 94756 508131 94824 508187
rect 94880 508131 94948 508187
rect 95004 508131 95072 508187
rect 95128 508131 95196 508187
rect 95252 508131 95320 508187
rect 95376 508131 95444 508187
rect 95500 508131 95568 508187
rect 95624 508131 95692 508187
rect 95748 508131 95816 508187
rect 95872 508131 95940 508187
rect 95996 508131 96064 508187
rect 96120 508131 96188 508187
rect 96244 508131 96312 508187
rect 96368 508131 96436 508187
rect 96492 508131 96560 508187
rect 96616 508131 96684 508187
rect 96740 508131 96808 508187
rect 96864 508131 96932 508187
rect 96988 508131 97056 508187
rect 97112 508131 97180 508187
rect 97236 508131 97304 508187
rect 97360 508131 97428 508187
rect 97484 508131 97552 508187
rect 97608 508131 97676 508187
rect 97732 508131 97800 508187
rect 97856 508131 97924 508187
rect 97980 508131 98048 508187
rect 98104 508131 98172 508187
rect 98228 508131 98296 508187
rect 98352 508131 98420 508187
rect 98476 508131 98544 508187
rect 98600 508131 98668 508187
rect 98724 508131 98792 508187
rect 98848 508131 98916 508187
rect 98972 508131 99040 508187
rect 99096 508131 99164 508187
rect 99220 508131 99288 508187
rect 99344 508131 99412 508187
rect 99468 508131 99536 508187
rect 99592 508131 99660 508187
rect 99716 508131 99784 508187
rect 99840 508131 99908 508187
rect 99964 508131 100032 508187
rect 100088 508170 159114 508187
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect 100088 508131 597980 508170
rect -1916 508102 597980 508131
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507911 597980 507922
rect -1916 507855 89904 507911
rect 89960 507855 90028 507911
rect 90084 507855 90152 507911
rect 90208 507855 90276 507911
rect 90332 507855 90400 507911
rect 90456 507855 90524 507911
rect 90580 507855 90648 507911
rect 90704 507855 90772 507911
rect 90828 507855 90896 507911
rect 90952 507855 91020 507911
rect 91076 507855 91144 507911
rect 91200 507855 91268 507911
rect 91324 507855 91392 507911
rect 91448 507855 91516 507911
rect 91572 507855 91640 507911
rect 91696 507855 91764 507911
rect 91820 507855 91888 507911
rect 91944 507855 92012 507911
rect 92068 507855 92136 507911
rect 92192 507855 92260 507911
rect 92316 507855 92384 507911
rect 92440 507855 92508 507911
rect 92564 507855 92632 507911
rect 92688 507855 92756 507911
rect 92812 507855 92880 507911
rect 92936 507855 93004 507911
rect 93060 507855 93128 507911
rect 93184 507855 93252 507911
rect 93308 507855 93376 507911
rect 93432 507855 93500 507911
rect 93556 507855 93624 507911
rect 93680 507855 93748 507911
rect 93804 507855 93872 507911
rect 93928 507855 93996 507911
rect 94052 507855 94120 507911
rect 94176 507855 94244 507911
rect 94300 507855 94368 507911
rect 94424 507855 94492 507911
rect 94548 507855 94616 507911
rect 94672 507855 94740 507911
rect 94796 507855 94864 507911
rect 94920 507855 94988 507911
rect 95044 507855 95112 507911
rect 95168 507855 95236 507911
rect 95292 507855 95360 507911
rect 95416 507855 95484 507911
rect 95540 507855 95608 507911
rect 95664 507855 95732 507911
rect 95788 507855 95856 507911
rect 95912 507855 95980 507911
rect 96036 507855 96104 507911
rect 96160 507855 96228 507911
rect 96284 507855 96352 507911
rect 96408 507855 96476 507911
rect 96532 507855 96600 507911
rect 96656 507855 96724 507911
rect 96780 507855 96848 507911
rect 96904 507855 96972 507911
rect 97028 507855 97096 507911
rect 97152 507855 97220 507911
rect 97276 507855 97344 507911
rect 97400 507855 97468 507911
rect 97524 507855 97592 507911
rect 97648 507855 97716 507911
rect 97772 507855 97840 507911
rect 97896 507855 97964 507911
rect 98020 507855 98088 507911
rect 98144 507855 98212 507911
rect 98268 507855 98336 507911
rect 98392 507855 98460 507911
rect 98516 507855 98584 507911
rect 98640 507855 98708 507911
rect 98764 507855 98832 507911
rect 98888 507855 98956 507911
rect 99012 507855 99080 507911
rect 99136 507855 99204 507911
rect 99260 507855 99328 507911
rect 99384 507855 99452 507911
rect 99508 507855 99576 507911
rect 99632 507855 99700 507911
rect 99756 507855 597980 507911
rect -1916 507826 597980 507855
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496212 162834 496226
rect 40382 496170 63430 496212
rect -1916 496156 63430 496170
rect 63486 496156 63554 496212
rect 63610 496156 63678 496212
rect 63734 496156 63802 496212
rect 63858 496156 63926 496212
rect 63982 496156 64050 496212
rect 64106 496156 64174 496212
rect 64230 496156 64298 496212
rect 64354 496156 64422 496212
rect 64478 496156 64546 496212
rect 64602 496156 64670 496212
rect 64726 496156 64794 496212
rect 64850 496156 64918 496212
rect 64974 496156 65042 496212
rect 65098 496156 65166 496212
rect 65222 496156 65290 496212
rect 65346 496156 65414 496212
rect 65470 496156 65538 496212
rect 65594 496156 65662 496212
rect 65718 496156 65786 496212
rect 65842 496156 65910 496212
rect 65966 496156 66034 496212
rect 66090 496156 66158 496212
rect 66214 496156 66282 496212
rect 66338 496156 66406 496212
rect 66462 496156 66530 496212
rect 66586 496156 66654 496212
rect 66710 496156 66778 496212
rect 66834 496156 66902 496212
rect 66958 496156 67026 496212
rect 67082 496156 67150 496212
rect 67206 496156 67274 496212
rect 67330 496156 67398 496212
rect 67454 496156 67522 496212
rect 67578 496156 67646 496212
rect 67702 496156 67770 496212
rect 67826 496156 67894 496212
rect 67950 496156 68018 496212
rect 68074 496156 68142 496212
rect 68198 496156 68266 496212
rect 68322 496156 68390 496212
rect 68446 496156 68514 496212
rect 68570 496156 68638 496212
rect 68694 496156 68762 496212
rect 68818 496156 68886 496212
rect 68942 496156 69010 496212
rect 69066 496156 69134 496212
rect 69190 496156 69258 496212
rect 69314 496156 69382 496212
rect 69438 496156 69506 496212
rect 69562 496156 69630 496212
rect 69686 496156 69754 496212
rect 69810 496156 69878 496212
rect 69934 496156 70002 496212
rect 70058 496156 70126 496212
rect 70182 496156 70250 496212
rect 70306 496156 70374 496212
rect 70430 496170 162834 496212
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 70430 496156 597980 496170
rect -1916 496102 597980 496156
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496088 162834 496102
rect 40382 496046 63430 496088
rect -1916 496032 63430 496046
rect 63486 496032 63554 496088
rect 63610 496032 63678 496088
rect 63734 496032 63802 496088
rect 63858 496032 63926 496088
rect 63982 496032 64050 496088
rect 64106 496032 64174 496088
rect 64230 496032 64298 496088
rect 64354 496032 64422 496088
rect 64478 496032 64546 496088
rect 64602 496032 64670 496088
rect 64726 496032 64794 496088
rect 64850 496032 64918 496088
rect 64974 496032 65042 496088
rect 65098 496032 65166 496088
rect 65222 496032 65290 496088
rect 65346 496032 65414 496088
rect 65470 496032 65538 496088
rect 65594 496032 65662 496088
rect 65718 496032 65786 496088
rect 65842 496032 65910 496088
rect 65966 496032 66034 496088
rect 66090 496032 66158 496088
rect 66214 496032 66282 496088
rect 66338 496032 66406 496088
rect 66462 496032 66530 496088
rect 66586 496032 66654 496088
rect 66710 496032 66778 496088
rect 66834 496032 66902 496088
rect 66958 496032 67026 496088
rect 67082 496032 67150 496088
rect 67206 496032 67274 496088
rect 67330 496032 67398 496088
rect 67454 496032 67522 496088
rect 67578 496032 67646 496088
rect 67702 496032 67770 496088
rect 67826 496032 67894 496088
rect 67950 496032 68018 496088
rect 68074 496032 68142 496088
rect 68198 496032 68266 496088
rect 68322 496032 68390 496088
rect 68446 496032 68514 496088
rect 68570 496032 68638 496088
rect 68694 496032 68762 496088
rect 68818 496032 68886 496088
rect 68942 496032 69010 496088
rect 69066 496032 69134 496088
rect 69190 496032 69258 496088
rect 69314 496032 69382 496088
rect 69438 496032 69506 496088
rect 69562 496032 69630 496088
rect 69686 496032 69754 496088
rect 69810 496032 69878 496088
rect 69934 496032 70002 496088
rect 70058 496032 70126 496088
rect 70182 496032 70250 496088
rect 70306 496032 70374 496088
rect 70430 496046 162834 496088
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 70430 496032 597980 496046
rect -1916 495978 597980 496032
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495964 162834 495978
rect 40382 495922 63430 495964
rect -1916 495908 63430 495922
rect 63486 495908 63554 495964
rect 63610 495908 63678 495964
rect 63734 495908 63802 495964
rect 63858 495908 63926 495964
rect 63982 495908 64050 495964
rect 64106 495908 64174 495964
rect 64230 495908 64298 495964
rect 64354 495908 64422 495964
rect 64478 495908 64546 495964
rect 64602 495908 64670 495964
rect 64726 495908 64794 495964
rect 64850 495908 64918 495964
rect 64974 495908 65042 495964
rect 65098 495908 65166 495964
rect 65222 495908 65290 495964
rect 65346 495908 65414 495964
rect 65470 495908 65538 495964
rect 65594 495908 65662 495964
rect 65718 495908 65786 495964
rect 65842 495908 65910 495964
rect 65966 495908 66034 495964
rect 66090 495908 66158 495964
rect 66214 495908 66282 495964
rect 66338 495908 66406 495964
rect 66462 495908 66530 495964
rect 66586 495908 66654 495964
rect 66710 495908 66778 495964
rect 66834 495908 66902 495964
rect 66958 495908 67026 495964
rect 67082 495908 67150 495964
rect 67206 495908 67274 495964
rect 67330 495908 67398 495964
rect 67454 495908 67522 495964
rect 67578 495908 67646 495964
rect 67702 495908 67770 495964
rect 67826 495908 67894 495964
rect 67950 495908 68018 495964
rect 68074 495908 68142 495964
rect 68198 495908 68266 495964
rect 68322 495908 68390 495964
rect 68446 495908 68514 495964
rect 68570 495908 68638 495964
rect 68694 495908 68762 495964
rect 68818 495908 68886 495964
rect 68942 495908 69010 495964
rect 69066 495908 69134 495964
rect 69190 495908 69258 495964
rect 69314 495908 69382 495964
rect 69438 495908 69506 495964
rect 69562 495908 69630 495964
rect 69686 495908 69754 495964
rect 69810 495908 69878 495964
rect 69934 495908 70002 495964
rect 70058 495908 70126 495964
rect 70182 495908 70250 495964
rect 70306 495908 70374 495964
rect 70430 495922 162834 495964
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 70430 495908 597980 495922
rect -1916 495826 597980 495908
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490272 597980 490294
rect -1916 490226 85236 490272
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490216 85236 490226
rect 85292 490216 85360 490272
rect 85416 490216 85484 490272
rect 85540 490216 85608 490272
rect 85664 490216 85732 490272
rect 85788 490216 85856 490272
rect 85912 490216 85980 490272
rect 86036 490216 86104 490272
rect 86160 490216 86228 490272
rect 86284 490216 86352 490272
rect 86408 490216 86476 490272
rect 86532 490216 86600 490272
rect 86656 490216 86724 490272
rect 86780 490216 86848 490272
rect 86904 490216 86972 490272
rect 87028 490216 87096 490272
rect 87152 490216 87220 490272
rect 87276 490216 87344 490272
rect 87400 490216 87468 490272
rect 87524 490216 87592 490272
rect 87648 490216 87716 490272
rect 87772 490216 87840 490272
rect 87896 490216 87964 490272
rect 88020 490216 88088 490272
rect 88144 490216 88212 490272
rect 88268 490216 88336 490272
rect 88392 490216 88460 490272
rect 88516 490216 88584 490272
rect 88640 490216 88708 490272
rect 88764 490226 597980 490272
rect 88764 490216 159114 490226
rect 36662 490170 159114 490216
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490148 597980 490170
rect -1916 490102 85236 490148
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490092 85236 490102
rect 85292 490092 85360 490148
rect 85416 490092 85484 490148
rect 85540 490092 85608 490148
rect 85664 490092 85732 490148
rect 85788 490092 85856 490148
rect 85912 490092 85980 490148
rect 86036 490092 86104 490148
rect 86160 490092 86228 490148
rect 86284 490092 86352 490148
rect 86408 490092 86476 490148
rect 86532 490092 86600 490148
rect 86656 490092 86724 490148
rect 86780 490092 86848 490148
rect 86904 490092 86972 490148
rect 87028 490092 87096 490148
rect 87152 490092 87220 490148
rect 87276 490092 87344 490148
rect 87400 490092 87468 490148
rect 87524 490092 87592 490148
rect 87648 490092 87716 490148
rect 87772 490092 87840 490148
rect 87896 490092 87964 490148
rect 88020 490092 88088 490148
rect 88144 490092 88212 490148
rect 88268 490092 88336 490148
rect 88392 490092 88460 490148
rect 88516 490092 88584 490148
rect 88640 490092 88708 490148
rect 88764 490102 597980 490148
rect 88764 490092 159114 490102
rect 36662 490046 159114 490092
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 490024 597980 490046
rect -1916 489978 85236 490024
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489968 85236 489978
rect 85292 489968 85360 490024
rect 85416 489968 85484 490024
rect 85540 489968 85608 490024
rect 85664 489968 85732 490024
rect 85788 489968 85856 490024
rect 85912 489968 85980 490024
rect 86036 489968 86104 490024
rect 86160 489968 86228 490024
rect 86284 489968 86352 490024
rect 86408 489968 86476 490024
rect 86532 489968 86600 490024
rect 86656 489968 86724 490024
rect 86780 489968 86848 490024
rect 86904 489968 86972 490024
rect 87028 489968 87096 490024
rect 87152 489968 87220 490024
rect 87276 489968 87344 490024
rect 87400 489968 87468 490024
rect 87524 489968 87592 490024
rect 87648 489968 87716 490024
rect 87772 489968 87840 490024
rect 87896 489968 87964 490024
rect 88020 489968 88088 490024
rect 88144 489968 88212 490024
rect 88268 489968 88336 490024
rect 88392 489968 88460 490024
rect 88516 489968 88584 490024
rect 88640 489968 88708 490024
rect 88764 489978 597980 490024
rect 88764 489968 159114 489978
rect 36662 489922 159114 489968
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478358 597980 478446
rect -1916 478350 80936 478358
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478302 80936 478350
rect 80992 478302 81060 478358
rect 81116 478302 81184 478358
rect 81240 478302 81308 478358
rect 81364 478350 597980 478358
rect 81364 478302 132114 478350
rect 71102 478294 132114 478302
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect 4156 416818 83988 416834
rect 4156 416762 4172 416818
rect 4228 416762 83916 416818
rect 83972 416762 83988 416818
rect 4156 416746 83988 416762
rect 4268 410698 202372 410714
rect 4268 410642 4284 410698
rect 4340 410642 202300 410698
rect 202356 410642 202372 410698
rect 4268 410626 202372 410642
rect 336908 410518 354692 410534
rect 336908 410462 336924 410518
rect 336980 410462 354620 410518
rect 354676 410462 354692 410518
rect 336908 410446 354692 410462
rect 359980 410518 366004 410534
rect 359980 410462 359996 410518
rect 360052 410462 365932 410518
rect 365988 410462 366004 410518
rect 359980 410446 366004 410462
rect 297260 410338 499396 410354
rect 297260 410282 297276 410338
rect 297332 410282 499324 410338
rect 499380 410282 499396 410338
rect 297260 410266 499396 410282
rect 352812 410158 359844 410174
rect 352812 410102 352828 410158
rect 352884 410102 359772 410158
rect 359828 410102 359844 410158
rect 352812 410086 359844 410102
rect 366252 410158 371380 410174
rect 366252 410102 366268 410158
rect 366324 410102 371308 410158
rect 371364 410102 371380 410158
rect 366252 410086 371380 410102
rect 386188 410158 404980 410174
rect 386188 410102 386204 410158
rect 386260 410102 404908 410158
rect 404964 410102 404980 410158
rect 386188 410086 404980 410102
rect 354716 409978 359732 409994
rect 354716 409922 354732 409978
rect 354788 409922 359660 409978
rect 359716 409922 359732 409978
rect 354716 409906 359732 409922
rect 369612 409978 386164 409994
rect 369612 409922 369628 409978
rect 369684 409922 386092 409978
rect 386148 409922 386164 409978
rect 369612 409906 386164 409922
rect 261980 409618 359620 409634
rect 261980 409562 261996 409618
rect 262052 409562 359548 409618
rect 359604 409562 359620 409618
rect 261980 409546 359620 409562
rect 4380 409438 278980 409454
rect 4380 409382 4396 409438
rect 4452 409382 278908 409438
rect 278964 409382 278980 409438
rect 4380 409366 278980 409382
rect 4492 409258 288164 409274
rect 4492 409202 4508 409258
rect 4564 409202 288092 409258
rect 288148 409202 288164 409258
rect 4492 409186 288164 409202
rect 243500 409078 532660 409094
rect 243500 409022 243516 409078
rect 243572 409022 532588 409078
rect 532644 409022 532660 409078
rect 243500 409006 532660 409022
rect 340828 408898 356260 408914
rect 340828 408842 340844 408898
rect 340900 408842 356188 408898
rect 356244 408842 356260 408898
rect 340828 408826 356260 408842
rect 295580 408718 366228 408734
rect 295580 408662 295596 408718
rect 295652 408662 366156 408718
rect 366212 408662 366228 408718
rect 295580 408646 366228 408662
rect 356620 408538 496484 408554
rect 356620 408482 356636 408538
rect 356692 408482 496412 408538
rect 496468 408482 496484 408538
rect 356620 408466 496484 408482
rect 298940 408358 514180 408374
rect 298940 408302 298956 408358
rect 299012 408302 514108 408358
rect 514164 408302 514180 408358
rect 298940 408286 514180 408302
rect 354492 408178 558308 408194
rect 354492 408122 354508 408178
rect 354564 408122 558236 408178
rect 558292 408122 558308 408178
rect 354492 408106 558308 408122
rect 305660 407638 580708 407654
rect 305660 407582 305676 407638
rect 305732 407582 580636 407638
rect 580692 407582 580708 407638
rect 305660 407566 580708 407582
rect 240252 407458 335204 407474
rect 240252 407402 240268 407458
rect 240324 407402 335132 407458
rect 335188 407402 335204 407458
rect 240252 407386 335204 407402
rect 246860 407278 336100 407294
rect 246860 407222 246876 407278
rect 246932 407222 336028 407278
rect 336084 407222 336100 407278
rect 246860 407206 336100 407222
rect 339596 407278 528964 407294
rect 339596 407222 339612 407278
rect 339668 407222 528892 407278
rect 528948 407222 528964 407278
rect 339596 407206 528964 407222
rect 302300 407098 543748 407114
rect 302300 407042 302316 407098
rect 302372 407042 543676 407098
rect 543732 407042 543748 407098
rect 302300 407026 543748 407042
rect 302188 406918 551140 406934
rect 302188 406862 302204 406918
rect 302260 406862 551068 406918
rect 551124 406862 551140 406918
rect 302188 406846 551140 406862
rect 203292 406738 232388 406754
rect 203292 406682 203308 406738
rect 203364 406682 232316 406738
rect 232372 406682 232388 406738
rect 203292 406666 232388 406682
rect 337468 406738 352228 406754
rect 337468 406682 337484 406738
rect 337540 406682 352156 406738
rect 352212 406682 352228 406738
rect 337468 406666 352228 406682
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 66574 406350
rect 66630 406294 66698 406350
rect 66754 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71894 406350
rect 71950 406294 72018 406350
rect 72074 406294 77214 406350
rect 77270 406294 77338 406350
rect 77394 406294 82534 406350
rect 82590 406294 82658 406350
rect 82714 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 66574 406226
rect 66630 406170 66698 406226
rect 66754 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71894 406226
rect 71950 406170 72018 406226
rect 72074 406170 77214 406226
rect 77270 406170 77338 406226
rect 77394 406170 82534 406226
rect 82590 406170 82658 406226
rect 82714 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 66574 406102
rect 66630 406046 66698 406102
rect 66754 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71894 406102
rect 71950 406046 72018 406102
rect 72074 406046 77214 406102
rect 77270 406046 77338 406102
rect 77394 406046 82534 406102
rect 82590 406046 82658 406102
rect 82714 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 66574 405978
rect 66630 405922 66698 405978
rect 66754 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71894 405978
rect 71950 405922 72018 405978
rect 72074 405922 77214 405978
rect 77270 405922 77338 405978
rect 77394 405922 82534 405978
rect 82590 405922 82658 405978
rect 82714 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect 303980 405658 383140 405674
rect 303980 405602 303996 405658
rect 304052 405602 383068 405658
rect 383124 405602 383140 405658
rect 303980 405586 383140 405602
rect 340156 404938 357380 404954
rect 340156 404882 340172 404938
rect 340228 404882 357308 404938
rect 357364 404882 357380 404938
rect 340156 404866 357380 404882
rect 338476 404758 366116 404774
rect 338476 404702 338492 404758
rect 338548 404702 366044 404758
rect 366100 404702 366116 404758
rect 338476 404686 366116 404702
rect 346092 404398 354580 404414
rect 346092 404342 346108 404398
rect 346164 404342 354508 404398
rect 354564 404342 354580 404398
rect 346092 404326 354580 404342
rect 189180 404218 200020 404234
rect 189180 404162 189196 404218
rect 189252 404162 199948 404218
rect 200004 404162 200020 404218
rect 189180 404146 200020 404162
rect 339484 404218 522244 404234
rect 339484 404162 339500 404218
rect 339556 404162 522172 404218
rect 522228 404162 522244 404218
rect 339484 404146 522244 404162
rect 57916 404038 206740 404054
rect 57916 403982 57932 404038
rect 57988 403982 206668 404038
rect 206724 403982 206740 404038
rect 57916 403966 206740 403982
rect 300620 404038 366228 404054
rect 300620 403982 300636 404038
rect 300692 403982 366156 404038
rect 366212 403982 366228 404038
rect 300620 403966 366228 403982
rect 372916 404038 582164 404054
rect 372916 403982 582092 404038
rect 582148 403982 582164 404038
rect 372916 403966 582164 403982
rect 372916 403874 373004 403966
rect 365916 403858 373004 403874
rect 365916 403802 365932 403858
rect 365988 403802 373004 403858
rect 365916 403786 373004 403802
rect 341500 403498 347972 403514
rect 341500 403442 341516 403498
rect 341572 403442 347900 403498
rect 347956 403442 347972 403498
rect 341500 403426 347972 403442
rect 340940 403318 342932 403334
rect 340940 403262 340956 403318
rect 341012 403262 342932 403318
rect 340940 403246 342932 403262
rect 342844 403154 342932 403246
rect 376220 403318 383140 403334
rect 376220 403262 383068 403318
rect 383124 403262 383140 403318
rect 376220 403246 383140 403262
rect 342844 403138 350996 403154
rect 342844 403082 350924 403138
rect 350980 403082 350996 403138
rect 342844 403066 350996 403082
rect 364796 403138 373004 403154
rect 364796 403082 364812 403138
rect 364868 403082 373004 403138
rect 364796 403066 373004 403082
rect 372916 402974 373004 403066
rect 376220 402974 376308 403246
rect 338700 402958 350548 402974
rect 338700 402902 338716 402958
rect 338772 402902 350476 402958
rect 350532 402902 350548 402958
rect 338700 402886 350548 402902
rect 350684 402958 366228 402974
rect 350684 402902 350700 402958
rect 350756 402902 366156 402958
rect 366212 402902 366228 402958
rect 350684 402886 366228 402902
rect 372916 402886 376308 402974
rect 384676 403138 565924 403154
rect 384676 403082 565852 403138
rect 565908 403082 565924 403138
rect 384676 403066 565924 403082
rect 384676 402794 384764 403066
rect 293900 402778 350884 402794
rect 293900 402722 293916 402778
rect 293972 402722 350812 402778
rect 350868 402722 350884 402778
rect 293900 402706 350884 402722
rect 367932 402778 384764 402794
rect 367932 402722 367948 402778
rect 368004 402722 384764 402778
rect 367932 402706 384764 402722
rect 339036 402598 511940 402614
rect 339036 402542 339052 402598
rect 339108 402542 511868 402598
rect 511924 402542 511940 402598
rect 339036 402526 511940 402542
rect 12556 402418 208420 402434
rect 12556 402362 12572 402418
rect 12628 402362 208348 402418
rect 208404 402362 208420 402418
rect 12556 402346 208420 402362
rect 278780 402418 517092 402434
rect 278780 402362 278796 402418
rect 278852 402362 517020 402418
rect 517076 402362 517092 402418
rect 278780 402346 517092 402362
rect 352700 401518 358612 401534
rect 352700 401462 352716 401518
rect 352772 401462 358540 401518
rect 358596 401462 358612 401518
rect 352700 401446 358612 401462
rect 361212 401518 367908 401534
rect 361212 401462 361228 401518
rect 361284 401462 367836 401518
rect 367892 401462 367908 401518
rect 361212 401446 367908 401462
rect 337636 401158 346180 401174
rect 337636 401102 346108 401158
rect 346164 401102 346180 401158
rect 337636 401086 346180 401102
rect 337636 400814 337724 401086
rect 303868 400798 337724 400814
rect 303868 400742 303884 400798
rect 303940 400742 337724 400798
rect 303868 400726 337724 400742
rect 263660 400618 341588 400634
rect 263660 400562 263676 400618
rect 263732 400562 341516 400618
rect 341572 400562 341588 400618
rect 263660 400546 341588 400562
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 63914 400350
rect 63970 400294 64038 400350
rect 64094 400294 69234 400350
rect 69290 400294 69358 400350
rect 69414 400294 74554 400350
rect 74610 400294 74678 400350
rect 74734 400294 79874 400350
rect 79930 400294 79998 400350
rect 80054 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 344518 400350
rect 344574 400294 344642 400350
rect 344698 400294 375238 400350
rect 375294 400294 375362 400350
rect 375418 400294 405958 400350
rect 406014 400294 406082 400350
rect 406138 400294 436678 400350
rect 436734 400294 436802 400350
rect 436858 400294 467398 400350
rect 467454 400294 467522 400350
rect 467578 400294 498118 400350
rect 498174 400294 498242 400350
rect 498298 400294 528838 400350
rect 528894 400294 528962 400350
rect 529018 400294 559558 400350
rect 559614 400294 559682 400350
rect 559738 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 63914 400226
rect 63970 400170 64038 400226
rect 64094 400170 69234 400226
rect 69290 400170 69358 400226
rect 69414 400170 74554 400226
rect 74610 400170 74678 400226
rect 74734 400170 79874 400226
rect 79930 400170 79998 400226
rect 80054 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 344518 400226
rect 344574 400170 344642 400226
rect 344698 400170 375238 400226
rect 375294 400170 375362 400226
rect 375418 400170 405958 400226
rect 406014 400170 406082 400226
rect 406138 400170 436678 400226
rect 436734 400170 436802 400226
rect 436858 400170 467398 400226
rect 467454 400170 467522 400226
rect 467578 400170 498118 400226
rect 498174 400170 498242 400226
rect 498298 400170 528838 400226
rect 528894 400170 528962 400226
rect 529018 400170 559558 400226
rect 559614 400170 559682 400226
rect 559738 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 63914 400102
rect 63970 400046 64038 400102
rect 64094 400046 69234 400102
rect 69290 400046 69358 400102
rect 69414 400046 74554 400102
rect 74610 400046 74678 400102
rect 74734 400046 79874 400102
rect 79930 400046 79998 400102
rect 80054 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 344518 400102
rect 344574 400046 344642 400102
rect 344698 400046 375238 400102
rect 375294 400046 375362 400102
rect 375418 400046 405958 400102
rect 406014 400046 406082 400102
rect 406138 400046 436678 400102
rect 436734 400046 436802 400102
rect 436858 400046 467398 400102
rect 467454 400046 467522 400102
rect 467578 400046 498118 400102
rect 498174 400046 498242 400102
rect 498298 400046 528838 400102
rect 528894 400046 528962 400102
rect 529018 400046 559558 400102
rect 559614 400046 559682 400102
rect 559738 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 63914 399978
rect 63970 399922 64038 399978
rect 64094 399922 69234 399978
rect 69290 399922 69358 399978
rect 69414 399922 74554 399978
rect 74610 399922 74678 399978
rect 74734 399922 79874 399978
rect 79930 399922 79998 399978
rect 80054 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 344518 399978
rect 344574 399922 344642 399978
rect 344698 399922 375238 399978
rect 375294 399922 375362 399978
rect 375418 399922 405958 399978
rect 406014 399922 406082 399978
rect 406138 399922 436678 399978
rect 436734 399922 436802 399978
rect 436858 399922 467398 399978
rect 467454 399922 467522 399978
rect 467578 399922 498118 399978
rect 498174 399922 498242 399978
rect 498298 399922 528838 399978
rect 528894 399922 528962 399978
rect 529018 399922 559558 399978
rect 559614 399922 559682 399978
rect 559738 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 337692 399718 341252 399734
rect 337692 399662 337708 399718
rect 337764 399662 341180 399718
rect 341236 399662 341252 399718
rect 337692 399646 341252 399662
rect 184700 397378 332852 397394
rect 184700 397322 184716 397378
rect 184772 397322 332780 397378
rect 332836 397322 332852 397378
rect 184700 397306 332852 397322
rect 62060 395578 313476 395594
rect 62060 395522 62076 395578
rect 62132 395522 313404 395578
rect 313460 395522 313476 395578
rect 62060 395506 313476 395522
rect 197692 392338 338788 392354
rect 197692 392282 197708 392338
rect 197764 392282 338716 392338
rect 338772 392282 338788 392338
rect 197692 392266 338788 392282
rect 191532 391618 333300 391634
rect 191532 391562 191548 391618
rect 191604 391562 192892 391618
rect 192948 391562 333228 391618
rect 333284 391562 333300 391618
rect 191532 391546 333300 391562
rect 582076 391438 587204 391454
rect 582076 391382 582092 391438
rect 582148 391382 587132 391438
rect 587188 391382 587204 391438
rect 582076 391366 587204 391382
rect 189404 390538 203380 390554
rect 189404 390482 189420 390538
rect 189476 390482 203308 390538
rect 203364 390482 203380 390538
rect 189404 390466 203380 390482
rect 201052 389998 333076 390014
rect 201052 389942 201068 389998
rect 201124 389942 333004 389998
rect 333060 389942 333076 389998
rect 201052 389926 333076 389942
rect 199596 389818 332964 389834
rect 199596 389762 199612 389818
rect 199668 389762 332892 389818
rect 332948 389762 332964 389818
rect 199596 389746 332964 389762
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 359878 388350
rect 359934 388294 360002 388350
rect 360058 388294 390598 388350
rect 390654 388294 390722 388350
rect 390778 388294 421318 388350
rect 421374 388294 421442 388350
rect 421498 388294 452038 388350
rect 452094 388294 452162 388350
rect 452218 388294 482758 388350
rect 482814 388294 482882 388350
rect 482938 388294 513478 388350
rect 513534 388294 513602 388350
rect 513658 388294 544198 388350
rect 544254 388294 544322 388350
rect 544378 388294 574918 388350
rect 574974 388294 575042 388350
rect 575098 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 359878 388226
rect 359934 388170 360002 388226
rect 360058 388170 390598 388226
rect 390654 388170 390722 388226
rect 390778 388170 421318 388226
rect 421374 388170 421442 388226
rect 421498 388170 452038 388226
rect 452094 388170 452162 388226
rect 452218 388170 482758 388226
rect 482814 388170 482882 388226
rect 482938 388170 513478 388226
rect 513534 388170 513602 388226
rect 513658 388170 544198 388226
rect 544254 388170 544322 388226
rect 544378 388170 574918 388226
rect 574974 388170 575042 388226
rect 575098 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 359878 388102
rect 359934 388046 360002 388102
rect 360058 388046 390598 388102
rect 390654 388046 390722 388102
rect 390778 388046 421318 388102
rect 421374 388046 421442 388102
rect 421498 388046 452038 388102
rect 452094 388046 452162 388102
rect 452218 388046 482758 388102
rect 482814 388046 482882 388102
rect 482938 388046 513478 388102
rect 513534 388046 513602 388102
rect 513658 388046 544198 388102
rect 544254 388046 544322 388102
rect 544378 388046 574918 388102
rect 574974 388046 575042 388102
rect 575098 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 359878 387978
rect 359934 387922 360002 387978
rect 360058 387922 390598 387978
rect 390654 387922 390722 387978
rect 390778 387922 421318 387978
rect 421374 387922 421442 387978
rect 421498 387922 452038 387978
rect 452094 387922 452162 387978
rect 452218 387922 482758 387978
rect 482814 387922 482882 387978
rect 482938 387922 513478 387978
rect 513534 387922 513602 387978
rect 513658 387922 544198 387978
rect 544254 387922 544322 387978
rect 544378 387922 574918 387978
rect 574974 387922 575042 387978
rect 575098 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect 202508 387298 317508 387314
rect 202508 387242 202524 387298
rect 202580 387242 317436 387298
rect 317492 387242 317508 387298
rect 202508 387226 317508 387242
rect 197804 386578 331620 386594
rect 197804 386522 197820 386578
rect 197876 386522 331548 386578
rect 331604 386522 331620 386578
rect 197804 386506 331620 386522
rect 202732 384958 336212 384974
rect 202732 384902 202748 384958
rect 202804 384902 336140 384958
rect 336196 384902 336212 384958
rect 202732 384886 336212 384902
rect 20060 384778 334644 384794
rect 20060 384722 20076 384778
rect 20132 384722 334572 384778
rect 334628 384722 334644 384778
rect 20060 384706 334644 384722
rect 18380 383698 331844 383714
rect 18380 383642 18396 383698
rect 18452 383642 331772 383698
rect 331828 383642 331844 383698
rect 18380 383626 331844 383642
rect 203068 383518 335988 383534
rect 203068 383462 203084 383518
rect 203140 383462 335916 383518
rect 335972 383462 335988 383518
rect 203068 383446 335988 383462
rect 14236 383338 214580 383354
rect 14236 383282 14252 383338
rect 14308 383282 214508 383338
rect 214564 383282 214580 383338
rect 14236 383266 214580 383282
rect 200828 383158 216596 383174
rect 200828 383102 200844 383158
rect 200900 383102 216524 383158
rect 216580 383102 216596 383158
rect 200828 383086 216596 383102
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 344518 382350
rect 344574 382294 344642 382350
rect 344698 382294 375238 382350
rect 375294 382294 375362 382350
rect 375418 382294 405958 382350
rect 406014 382294 406082 382350
rect 406138 382294 436678 382350
rect 436734 382294 436802 382350
rect 436858 382294 467398 382350
rect 467454 382294 467522 382350
rect 467578 382294 498118 382350
rect 498174 382294 498242 382350
rect 498298 382294 528838 382350
rect 528894 382294 528962 382350
rect 529018 382294 559558 382350
rect 559614 382294 559682 382350
rect 559738 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 344518 382226
rect 344574 382170 344642 382226
rect 344698 382170 375238 382226
rect 375294 382170 375362 382226
rect 375418 382170 405958 382226
rect 406014 382170 406082 382226
rect 406138 382170 436678 382226
rect 436734 382170 436802 382226
rect 436858 382170 467398 382226
rect 467454 382170 467522 382226
rect 467578 382170 498118 382226
rect 498174 382170 498242 382226
rect 498298 382170 528838 382226
rect 528894 382170 528962 382226
rect 529018 382170 559558 382226
rect 559614 382170 559682 382226
rect 559738 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 344518 382102
rect 344574 382046 344642 382102
rect 344698 382046 375238 382102
rect 375294 382046 375362 382102
rect 375418 382046 405958 382102
rect 406014 382046 406082 382102
rect 406138 382046 436678 382102
rect 436734 382046 436802 382102
rect 436858 382046 467398 382102
rect 467454 382046 467522 382102
rect 467578 382046 498118 382102
rect 498174 382046 498242 382102
rect 498298 382046 528838 382102
rect 528894 382046 528962 382102
rect 529018 382046 559558 382102
rect 559614 382046 559682 382102
rect 559738 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 344518 381978
rect 344574 381922 344642 381978
rect 344698 381922 375238 381978
rect 375294 381922 375362 381978
rect 375418 381922 405958 381978
rect 406014 381922 406082 381978
rect 406138 381922 436678 381978
rect 436734 381922 436802 381978
rect 436858 381922 467398 381978
rect 467454 381922 467522 381978
rect 467578 381922 498118 381978
rect 498174 381922 498242 381978
rect 498298 381922 528838 381978
rect 528894 381922 528962 381978
rect 529018 381922 559558 381978
rect 559614 381922 559682 381978
rect 559738 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect 4044 380278 215924 380294
rect 4044 380222 4060 380278
rect 4116 380222 215852 380278
rect 215908 380222 215924 380278
rect 4044 380206 215924 380222
rect 198140 380098 336324 380114
rect 198140 380042 198156 380098
rect 198212 380042 336252 380098
rect 336308 380042 336324 380098
rect 198140 380026 336324 380042
rect 204860 379918 218612 379934
rect 204860 379862 204876 379918
rect 204932 379862 218540 379918
rect 218596 379862 218612 379918
rect 204860 379846 218612 379862
rect 199148 379738 328484 379754
rect 199148 379682 199164 379738
rect 199220 379682 328412 379738
rect 328468 379682 328484 379738
rect 199148 379666 328484 379682
rect 204636 379378 217268 379394
rect 204636 379322 204652 379378
rect 204708 379322 217196 379378
rect 217252 379322 217268 379378
rect 204636 379306 217268 379322
rect 31036 379198 213236 379214
rect 31036 379142 31052 379198
rect 31108 379142 213164 379198
rect 213220 379142 213236 379198
rect 31036 379126 213236 379142
rect 32716 379018 215252 379034
rect 32716 378962 32732 379018
rect 32788 378962 215180 379018
rect 215236 378962 215252 379018
rect 32716 378946 215252 378962
rect 7516 378838 213908 378854
rect 7516 378782 7532 378838
rect 7588 378782 213836 378838
rect 213892 378782 213908 378838
rect 7516 378766 213908 378782
rect 208276 378118 337780 378134
rect 208276 378062 337708 378118
rect 337764 378062 337780 378118
rect 208276 378046 337780 378062
rect 208276 377954 208364 378046
rect 202620 377938 208364 377954
rect 202620 377882 202636 377938
rect 202692 377882 208364 377938
rect 202620 377866 208364 377882
rect 108316 376498 332740 376514
rect 108316 376442 108332 376498
rect 108388 376442 332668 376498
rect 332724 376442 332740 376498
rect 108316 376426 332740 376442
rect 4156 376318 202596 376334
rect 4156 376262 4172 376318
rect 4228 376262 202524 376318
rect 202580 376262 202596 376318
rect 4156 376246 202596 376262
rect 16700 372178 202708 372194
rect 16700 372122 16716 372178
rect 16772 372122 202636 372178
rect 202692 372122 202708 372178
rect 16700 372106 202708 372122
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 199878 370350
rect 199934 370294 200002 370350
rect 200058 370294 230598 370350
rect 230654 370294 230722 370350
rect 230778 370294 261318 370350
rect 261374 370294 261442 370350
rect 261498 370294 292038 370350
rect 292094 370294 292162 370350
rect 292218 370294 322758 370350
rect 322814 370294 322882 370350
rect 322938 370294 359878 370350
rect 359934 370294 360002 370350
rect 360058 370294 390598 370350
rect 390654 370294 390722 370350
rect 390778 370294 421318 370350
rect 421374 370294 421442 370350
rect 421498 370294 452038 370350
rect 452094 370294 452162 370350
rect 452218 370294 482758 370350
rect 482814 370294 482882 370350
rect 482938 370294 513478 370350
rect 513534 370294 513602 370350
rect 513658 370294 544198 370350
rect 544254 370294 544322 370350
rect 544378 370294 574918 370350
rect 574974 370294 575042 370350
rect 575098 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 199878 370226
rect 199934 370170 200002 370226
rect 200058 370170 230598 370226
rect 230654 370170 230722 370226
rect 230778 370170 261318 370226
rect 261374 370170 261442 370226
rect 261498 370170 292038 370226
rect 292094 370170 292162 370226
rect 292218 370170 322758 370226
rect 322814 370170 322882 370226
rect 322938 370170 359878 370226
rect 359934 370170 360002 370226
rect 360058 370170 390598 370226
rect 390654 370170 390722 370226
rect 390778 370170 421318 370226
rect 421374 370170 421442 370226
rect 421498 370170 452038 370226
rect 452094 370170 452162 370226
rect 452218 370170 482758 370226
rect 482814 370170 482882 370226
rect 482938 370170 513478 370226
rect 513534 370170 513602 370226
rect 513658 370170 544198 370226
rect 544254 370170 544322 370226
rect 544378 370170 574918 370226
rect 574974 370170 575042 370226
rect 575098 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 199878 370102
rect 199934 370046 200002 370102
rect 200058 370046 230598 370102
rect 230654 370046 230722 370102
rect 230778 370046 261318 370102
rect 261374 370046 261442 370102
rect 261498 370046 292038 370102
rect 292094 370046 292162 370102
rect 292218 370046 322758 370102
rect 322814 370046 322882 370102
rect 322938 370046 359878 370102
rect 359934 370046 360002 370102
rect 360058 370046 390598 370102
rect 390654 370046 390722 370102
rect 390778 370046 421318 370102
rect 421374 370046 421442 370102
rect 421498 370046 452038 370102
rect 452094 370046 452162 370102
rect 452218 370046 482758 370102
rect 482814 370046 482882 370102
rect 482938 370046 513478 370102
rect 513534 370046 513602 370102
rect 513658 370046 544198 370102
rect 544254 370046 544322 370102
rect 544378 370046 574918 370102
rect 574974 370046 575042 370102
rect 575098 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 199878 369978
rect 199934 369922 200002 369978
rect 200058 369922 230598 369978
rect 230654 369922 230722 369978
rect 230778 369922 261318 369978
rect 261374 369922 261442 369978
rect 261498 369922 292038 369978
rect 292094 369922 292162 369978
rect 292218 369922 322758 369978
rect 322814 369922 322882 369978
rect 322938 369922 359878 369978
rect 359934 369922 360002 369978
rect 360058 369922 390598 369978
rect 390654 369922 390722 369978
rect 390778 369922 421318 369978
rect 421374 369922 421442 369978
rect 421498 369922 452038 369978
rect 452094 369922 452162 369978
rect 452218 369922 482758 369978
rect 482814 369922 482882 369978
rect 482938 369922 513478 369978
rect 513534 369922 513602 369978
rect 513658 369922 544198 369978
rect 544254 369922 544322 369978
rect 544378 369922 574918 369978
rect 574974 369922 575042 369978
rect 575098 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect 329068 369658 335428 369674
rect 329068 369602 329084 369658
rect 329140 369602 335356 369658
rect 335412 369602 335428 369658
rect 329068 369586 335428 369602
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 184518 364350
rect 184574 364294 184642 364350
rect 184698 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 215238 364350
rect 215294 364294 215362 364350
rect 215418 364294 245958 364350
rect 246014 364294 246082 364350
rect 246138 364294 276678 364350
rect 276734 364294 276802 364350
rect 276858 364294 307398 364350
rect 307454 364294 307522 364350
rect 307578 364294 344518 364350
rect 344574 364294 344642 364350
rect 344698 364294 375238 364350
rect 375294 364294 375362 364350
rect 375418 364294 405958 364350
rect 406014 364294 406082 364350
rect 406138 364294 436678 364350
rect 436734 364294 436802 364350
rect 436858 364294 467398 364350
rect 467454 364294 467522 364350
rect 467578 364294 498118 364350
rect 498174 364294 498242 364350
rect 498298 364294 528838 364350
rect 528894 364294 528962 364350
rect 529018 364294 559558 364350
rect 559614 364294 559682 364350
rect 559738 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 184518 364226
rect 184574 364170 184642 364226
rect 184698 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 215238 364226
rect 215294 364170 215362 364226
rect 215418 364170 245958 364226
rect 246014 364170 246082 364226
rect 246138 364170 276678 364226
rect 276734 364170 276802 364226
rect 276858 364170 307398 364226
rect 307454 364170 307522 364226
rect 307578 364170 344518 364226
rect 344574 364170 344642 364226
rect 344698 364170 375238 364226
rect 375294 364170 375362 364226
rect 375418 364170 405958 364226
rect 406014 364170 406082 364226
rect 406138 364170 436678 364226
rect 436734 364170 436802 364226
rect 436858 364170 467398 364226
rect 467454 364170 467522 364226
rect 467578 364170 498118 364226
rect 498174 364170 498242 364226
rect 498298 364170 528838 364226
rect 528894 364170 528962 364226
rect 529018 364170 559558 364226
rect 559614 364170 559682 364226
rect 559738 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 184518 364102
rect 184574 364046 184642 364102
rect 184698 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 215238 364102
rect 215294 364046 215362 364102
rect 215418 364046 245958 364102
rect 246014 364046 246082 364102
rect 246138 364046 276678 364102
rect 276734 364046 276802 364102
rect 276858 364046 307398 364102
rect 307454 364046 307522 364102
rect 307578 364046 344518 364102
rect 344574 364046 344642 364102
rect 344698 364046 375238 364102
rect 375294 364046 375362 364102
rect 375418 364046 405958 364102
rect 406014 364046 406082 364102
rect 406138 364046 436678 364102
rect 436734 364046 436802 364102
rect 436858 364046 467398 364102
rect 467454 364046 467522 364102
rect 467578 364046 498118 364102
rect 498174 364046 498242 364102
rect 498298 364046 528838 364102
rect 528894 364046 528962 364102
rect 529018 364046 559558 364102
rect 559614 364046 559682 364102
rect 559738 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 184518 363978
rect 184574 363922 184642 363978
rect 184698 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 215238 363978
rect 215294 363922 215362 363978
rect 215418 363922 245958 363978
rect 246014 363922 246082 363978
rect 246138 363922 276678 363978
rect 276734 363922 276802 363978
rect 276858 363922 307398 363978
rect 307454 363922 307522 363978
rect 307578 363922 344518 363978
rect 344574 363922 344642 363978
rect 344698 363922 375238 363978
rect 375294 363922 375362 363978
rect 375418 363922 405958 363978
rect 406014 363922 406082 363978
rect 406138 363922 436678 363978
rect 436734 363922 436802 363978
rect 436858 363922 467398 363978
rect 467454 363922 467522 363978
rect 467578 363922 498118 363978
rect 498174 363922 498242 363978
rect 498298 363922 528838 363978
rect 528894 363922 528962 363978
rect 529018 363922 559558 363978
rect 559614 363922 559682 363978
rect 559738 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect 327388 360838 336436 360854
rect 327388 360782 327404 360838
rect 327460 360782 336364 360838
rect 336420 360782 336436 360838
rect 327388 360766 336436 360782
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 64878 352350
rect 64934 352294 65002 352350
rect 65058 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 134878 352350
rect 134934 352294 135002 352350
rect 135058 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 199878 352350
rect 199934 352294 200002 352350
rect 200058 352294 230598 352350
rect 230654 352294 230722 352350
rect 230778 352294 261318 352350
rect 261374 352294 261442 352350
rect 261498 352294 292038 352350
rect 292094 352294 292162 352350
rect 292218 352294 322758 352350
rect 322814 352294 322882 352350
rect 322938 352294 359878 352350
rect 359934 352294 360002 352350
rect 360058 352294 390598 352350
rect 390654 352294 390722 352350
rect 390778 352294 421318 352350
rect 421374 352294 421442 352350
rect 421498 352294 452038 352350
rect 452094 352294 452162 352350
rect 452218 352294 482758 352350
rect 482814 352294 482882 352350
rect 482938 352294 513478 352350
rect 513534 352294 513602 352350
rect 513658 352294 544198 352350
rect 544254 352294 544322 352350
rect 544378 352294 574918 352350
rect 574974 352294 575042 352350
rect 575098 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 64878 352226
rect 64934 352170 65002 352226
rect 65058 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 134878 352226
rect 134934 352170 135002 352226
rect 135058 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 199878 352226
rect 199934 352170 200002 352226
rect 200058 352170 230598 352226
rect 230654 352170 230722 352226
rect 230778 352170 261318 352226
rect 261374 352170 261442 352226
rect 261498 352170 292038 352226
rect 292094 352170 292162 352226
rect 292218 352170 322758 352226
rect 322814 352170 322882 352226
rect 322938 352170 359878 352226
rect 359934 352170 360002 352226
rect 360058 352170 390598 352226
rect 390654 352170 390722 352226
rect 390778 352170 421318 352226
rect 421374 352170 421442 352226
rect 421498 352170 452038 352226
rect 452094 352170 452162 352226
rect 452218 352170 482758 352226
rect 482814 352170 482882 352226
rect 482938 352170 513478 352226
rect 513534 352170 513602 352226
rect 513658 352170 544198 352226
rect 544254 352170 544322 352226
rect 544378 352170 574918 352226
rect 574974 352170 575042 352226
rect 575098 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 64878 352102
rect 64934 352046 65002 352102
rect 65058 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 134878 352102
rect 134934 352046 135002 352102
rect 135058 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 199878 352102
rect 199934 352046 200002 352102
rect 200058 352046 230598 352102
rect 230654 352046 230722 352102
rect 230778 352046 261318 352102
rect 261374 352046 261442 352102
rect 261498 352046 292038 352102
rect 292094 352046 292162 352102
rect 292218 352046 322758 352102
rect 322814 352046 322882 352102
rect 322938 352046 359878 352102
rect 359934 352046 360002 352102
rect 360058 352046 390598 352102
rect 390654 352046 390722 352102
rect 390778 352046 421318 352102
rect 421374 352046 421442 352102
rect 421498 352046 452038 352102
rect 452094 352046 452162 352102
rect 452218 352046 482758 352102
rect 482814 352046 482882 352102
rect 482938 352046 513478 352102
rect 513534 352046 513602 352102
rect 513658 352046 544198 352102
rect 544254 352046 544322 352102
rect 544378 352046 574918 352102
rect 574974 352046 575042 352102
rect 575098 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 64878 351978
rect 64934 351922 65002 351978
rect 65058 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 134878 351978
rect 134934 351922 135002 351978
rect 135058 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 199878 351978
rect 199934 351922 200002 351978
rect 200058 351922 230598 351978
rect 230654 351922 230722 351978
rect 230778 351922 261318 351978
rect 261374 351922 261442 351978
rect 261498 351922 292038 351978
rect 292094 351922 292162 351978
rect 292218 351922 322758 351978
rect 322814 351922 322882 351978
rect 322938 351922 359878 351978
rect 359934 351922 360002 351978
rect 360058 351922 390598 351978
rect 390654 351922 390722 351978
rect 390778 351922 421318 351978
rect 421374 351922 421442 351978
rect 421498 351922 452038 351978
rect 452094 351922 452162 351978
rect 452218 351922 482758 351978
rect 482814 351922 482882 351978
rect 482938 351922 513478 351978
rect 513534 351922 513602 351978
rect 513658 351922 544198 351978
rect 544254 351922 544322 351978
rect 544378 351922 574918 351978
rect 574974 351922 575042 351978
rect 575098 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect 201052 351118 201700 351134
rect 201052 351062 201068 351118
rect 201124 351062 201628 351118
rect 201684 351062 201700 351118
rect 201052 351046 201700 351062
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 49518 346350
rect 49574 346294 49642 346350
rect 49698 346294 80238 346350
rect 80294 346294 80362 346350
rect 80418 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 119518 346350
rect 119574 346294 119642 346350
rect 119698 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 150238 346350
rect 150294 346294 150362 346350
rect 150418 346294 184518 346350
rect 184574 346294 184642 346350
rect 184698 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 215238 346350
rect 215294 346294 215362 346350
rect 215418 346294 245958 346350
rect 246014 346294 246082 346350
rect 246138 346294 276678 346350
rect 276734 346294 276802 346350
rect 276858 346294 307398 346350
rect 307454 346294 307522 346350
rect 307578 346294 344518 346350
rect 344574 346294 344642 346350
rect 344698 346294 375238 346350
rect 375294 346294 375362 346350
rect 375418 346294 405958 346350
rect 406014 346294 406082 346350
rect 406138 346294 436678 346350
rect 436734 346294 436802 346350
rect 436858 346294 467398 346350
rect 467454 346294 467522 346350
rect 467578 346294 498118 346350
rect 498174 346294 498242 346350
rect 498298 346294 528838 346350
rect 528894 346294 528962 346350
rect 529018 346294 559558 346350
rect 559614 346294 559682 346350
rect 559738 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 49518 346226
rect 49574 346170 49642 346226
rect 49698 346170 80238 346226
rect 80294 346170 80362 346226
rect 80418 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 119518 346226
rect 119574 346170 119642 346226
rect 119698 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 150238 346226
rect 150294 346170 150362 346226
rect 150418 346170 184518 346226
rect 184574 346170 184642 346226
rect 184698 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 215238 346226
rect 215294 346170 215362 346226
rect 215418 346170 245958 346226
rect 246014 346170 246082 346226
rect 246138 346170 276678 346226
rect 276734 346170 276802 346226
rect 276858 346170 307398 346226
rect 307454 346170 307522 346226
rect 307578 346170 344518 346226
rect 344574 346170 344642 346226
rect 344698 346170 375238 346226
rect 375294 346170 375362 346226
rect 375418 346170 405958 346226
rect 406014 346170 406082 346226
rect 406138 346170 436678 346226
rect 436734 346170 436802 346226
rect 436858 346170 467398 346226
rect 467454 346170 467522 346226
rect 467578 346170 498118 346226
rect 498174 346170 498242 346226
rect 498298 346170 528838 346226
rect 528894 346170 528962 346226
rect 529018 346170 559558 346226
rect 559614 346170 559682 346226
rect 559738 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 49518 346102
rect 49574 346046 49642 346102
rect 49698 346046 80238 346102
rect 80294 346046 80362 346102
rect 80418 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 119518 346102
rect 119574 346046 119642 346102
rect 119698 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 150238 346102
rect 150294 346046 150362 346102
rect 150418 346046 184518 346102
rect 184574 346046 184642 346102
rect 184698 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 215238 346102
rect 215294 346046 215362 346102
rect 215418 346046 245958 346102
rect 246014 346046 246082 346102
rect 246138 346046 276678 346102
rect 276734 346046 276802 346102
rect 276858 346046 307398 346102
rect 307454 346046 307522 346102
rect 307578 346046 344518 346102
rect 344574 346046 344642 346102
rect 344698 346046 375238 346102
rect 375294 346046 375362 346102
rect 375418 346046 405958 346102
rect 406014 346046 406082 346102
rect 406138 346046 436678 346102
rect 436734 346046 436802 346102
rect 436858 346046 467398 346102
rect 467454 346046 467522 346102
rect 467578 346046 498118 346102
rect 498174 346046 498242 346102
rect 498298 346046 528838 346102
rect 528894 346046 528962 346102
rect 529018 346046 559558 346102
rect 559614 346046 559682 346102
rect 559738 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 49518 345978
rect 49574 345922 49642 345978
rect 49698 345922 80238 345978
rect 80294 345922 80362 345978
rect 80418 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 119518 345978
rect 119574 345922 119642 345978
rect 119698 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 150238 345978
rect 150294 345922 150362 345978
rect 150418 345922 184518 345978
rect 184574 345922 184642 345978
rect 184698 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 215238 345978
rect 215294 345922 215362 345978
rect 215418 345922 245958 345978
rect 246014 345922 246082 345978
rect 246138 345922 276678 345978
rect 276734 345922 276802 345978
rect 276858 345922 307398 345978
rect 307454 345922 307522 345978
rect 307578 345922 344518 345978
rect 344574 345922 344642 345978
rect 344698 345922 375238 345978
rect 375294 345922 375362 345978
rect 375418 345922 405958 345978
rect 406014 345922 406082 345978
rect 406138 345922 436678 345978
rect 436734 345922 436802 345978
rect 436858 345922 467398 345978
rect 467454 345922 467522 345978
rect 467578 345922 498118 345978
rect 498174 345922 498242 345978
rect 498298 345922 528838 345978
rect 528894 345922 528962 345978
rect 529018 345922 559558 345978
rect 559614 345922 559682 345978
rect 559738 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 64878 334350
rect 64934 334294 65002 334350
rect 65058 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 134878 334350
rect 134934 334294 135002 334350
rect 135058 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 199878 334350
rect 199934 334294 200002 334350
rect 200058 334294 230598 334350
rect 230654 334294 230722 334350
rect 230778 334294 261318 334350
rect 261374 334294 261442 334350
rect 261498 334294 292038 334350
rect 292094 334294 292162 334350
rect 292218 334294 322758 334350
rect 322814 334294 322882 334350
rect 322938 334294 359878 334350
rect 359934 334294 360002 334350
rect 360058 334294 390598 334350
rect 390654 334294 390722 334350
rect 390778 334294 421318 334350
rect 421374 334294 421442 334350
rect 421498 334294 452038 334350
rect 452094 334294 452162 334350
rect 452218 334294 482758 334350
rect 482814 334294 482882 334350
rect 482938 334294 513478 334350
rect 513534 334294 513602 334350
rect 513658 334294 544198 334350
rect 544254 334294 544322 334350
rect 544378 334294 574918 334350
rect 574974 334294 575042 334350
rect 575098 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 64878 334226
rect 64934 334170 65002 334226
rect 65058 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 134878 334226
rect 134934 334170 135002 334226
rect 135058 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 199878 334226
rect 199934 334170 200002 334226
rect 200058 334170 230598 334226
rect 230654 334170 230722 334226
rect 230778 334170 261318 334226
rect 261374 334170 261442 334226
rect 261498 334170 292038 334226
rect 292094 334170 292162 334226
rect 292218 334170 322758 334226
rect 322814 334170 322882 334226
rect 322938 334170 359878 334226
rect 359934 334170 360002 334226
rect 360058 334170 390598 334226
rect 390654 334170 390722 334226
rect 390778 334170 421318 334226
rect 421374 334170 421442 334226
rect 421498 334170 452038 334226
rect 452094 334170 452162 334226
rect 452218 334170 482758 334226
rect 482814 334170 482882 334226
rect 482938 334170 513478 334226
rect 513534 334170 513602 334226
rect 513658 334170 544198 334226
rect 544254 334170 544322 334226
rect 544378 334170 574918 334226
rect 574974 334170 575042 334226
rect 575098 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 64878 334102
rect 64934 334046 65002 334102
rect 65058 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 134878 334102
rect 134934 334046 135002 334102
rect 135058 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 199878 334102
rect 199934 334046 200002 334102
rect 200058 334046 230598 334102
rect 230654 334046 230722 334102
rect 230778 334046 261318 334102
rect 261374 334046 261442 334102
rect 261498 334046 292038 334102
rect 292094 334046 292162 334102
rect 292218 334046 322758 334102
rect 322814 334046 322882 334102
rect 322938 334046 359878 334102
rect 359934 334046 360002 334102
rect 360058 334046 390598 334102
rect 390654 334046 390722 334102
rect 390778 334046 421318 334102
rect 421374 334046 421442 334102
rect 421498 334046 452038 334102
rect 452094 334046 452162 334102
rect 452218 334046 482758 334102
rect 482814 334046 482882 334102
rect 482938 334046 513478 334102
rect 513534 334046 513602 334102
rect 513658 334046 544198 334102
rect 544254 334046 544322 334102
rect 544378 334046 574918 334102
rect 574974 334046 575042 334102
rect 575098 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 64878 333978
rect 64934 333922 65002 333978
rect 65058 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 134878 333978
rect 134934 333922 135002 333978
rect 135058 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 199878 333978
rect 199934 333922 200002 333978
rect 200058 333922 230598 333978
rect 230654 333922 230722 333978
rect 230778 333922 261318 333978
rect 261374 333922 261442 333978
rect 261498 333922 292038 333978
rect 292094 333922 292162 333978
rect 292218 333922 322758 333978
rect 322814 333922 322882 333978
rect 322938 333922 359878 333978
rect 359934 333922 360002 333978
rect 360058 333922 390598 333978
rect 390654 333922 390722 333978
rect 390778 333922 421318 333978
rect 421374 333922 421442 333978
rect 421498 333922 452038 333978
rect 452094 333922 452162 333978
rect 452218 333922 482758 333978
rect 482814 333922 482882 333978
rect 482938 333922 513478 333978
rect 513534 333922 513602 333978
rect 513658 333922 544198 333978
rect 544254 333922 544322 333978
rect 544378 333922 574918 333978
rect 574974 333922 575042 333978
rect 575098 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 49518 328350
rect 49574 328294 49642 328350
rect 49698 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 80238 328350
rect 80294 328294 80362 328350
rect 80418 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 119518 328350
rect 119574 328294 119642 328350
rect 119698 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 150238 328350
rect 150294 328294 150362 328350
rect 150418 328294 184518 328350
rect 184574 328294 184642 328350
rect 184698 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 215238 328350
rect 215294 328294 215362 328350
rect 215418 328294 245958 328350
rect 246014 328294 246082 328350
rect 246138 328294 276678 328350
rect 276734 328294 276802 328350
rect 276858 328294 307398 328350
rect 307454 328294 307522 328350
rect 307578 328294 344518 328350
rect 344574 328294 344642 328350
rect 344698 328294 375238 328350
rect 375294 328294 375362 328350
rect 375418 328294 405958 328350
rect 406014 328294 406082 328350
rect 406138 328294 436678 328350
rect 436734 328294 436802 328350
rect 436858 328294 467398 328350
rect 467454 328294 467522 328350
rect 467578 328294 498118 328350
rect 498174 328294 498242 328350
rect 498298 328294 528838 328350
rect 528894 328294 528962 328350
rect 529018 328294 559558 328350
rect 559614 328294 559682 328350
rect 559738 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 49518 328226
rect 49574 328170 49642 328226
rect 49698 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 80238 328226
rect 80294 328170 80362 328226
rect 80418 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 119518 328226
rect 119574 328170 119642 328226
rect 119698 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 150238 328226
rect 150294 328170 150362 328226
rect 150418 328170 184518 328226
rect 184574 328170 184642 328226
rect 184698 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 215238 328226
rect 215294 328170 215362 328226
rect 215418 328170 245958 328226
rect 246014 328170 246082 328226
rect 246138 328170 276678 328226
rect 276734 328170 276802 328226
rect 276858 328170 307398 328226
rect 307454 328170 307522 328226
rect 307578 328170 344518 328226
rect 344574 328170 344642 328226
rect 344698 328170 375238 328226
rect 375294 328170 375362 328226
rect 375418 328170 405958 328226
rect 406014 328170 406082 328226
rect 406138 328170 436678 328226
rect 436734 328170 436802 328226
rect 436858 328170 467398 328226
rect 467454 328170 467522 328226
rect 467578 328170 498118 328226
rect 498174 328170 498242 328226
rect 498298 328170 528838 328226
rect 528894 328170 528962 328226
rect 529018 328170 559558 328226
rect 559614 328170 559682 328226
rect 559738 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 49518 328102
rect 49574 328046 49642 328102
rect 49698 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 80238 328102
rect 80294 328046 80362 328102
rect 80418 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 119518 328102
rect 119574 328046 119642 328102
rect 119698 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 150238 328102
rect 150294 328046 150362 328102
rect 150418 328046 184518 328102
rect 184574 328046 184642 328102
rect 184698 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 215238 328102
rect 215294 328046 215362 328102
rect 215418 328046 245958 328102
rect 246014 328046 246082 328102
rect 246138 328046 276678 328102
rect 276734 328046 276802 328102
rect 276858 328046 307398 328102
rect 307454 328046 307522 328102
rect 307578 328046 344518 328102
rect 344574 328046 344642 328102
rect 344698 328046 375238 328102
rect 375294 328046 375362 328102
rect 375418 328046 405958 328102
rect 406014 328046 406082 328102
rect 406138 328046 436678 328102
rect 436734 328046 436802 328102
rect 436858 328046 467398 328102
rect 467454 328046 467522 328102
rect 467578 328046 498118 328102
rect 498174 328046 498242 328102
rect 498298 328046 528838 328102
rect 528894 328046 528962 328102
rect 529018 328046 559558 328102
rect 559614 328046 559682 328102
rect 559738 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 49518 327978
rect 49574 327922 49642 327978
rect 49698 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 80238 327978
rect 80294 327922 80362 327978
rect 80418 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 119518 327978
rect 119574 327922 119642 327978
rect 119698 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 150238 327978
rect 150294 327922 150362 327978
rect 150418 327922 184518 327978
rect 184574 327922 184642 327978
rect 184698 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 215238 327978
rect 215294 327922 215362 327978
rect 215418 327922 245958 327978
rect 246014 327922 246082 327978
rect 246138 327922 276678 327978
rect 276734 327922 276802 327978
rect 276858 327922 307398 327978
rect 307454 327922 307522 327978
rect 307578 327922 344518 327978
rect 344574 327922 344642 327978
rect 344698 327922 375238 327978
rect 375294 327922 375362 327978
rect 375418 327922 405958 327978
rect 406014 327922 406082 327978
rect 406138 327922 436678 327978
rect 436734 327922 436802 327978
rect 436858 327922 467398 327978
rect 467454 327922 467522 327978
rect 467578 327922 498118 327978
rect 498174 327922 498242 327978
rect 498298 327922 528838 327978
rect 528894 327922 528962 327978
rect 529018 327922 559558 327978
rect 559614 327922 559682 327978
rect 559738 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect 328620 321058 329380 321074
rect 328620 321002 328636 321058
rect 328692 321002 329308 321058
rect 329364 321002 329380 321058
rect 328620 320986 329380 321002
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 199878 316350
rect 199934 316294 200002 316350
rect 200058 316294 230598 316350
rect 230654 316294 230722 316350
rect 230778 316294 261318 316350
rect 261374 316294 261442 316350
rect 261498 316294 292038 316350
rect 292094 316294 292162 316350
rect 292218 316294 322758 316350
rect 322814 316294 322882 316350
rect 322938 316294 359878 316350
rect 359934 316294 360002 316350
rect 360058 316294 390598 316350
rect 390654 316294 390722 316350
rect 390778 316294 421318 316350
rect 421374 316294 421442 316350
rect 421498 316294 452038 316350
rect 452094 316294 452162 316350
rect 452218 316294 482758 316350
rect 482814 316294 482882 316350
rect 482938 316294 513478 316350
rect 513534 316294 513602 316350
rect 513658 316294 544198 316350
rect 544254 316294 544322 316350
rect 544378 316294 574918 316350
rect 574974 316294 575042 316350
rect 575098 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 199878 316226
rect 199934 316170 200002 316226
rect 200058 316170 230598 316226
rect 230654 316170 230722 316226
rect 230778 316170 261318 316226
rect 261374 316170 261442 316226
rect 261498 316170 292038 316226
rect 292094 316170 292162 316226
rect 292218 316170 322758 316226
rect 322814 316170 322882 316226
rect 322938 316170 359878 316226
rect 359934 316170 360002 316226
rect 360058 316170 390598 316226
rect 390654 316170 390722 316226
rect 390778 316170 421318 316226
rect 421374 316170 421442 316226
rect 421498 316170 452038 316226
rect 452094 316170 452162 316226
rect 452218 316170 482758 316226
rect 482814 316170 482882 316226
rect 482938 316170 513478 316226
rect 513534 316170 513602 316226
rect 513658 316170 544198 316226
rect 544254 316170 544322 316226
rect 544378 316170 574918 316226
rect 574974 316170 575042 316226
rect 575098 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 199878 316102
rect 199934 316046 200002 316102
rect 200058 316046 230598 316102
rect 230654 316046 230722 316102
rect 230778 316046 261318 316102
rect 261374 316046 261442 316102
rect 261498 316046 292038 316102
rect 292094 316046 292162 316102
rect 292218 316046 322758 316102
rect 322814 316046 322882 316102
rect 322938 316046 359878 316102
rect 359934 316046 360002 316102
rect 360058 316046 390598 316102
rect 390654 316046 390722 316102
rect 390778 316046 421318 316102
rect 421374 316046 421442 316102
rect 421498 316046 452038 316102
rect 452094 316046 452162 316102
rect 452218 316046 482758 316102
rect 482814 316046 482882 316102
rect 482938 316046 513478 316102
rect 513534 316046 513602 316102
rect 513658 316046 544198 316102
rect 544254 316046 544322 316102
rect 544378 316046 574918 316102
rect 574974 316046 575042 316102
rect 575098 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 199878 315978
rect 199934 315922 200002 315978
rect 200058 315922 230598 315978
rect 230654 315922 230722 315978
rect 230778 315922 261318 315978
rect 261374 315922 261442 315978
rect 261498 315922 292038 315978
rect 292094 315922 292162 315978
rect 292218 315922 322758 315978
rect 322814 315922 322882 315978
rect 322938 315922 359878 315978
rect 359934 315922 360002 315978
rect 360058 315922 390598 315978
rect 390654 315922 390722 315978
rect 390778 315922 421318 315978
rect 421374 315922 421442 315978
rect 421498 315922 452038 315978
rect 452094 315922 452162 315978
rect 452218 315922 482758 315978
rect 482814 315922 482882 315978
rect 482938 315922 513478 315978
rect 513534 315922 513602 315978
rect 513658 315922 544198 315978
rect 544254 315922 544322 315978
rect 544378 315922 574918 315978
rect 574974 315922 575042 315978
rect 575098 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect 328508 313318 336996 313334
rect 328508 313262 328524 313318
rect 328580 313262 336924 313318
rect 336980 313262 336996 313318
rect 328508 313246 336996 313262
rect 328508 313138 329380 313154
rect 328508 313082 328524 313138
rect 328580 313082 329308 313138
rect 329364 313082 329380 313138
rect 328508 313066 329380 313082
rect 328060 311698 338116 311714
rect 328060 311642 328076 311698
rect 328132 311642 338044 311698
rect 338100 311642 338116 311698
rect 328060 311626 338116 311642
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 184518 310350
rect 184574 310294 184642 310350
rect 184698 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 215238 310350
rect 215294 310294 215362 310350
rect 215418 310294 245958 310350
rect 246014 310294 246082 310350
rect 246138 310294 276678 310350
rect 276734 310294 276802 310350
rect 276858 310294 307398 310350
rect 307454 310294 307522 310350
rect 307578 310294 344518 310350
rect 344574 310294 344642 310350
rect 344698 310294 375238 310350
rect 375294 310294 375362 310350
rect 375418 310294 405958 310350
rect 406014 310294 406082 310350
rect 406138 310294 436678 310350
rect 436734 310294 436802 310350
rect 436858 310294 467398 310350
rect 467454 310294 467522 310350
rect 467578 310294 498118 310350
rect 498174 310294 498242 310350
rect 498298 310294 528838 310350
rect 528894 310294 528962 310350
rect 529018 310294 559558 310350
rect 559614 310294 559682 310350
rect 559738 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 184518 310226
rect 184574 310170 184642 310226
rect 184698 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 215238 310226
rect 215294 310170 215362 310226
rect 215418 310170 245958 310226
rect 246014 310170 246082 310226
rect 246138 310170 276678 310226
rect 276734 310170 276802 310226
rect 276858 310170 307398 310226
rect 307454 310170 307522 310226
rect 307578 310170 344518 310226
rect 344574 310170 344642 310226
rect 344698 310170 375238 310226
rect 375294 310170 375362 310226
rect 375418 310170 405958 310226
rect 406014 310170 406082 310226
rect 406138 310170 436678 310226
rect 436734 310170 436802 310226
rect 436858 310170 467398 310226
rect 467454 310170 467522 310226
rect 467578 310170 498118 310226
rect 498174 310170 498242 310226
rect 498298 310170 528838 310226
rect 528894 310170 528962 310226
rect 529018 310170 559558 310226
rect 559614 310170 559682 310226
rect 559738 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 184518 310102
rect 184574 310046 184642 310102
rect 184698 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 215238 310102
rect 215294 310046 215362 310102
rect 215418 310046 245958 310102
rect 246014 310046 246082 310102
rect 246138 310046 276678 310102
rect 276734 310046 276802 310102
rect 276858 310046 307398 310102
rect 307454 310046 307522 310102
rect 307578 310046 344518 310102
rect 344574 310046 344642 310102
rect 344698 310046 375238 310102
rect 375294 310046 375362 310102
rect 375418 310046 405958 310102
rect 406014 310046 406082 310102
rect 406138 310046 436678 310102
rect 436734 310046 436802 310102
rect 436858 310046 467398 310102
rect 467454 310046 467522 310102
rect 467578 310046 498118 310102
rect 498174 310046 498242 310102
rect 498298 310046 528838 310102
rect 528894 310046 528962 310102
rect 529018 310046 559558 310102
rect 559614 310046 559682 310102
rect 559738 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 184518 309978
rect 184574 309922 184642 309978
rect 184698 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 215238 309978
rect 215294 309922 215362 309978
rect 215418 309922 245958 309978
rect 246014 309922 246082 309978
rect 246138 309922 276678 309978
rect 276734 309922 276802 309978
rect 276858 309922 307398 309978
rect 307454 309922 307522 309978
rect 307578 309922 344518 309978
rect 344574 309922 344642 309978
rect 344698 309922 375238 309978
rect 375294 309922 375362 309978
rect 375418 309922 405958 309978
rect 406014 309922 406082 309978
rect 406138 309922 436678 309978
rect 436734 309922 436802 309978
rect 436858 309922 467398 309978
rect 467454 309922 467522 309978
rect 467578 309922 498118 309978
rect 498174 309922 498242 309978
rect 498298 309922 528838 309978
rect 528894 309922 528962 309978
rect 529018 309922 559558 309978
rect 559614 309922 559682 309978
rect 559738 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect 328844 308278 330052 308294
rect 328844 308222 328860 308278
rect 328916 308222 329980 308278
rect 330036 308222 330052 308278
rect 328844 308206 330052 308222
rect 201052 307378 202484 307394
rect 201052 307322 201068 307378
rect 201124 307322 202412 307378
rect 202468 307322 202484 307378
rect 201052 307306 202484 307322
rect 85580 305938 201140 305954
rect 85580 305882 85596 305938
rect 85652 305882 201068 305938
rect 201124 305882 201140 305938
rect 85580 305866 201140 305882
rect 72140 302518 204164 302534
rect 72140 302462 72156 302518
rect 72212 302462 204092 302518
rect 204148 302462 204164 302518
rect 72140 302446 204164 302462
rect 331756 301618 341140 301634
rect 331756 301562 331772 301618
rect 331828 301562 341068 301618
rect 341124 301562 341140 301618
rect 331756 301546 341140 301562
rect 201164 300898 201812 300914
rect 201164 300842 201180 300898
rect 201236 300842 201740 300898
rect 201796 300842 201812 300898
rect 201164 300826 201812 300842
rect 329068 300898 336100 300914
rect 329068 300842 329084 300898
rect 329140 300842 336028 300898
rect 336084 300842 336100 300898
rect 329068 300826 336100 300842
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 199878 298350
rect 199934 298294 200002 298350
rect 200058 298294 230598 298350
rect 230654 298294 230722 298350
rect 230778 298294 261318 298350
rect 261374 298294 261442 298350
rect 261498 298294 292038 298350
rect 292094 298294 292162 298350
rect 292218 298294 322758 298350
rect 322814 298294 322882 298350
rect 322938 298294 359878 298350
rect 359934 298294 360002 298350
rect 360058 298294 390598 298350
rect 390654 298294 390722 298350
rect 390778 298294 421318 298350
rect 421374 298294 421442 298350
rect 421498 298294 452038 298350
rect 452094 298294 452162 298350
rect 452218 298294 482758 298350
rect 482814 298294 482882 298350
rect 482938 298294 513478 298350
rect 513534 298294 513602 298350
rect 513658 298294 544198 298350
rect 544254 298294 544322 298350
rect 544378 298294 574918 298350
rect 574974 298294 575042 298350
rect 575098 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 199878 298226
rect 199934 298170 200002 298226
rect 200058 298170 230598 298226
rect 230654 298170 230722 298226
rect 230778 298170 261318 298226
rect 261374 298170 261442 298226
rect 261498 298170 292038 298226
rect 292094 298170 292162 298226
rect 292218 298170 322758 298226
rect 322814 298170 322882 298226
rect 322938 298170 359878 298226
rect 359934 298170 360002 298226
rect 360058 298170 390598 298226
rect 390654 298170 390722 298226
rect 390778 298170 421318 298226
rect 421374 298170 421442 298226
rect 421498 298170 452038 298226
rect 452094 298170 452162 298226
rect 452218 298170 482758 298226
rect 482814 298170 482882 298226
rect 482938 298170 513478 298226
rect 513534 298170 513602 298226
rect 513658 298170 544198 298226
rect 544254 298170 544322 298226
rect 544378 298170 574918 298226
rect 574974 298170 575042 298226
rect 575098 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 199878 298102
rect 199934 298046 200002 298102
rect 200058 298046 230598 298102
rect 230654 298046 230722 298102
rect 230778 298046 261318 298102
rect 261374 298046 261442 298102
rect 261498 298046 292038 298102
rect 292094 298046 292162 298102
rect 292218 298046 322758 298102
rect 322814 298046 322882 298102
rect 322938 298046 359878 298102
rect 359934 298046 360002 298102
rect 360058 298046 390598 298102
rect 390654 298046 390722 298102
rect 390778 298046 421318 298102
rect 421374 298046 421442 298102
rect 421498 298046 452038 298102
rect 452094 298046 452162 298102
rect 452218 298046 482758 298102
rect 482814 298046 482882 298102
rect 482938 298046 513478 298102
rect 513534 298046 513602 298102
rect 513658 298046 544198 298102
rect 544254 298046 544322 298102
rect 544378 298046 574918 298102
rect 574974 298046 575042 298102
rect 575098 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 199878 297978
rect 199934 297922 200002 297978
rect 200058 297922 230598 297978
rect 230654 297922 230722 297978
rect 230778 297922 261318 297978
rect 261374 297922 261442 297978
rect 261498 297922 292038 297978
rect 292094 297922 292162 297978
rect 292218 297922 322758 297978
rect 322814 297922 322882 297978
rect 322938 297922 359878 297978
rect 359934 297922 360002 297978
rect 360058 297922 390598 297978
rect 390654 297922 390722 297978
rect 390778 297922 421318 297978
rect 421374 297922 421442 297978
rect 421498 297922 452038 297978
rect 452094 297922 452162 297978
rect 452218 297922 482758 297978
rect 482814 297922 482882 297978
rect 482938 297922 513478 297978
rect 513534 297922 513602 297978
rect 513658 297922 544198 297978
rect 544254 297922 544322 297978
rect 544378 297922 574918 297978
rect 574974 297922 575042 297978
rect 575098 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect 328844 296578 330500 296594
rect 328844 296522 328860 296578
rect 328916 296522 330428 296578
rect 330484 296522 330500 296578
rect 328844 296506 330500 296522
rect 340380 294598 341028 294614
rect 340380 294542 340396 294598
rect 340452 294542 340956 294598
rect 341012 294542 341028 294598
rect 340380 294526 341028 294542
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 184518 292350
rect 184574 292294 184642 292350
rect 184698 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 215238 292350
rect 215294 292294 215362 292350
rect 215418 292294 245958 292350
rect 246014 292294 246082 292350
rect 246138 292294 276678 292350
rect 276734 292294 276802 292350
rect 276858 292294 307398 292350
rect 307454 292294 307522 292350
rect 307578 292294 344518 292350
rect 344574 292294 344642 292350
rect 344698 292294 375238 292350
rect 375294 292294 375362 292350
rect 375418 292294 405958 292350
rect 406014 292294 406082 292350
rect 406138 292294 436678 292350
rect 436734 292294 436802 292350
rect 436858 292294 467398 292350
rect 467454 292294 467522 292350
rect 467578 292294 498118 292350
rect 498174 292294 498242 292350
rect 498298 292294 528838 292350
rect 528894 292294 528962 292350
rect 529018 292294 559558 292350
rect 559614 292294 559682 292350
rect 559738 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 184518 292226
rect 184574 292170 184642 292226
rect 184698 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 215238 292226
rect 215294 292170 215362 292226
rect 215418 292170 245958 292226
rect 246014 292170 246082 292226
rect 246138 292170 276678 292226
rect 276734 292170 276802 292226
rect 276858 292170 307398 292226
rect 307454 292170 307522 292226
rect 307578 292170 344518 292226
rect 344574 292170 344642 292226
rect 344698 292170 375238 292226
rect 375294 292170 375362 292226
rect 375418 292170 405958 292226
rect 406014 292170 406082 292226
rect 406138 292170 436678 292226
rect 436734 292170 436802 292226
rect 436858 292170 467398 292226
rect 467454 292170 467522 292226
rect 467578 292170 498118 292226
rect 498174 292170 498242 292226
rect 498298 292170 528838 292226
rect 528894 292170 528962 292226
rect 529018 292170 559558 292226
rect 559614 292170 559682 292226
rect 559738 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 184518 292102
rect 184574 292046 184642 292102
rect 184698 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 215238 292102
rect 215294 292046 215362 292102
rect 215418 292046 245958 292102
rect 246014 292046 246082 292102
rect 246138 292046 276678 292102
rect 276734 292046 276802 292102
rect 276858 292046 307398 292102
rect 307454 292046 307522 292102
rect 307578 292046 344518 292102
rect 344574 292046 344642 292102
rect 344698 292046 375238 292102
rect 375294 292046 375362 292102
rect 375418 292046 405958 292102
rect 406014 292046 406082 292102
rect 406138 292046 436678 292102
rect 436734 292046 436802 292102
rect 436858 292046 467398 292102
rect 467454 292046 467522 292102
rect 467578 292046 498118 292102
rect 498174 292046 498242 292102
rect 498298 292046 528838 292102
rect 528894 292046 528962 292102
rect 529018 292046 559558 292102
rect 559614 292046 559682 292102
rect 559738 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 184518 291978
rect 184574 291922 184642 291978
rect 184698 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 215238 291978
rect 215294 291922 215362 291978
rect 215418 291922 245958 291978
rect 246014 291922 246082 291978
rect 246138 291922 276678 291978
rect 276734 291922 276802 291978
rect 276858 291922 307398 291978
rect 307454 291922 307522 291978
rect 307578 291922 344518 291978
rect 344574 291922 344642 291978
rect 344698 291922 375238 291978
rect 375294 291922 375362 291978
rect 375418 291922 405958 291978
rect 406014 291922 406082 291978
rect 406138 291922 436678 291978
rect 436734 291922 436802 291978
rect 436858 291922 467398 291978
rect 467454 291922 467522 291978
rect 467578 291922 498118 291978
rect 498174 291922 498242 291978
rect 498298 291922 528838 291978
rect 528894 291922 528962 291978
rect 529018 291922 559558 291978
rect 559614 291922 559682 291978
rect 559738 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect 137772 290638 185684 290654
rect 137772 290582 137788 290638
rect 137844 290582 139244 290638
rect 139300 290582 184828 290638
rect 184884 290582 185612 290638
rect 185668 290582 185684 290638
rect 137772 290566 185684 290582
rect 189292 289018 195316 289034
rect 189292 288962 189308 289018
rect 189364 288962 195244 289018
rect 195300 288962 195316 289018
rect 189292 288946 195316 288962
rect 180444 288838 199012 288854
rect 180444 288782 180460 288838
rect 180516 288782 196028 288838
rect 196084 288782 198940 288838
rect 198996 288782 199012 288838
rect 180444 288766 199012 288782
rect 183916 287218 187364 287234
rect 183916 287162 183932 287218
rect 183988 287162 187292 287218
rect 187348 287162 187364 287218
rect 183916 287146 187364 287162
rect 168908 286498 195988 286514
rect 168908 286442 168924 286498
rect 168980 286442 188076 286498
rect 188132 286442 195916 286498
rect 195972 286442 195988 286498
rect 168908 286426 195988 286442
rect 187164 285778 195764 285794
rect 187164 285722 187180 285778
rect 187236 285722 188076 285778
rect 188132 285722 195692 285778
rect 195748 285722 195764 285778
rect 187164 285706 195764 285722
rect 329068 285778 330276 285794
rect 329068 285722 329084 285778
rect 329140 285722 330204 285778
rect 330260 285722 330276 285778
rect 329068 285706 330276 285722
rect 164092 284698 188148 284714
rect 164092 284642 164108 284698
rect 164164 284642 188076 284698
rect 188132 284642 188148 284698
rect 164092 284626 188148 284642
rect 335564 283978 341364 283994
rect 335564 283922 335580 283978
rect 335636 283922 341292 283978
rect 341348 283922 341364 283978
rect 335564 283906 341364 283922
rect 187276 283798 199236 283814
rect 187276 283742 187292 283798
rect 187348 283742 187852 283798
rect 187908 283742 199164 283798
rect 199220 283742 199236 283798
rect 187276 283726 199236 283742
rect 328732 283798 332964 283814
rect 328732 283742 328748 283798
rect 328804 283742 332892 283798
rect 332948 283742 332964 283798
rect 328732 283726 332964 283742
rect 340380 283798 341140 283814
rect 340380 283742 340396 283798
rect 340452 283742 341068 283798
rect 341124 283742 341140 283798
rect 340380 283726 341140 283742
rect 169020 283258 202596 283274
rect 169020 283202 169036 283258
rect 169092 283202 187964 283258
rect 188020 283202 202524 283258
rect 202580 283202 202596 283258
rect 169020 283186 202596 283202
rect 165548 283078 187364 283094
rect 165548 283022 165564 283078
rect 165620 283022 187292 283078
rect 187348 283022 187364 283078
rect 165548 283006 187364 283022
rect 328732 283078 335764 283094
rect 328732 283022 328748 283078
rect 328804 283022 335692 283078
rect 335748 283022 335764 283078
rect 328732 283006 335764 283022
rect 328396 282718 329380 282734
rect 328396 282662 328412 282718
rect 328468 282662 329308 282718
rect 329364 282662 329380 282718
rect 328396 282646 329380 282662
rect 195900 282358 199460 282374
rect 195900 282302 195916 282358
rect 195972 282302 199388 282358
rect 199444 282302 199460 282358
rect 195900 282286 199460 282302
rect 186380 282178 187476 282194
rect 186380 282122 186396 282178
rect 186452 282122 187404 282178
rect 187460 282122 187476 282178
rect 186380 282106 187476 282122
rect 167228 281458 202484 281474
rect 167228 281402 167244 281458
rect 167300 281402 187740 281458
rect 187796 281402 202412 281458
rect 202468 281402 202484 281458
rect 167228 281386 202484 281402
rect 163420 280738 186468 280754
rect 163420 280682 163436 280738
rect 163492 280682 186396 280738
rect 186452 280682 186468 280738
rect 163420 280666 186468 280682
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 142078 280350
rect 142134 280294 142202 280350
rect 142258 280294 147902 280350
rect 147958 280294 148026 280350
rect 148082 280294 153726 280350
rect 153782 280294 153850 280350
rect 153906 280294 159550 280350
rect 159606 280294 159674 280350
rect 159730 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 199878 280350
rect 199934 280294 200002 280350
rect 200058 280294 230598 280350
rect 230654 280294 230722 280350
rect 230778 280294 261318 280350
rect 261374 280294 261442 280350
rect 261498 280294 292038 280350
rect 292094 280294 292162 280350
rect 292218 280294 322758 280350
rect 322814 280294 322882 280350
rect 322938 280294 359878 280350
rect 359934 280294 360002 280350
rect 360058 280294 390598 280350
rect 390654 280294 390722 280350
rect 390778 280294 421318 280350
rect 421374 280294 421442 280350
rect 421498 280294 452038 280350
rect 452094 280294 452162 280350
rect 452218 280294 482758 280350
rect 482814 280294 482882 280350
rect 482938 280294 513478 280350
rect 513534 280294 513602 280350
rect 513658 280294 544198 280350
rect 544254 280294 544322 280350
rect 544378 280294 574918 280350
rect 574974 280294 575042 280350
rect 575098 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 142078 280226
rect 142134 280170 142202 280226
rect 142258 280170 147902 280226
rect 147958 280170 148026 280226
rect 148082 280170 153726 280226
rect 153782 280170 153850 280226
rect 153906 280170 159550 280226
rect 159606 280170 159674 280226
rect 159730 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 199878 280226
rect 199934 280170 200002 280226
rect 200058 280170 230598 280226
rect 230654 280170 230722 280226
rect 230778 280170 261318 280226
rect 261374 280170 261442 280226
rect 261498 280170 292038 280226
rect 292094 280170 292162 280226
rect 292218 280170 322758 280226
rect 322814 280170 322882 280226
rect 322938 280170 359878 280226
rect 359934 280170 360002 280226
rect 360058 280170 390598 280226
rect 390654 280170 390722 280226
rect 390778 280170 421318 280226
rect 421374 280170 421442 280226
rect 421498 280170 452038 280226
rect 452094 280170 452162 280226
rect 452218 280170 482758 280226
rect 482814 280170 482882 280226
rect 482938 280170 513478 280226
rect 513534 280170 513602 280226
rect 513658 280170 544198 280226
rect 544254 280170 544322 280226
rect 544378 280170 574918 280226
rect 574974 280170 575042 280226
rect 575098 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 142078 280102
rect 142134 280046 142202 280102
rect 142258 280046 147902 280102
rect 147958 280046 148026 280102
rect 148082 280046 153726 280102
rect 153782 280046 153850 280102
rect 153906 280046 159550 280102
rect 159606 280046 159674 280102
rect 159730 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 199878 280102
rect 199934 280046 200002 280102
rect 200058 280046 230598 280102
rect 230654 280046 230722 280102
rect 230778 280046 261318 280102
rect 261374 280046 261442 280102
rect 261498 280046 292038 280102
rect 292094 280046 292162 280102
rect 292218 280046 322758 280102
rect 322814 280046 322882 280102
rect 322938 280046 359878 280102
rect 359934 280046 360002 280102
rect 360058 280046 390598 280102
rect 390654 280046 390722 280102
rect 390778 280046 421318 280102
rect 421374 280046 421442 280102
rect 421498 280046 452038 280102
rect 452094 280046 452162 280102
rect 452218 280046 482758 280102
rect 482814 280046 482882 280102
rect 482938 280046 513478 280102
rect 513534 280046 513602 280102
rect 513658 280046 544198 280102
rect 544254 280046 544322 280102
rect 544378 280046 574918 280102
rect 574974 280046 575042 280102
rect 575098 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 142078 279978
rect 142134 279922 142202 279978
rect 142258 279922 147902 279978
rect 147958 279922 148026 279978
rect 148082 279922 153726 279978
rect 153782 279922 153850 279978
rect 153906 279922 159550 279978
rect 159606 279922 159674 279978
rect 159730 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 199878 279978
rect 199934 279922 200002 279978
rect 200058 279922 230598 279978
rect 230654 279922 230722 279978
rect 230778 279922 261318 279978
rect 261374 279922 261442 279978
rect 261498 279922 292038 279978
rect 292094 279922 292162 279978
rect 292218 279922 322758 279978
rect 322814 279922 322882 279978
rect 322938 279922 359878 279978
rect 359934 279922 360002 279978
rect 360058 279922 390598 279978
rect 390654 279922 390722 279978
rect 390778 279922 421318 279978
rect 421374 279922 421442 279978
rect 421498 279922 452038 279978
rect 452094 279922 452162 279978
rect 452218 279922 482758 279978
rect 482814 279922 482882 279978
rect 482938 279922 513478 279978
rect 513534 279922 513602 279978
rect 513658 279922 544198 279978
rect 544254 279922 544322 279978
rect 544378 279922 574918 279978
rect 574974 279922 575042 279978
rect 575098 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect 179884 279658 184004 279674
rect 179884 279602 179900 279658
rect 179956 279602 183932 279658
rect 183988 279602 184004 279658
rect 179884 279586 184004 279602
rect 186268 279658 187700 279674
rect 186268 279602 186284 279658
rect 186340 279602 187628 279658
rect 187684 279602 187700 279658
rect 186268 279586 187700 279602
rect 163868 278938 186356 278954
rect 163868 278882 163884 278938
rect 163940 278882 186284 278938
rect 186340 278882 186356 278938
rect 163868 278866 186356 278882
rect 163980 278038 187588 278054
rect 163980 277982 163996 278038
rect 164052 277982 187516 278038
rect 187572 277982 187588 278038
rect 163980 277966 187588 277982
rect 168460 277318 189156 277334
rect 168460 277262 168476 277318
rect 168532 277262 188076 277318
rect 188132 277262 189084 277318
rect 189140 277262 189156 277318
rect 168460 277246 189156 277262
rect 93980 275698 138756 275714
rect 93980 275642 93996 275698
rect 94052 275642 138684 275698
rect 138740 275642 138756 275698
rect 93980 275626 138756 275642
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 139166 274350
rect 139222 274294 139290 274350
rect 139346 274294 144990 274350
rect 145046 274294 145114 274350
rect 145170 274294 150814 274350
rect 150870 274294 150938 274350
rect 150994 274294 156638 274350
rect 156694 274294 156762 274350
rect 156818 274294 184518 274350
rect 184574 274294 184642 274350
rect 184698 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 215238 274350
rect 215294 274294 215362 274350
rect 215418 274294 245958 274350
rect 246014 274294 246082 274350
rect 246138 274294 276678 274350
rect 276734 274294 276802 274350
rect 276858 274294 307398 274350
rect 307454 274294 307522 274350
rect 307578 274294 344518 274350
rect 344574 274294 344642 274350
rect 344698 274294 375238 274350
rect 375294 274294 375362 274350
rect 375418 274294 405958 274350
rect 406014 274294 406082 274350
rect 406138 274294 436678 274350
rect 436734 274294 436802 274350
rect 436858 274294 467398 274350
rect 467454 274294 467522 274350
rect 467578 274294 498118 274350
rect 498174 274294 498242 274350
rect 498298 274294 528838 274350
rect 528894 274294 528962 274350
rect 529018 274294 559558 274350
rect 559614 274294 559682 274350
rect 559738 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 139166 274226
rect 139222 274170 139290 274226
rect 139346 274170 144990 274226
rect 145046 274170 145114 274226
rect 145170 274170 150814 274226
rect 150870 274170 150938 274226
rect 150994 274170 156638 274226
rect 156694 274170 156762 274226
rect 156818 274170 184518 274226
rect 184574 274170 184642 274226
rect 184698 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 215238 274226
rect 215294 274170 215362 274226
rect 215418 274170 245958 274226
rect 246014 274170 246082 274226
rect 246138 274170 276678 274226
rect 276734 274170 276802 274226
rect 276858 274170 307398 274226
rect 307454 274170 307522 274226
rect 307578 274170 344518 274226
rect 344574 274170 344642 274226
rect 344698 274170 375238 274226
rect 375294 274170 375362 274226
rect 375418 274170 405958 274226
rect 406014 274170 406082 274226
rect 406138 274170 436678 274226
rect 436734 274170 436802 274226
rect 436858 274170 467398 274226
rect 467454 274170 467522 274226
rect 467578 274170 498118 274226
rect 498174 274170 498242 274226
rect 498298 274170 528838 274226
rect 528894 274170 528962 274226
rect 529018 274170 559558 274226
rect 559614 274170 559682 274226
rect 559738 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 139166 274102
rect 139222 274046 139290 274102
rect 139346 274046 144990 274102
rect 145046 274046 145114 274102
rect 145170 274046 150814 274102
rect 150870 274046 150938 274102
rect 150994 274046 156638 274102
rect 156694 274046 156762 274102
rect 156818 274046 184518 274102
rect 184574 274046 184642 274102
rect 184698 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 215238 274102
rect 215294 274046 215362 274102
rect 215418 274046 245958 274102
rect 246014 274046 246082 274102
rect 246138 274046 276678 274102
rect 276734 274046 276802 274102
rect 276858 274046 307398 274102
rect 307454 274046 307522 274102
rect 307578 274046 344518 274102
rect 344574 274046 344642 274102
rect 344698 274046 375238 274102
rect 375294 274046 375362 274102
rect 375418 274046 405958 274102
rect 406014 274046 406082 274102
rect 406138 274046 436678 274102
rect 436734 274046 436802 274102
rect 436858 274046 467398 274102
rect 467454 274046 467522 274102
rect 467578 274046 498118 274102
rect 498174 274046 498242 274102
rect 498298 274046 528838 274102
rect 528894 274046 528962 274102
rect 529018 274046 559558 274102
rect 559614 274046 559682 274102
rect 559738 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 139166 273978
rect 139222 273922 139290 273978
rect 139346 273922 144990 273978
rect 145046 273922 145114 273978
rect 145170 273922 150814 273978
rect 150870 273922 150938 273978
rect 150994 273922 156638 273978
rect 156694 273922 156762 273978
rect 156818 273922 184518 273978
rect 184574 273922 184642 273978
rect 184698 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 215238 273978
rect 215294 273922 215362 273978
rect 215418 273922 245958 273978
rect 246014 273922 246082 273978
rect 246138 273922 276678 273978
rect 276734 273922 276802 273978
rect 276858 273922 307398 273978
rect 307454 273922 307522 273978
rect 307578 273922 344518 273978
rect 344574 273922 344642 273978
rect 344698 273922 375238 273978
rect 375294 273922 375362 273978
rect 375418 273922 405958 273978
rect 406014 273922 406082 273978
rect 406138 273922 436678 273978
rect 436734 273922 436802 273978
rect 436858 273922 467398 273978
rect 467454 273922 467522 273978
rect 467578 273922 498118 273978
rect 498174 273922 498242 273978
rect 498298 273922 528838 273978
rect 528894 273922 528962 273978
rect 529018 273922 559558 273978
rect 559614 273922 559682 273978
rect 559738 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect 329068 272998 330612 273014
rect 329068 272942 329084 272998
rect 329140 272942 330540 272998
rect 330596 272942 330612 272998
rect 329068 272926 330612 272942
rect 93420 270658 138644 270674
rect 93420 270602 93436 270658
rect 93492 270602 138572 270658
rect 138628 270602 138644 270658
rect 93420 270586 138644 270602
rect 201164 265618 201812 265634
rect 201164 265562 201180 265618
rect 201236 265562 201740 265618
rect 201796 265562 201812 265618
rect 201164 265546 201812 265562
rect 180556 265438 200804 265454
rect 180556 265382 180572 265438
rect 180628 265382 200732 265438
rect 200788 265382 200804 265438
rect 180556 265366 200804 265382
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 199878 262350
rect 199934 262294 200002 262350
rect 200058 262294 230598 262350
rect 230654 262294 230722 262350
rect 230778 262294 261318 262350
rect 261374 262294 261442 262350
rect 261498 262294 292038 262350
rect 292094 262294 292162 262350
rect 292218 262294 322758 262350
rect 322814 262294 322882 262350
rect 322938 262294 359878 262350
rect 359934 262294 360002 262350
rect 360058 262294 390598 262350
rect 390654 262294 390722 262350
rect 390778 262294 421318 262350
rect 421374 262294 421442 262350
rect 421498 262294 452038 262350
rect 452094 262294 452162 262350
rect 452218 262294 482758 262350
rect 482814 262294 482882 262350
rect 482938 262294 513478 262350
rect 513534 262294 513602 262350
rect 513658 262294 544198 262350
rect 544254 262294 544322 262350
rect 544378 262294 574918 262350
rect 574974 262294 575042 262350
rect 575098 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 199878 262226
rect 199934 262170 200002 262226
rect 200058 262170 230598 262226
rect 230654 262170 230722 262226
rect 230778 262170 261318 262226
rect 261374 262170 261442 262226
rect 261498 262170 292038 262226
rect 292094 262170 292162 262226
rect 292218 262170 322758 262226
rect 322814 262170 322882 262226
rect 322938 262170 359878 262226
rect 359934 262170 360002 262226
rect 360058 262170 390598 262226
rect 390654 262170 390722 262226
rect 390778 262170 421318 262226
rect 421374 262170 421442 262226
rect 421498 262170 452038 262226
rect 452094 262170 452162 262226
rect 452218 262170 482758 262226
rect 482814 262170 482882 262226
rect 482938 262170 513478 262226
rect 513534 262170 513602 262226
rect 513658 262170 544198 262226
rect 544254 262170 544322 262226
rect 544378 262170 574918 262226
rect 574974 262170 575042 262226
rect 575098 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 199878 262102
rect 199934 262046 200002 262102
rect 200058 262046 230598 262102
rect 230654 262046 230722 262102
rect 230778 262046 261318 262102
rect 261374 262046 261442 262102
rect 261498 262046 292038 262102
rect 292094 262046 292162 262102
rect 292218 262046 322758 262102
rect 322814 262046 322882 262102
rect 322938 262046 359878 262102
rect 359934 262046 360002 262102
rect 360058 262046 390598 262102
rect 390654 262046 390722 262102
rect 390778 262046 421318 262102
rect 421374 262046 421442 262102
rect 421498 262046 452038 262102
rect 452094 262046 452162 262102
rect 452218 262046 482758 262102
rect 482814 262046 482882 262102
rect 482938 262046 513478 262102
rect 513534 262046 513602 262102
rect 513658 262046 544198 262102
rect 544254 262046 544322 262102
rect 544378 262046 574918 262102
rect 574974 262046 575042 262102
rect 575098 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 199878 261978
rect 199934 261922 200002 261978
rect 200058 261922 230598 261978
rect 230654 261922 230722 261978
rect 230778 261922 261318 261978
rect 261374 261922 261442 261978
rect 261498 261922 292038 261978
rect 292094 261922 292162 261978
rect 292218 261922 322758 261978
rect 322814 261922 322882 261978
rect 322938 261922 359878 261978
rect 359934 261922 360002 261978
rect 360058 261922 390598 261978
rect 390654 261922 390722 261978
rect 390778 261922 421318 261978
rect 421374 261922 421442 261978
rect 421498 261922 452038 261978
rect 452094 261922 452162 261978
rect 452218 261922 482758 261978
rect 482814 261922 482882 261978
rect 482938 261922 513478 261978
rect 513534 261922 513602 261978
rect 513658 261922 544198 261978
rect 544254 261922 544322 261978
rect 544378 261922 574918 261978
rect 574974 261922 575042 261978
rect 575098 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect 180668 261118 187476 261134
rect 180668 261062 180684 261118
rect 180740 261062 187404 261118
rect 187460 261062 187476 261118
rect 180668 261046 187476 261062
rect 327948 260398 329492 260414
rect 327948 260342 327964 260398
rect 328020 260342 329420 260398
rect 329476 260342 329492 260398
rect 327948 260326 329492 260342
rect 180668 260038 187700 260054
rect 180668 259982 180684 260038
rect 180740 259982 187628 260038
rect 187684 259982 187700 260038
rect 180668 259966 187700 259982
rect 180668 258958 187364 258974
rect 180668 258902 180684 258958
rect 180740 258902 187292 258958
rect 187348 258902 187364 258958
rect 180668 258886 187364 258902
rect 328396 258598 332740 258614
rect 328396 258542 328412 258598
rect 328468 258542 332668 258598
rect 332724 258542 332740 258598
rect 328396 258526 332740 258542
rect 180556 257158 195876 257174
rect 180556 257102 180572 257158
rect 180628 257102 195804 257158
rect 195860 257102 195876 257158
rect 180556 257086 195876 257102
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 184518 256350
rect 184574 256294 184642 256350
rect 184698 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 215238 256350
rect 215294 256294 215362 256350
rect 215418 256294 245958 256350
rect 246014 256294 246082 256350
rect 246138 256294 276678 256350
rect 276734 256294 276802 256350
rect 276858 256294 307398 256350
rect 307454 256294 307522 256350
rect 307578 256294 344518 256350
rect 344574 256294 344642 256350
rect 344698 256294 375238 256350
rect 375294 256294 375362 256350
rect 375418 256294 405958 256350
rect 406014 256294 406082 256350
rect 406138 256294 436678 256350
rect 436734 256294 436802 256350
rect 436858 256294 467398 256350
rect 467454 256294 467522 256350
rect 467578 256294 498118 256350
rect 498174 256294 498242 256350
rect 498298 256294 528838 256350
rect 528894 256294 528962 256350
rect 529018 256294 559558 256350
rect 559614 256294 559682 256350
rect 559738 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 184518 256226
rect 184574 256170 184642 256226
rect 184698 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 215238 256226
rect 215294 256170 215362 256226
rect 215418 256170 245958 256226
rect 246014 256170 246082 256226
rect 246138 256170 276678 256226
rect 276734 256170 276802 256226
rect 276858 256170 307398 256226
rect 307454 256170 307522 256226
rect 307578 256170 344518 256226
rect 344574 256170 344642 256226
rect 344698 256170 375238 256226
rect 375294 256170 375362 256226
rect 375418 256170 405958 256226
rect 406014 256170 406082 256226
rect 406138 256170 436678 256226
rect 436734 256170 436802 256226
rect 436858 256170 467398 256226
rect 467454 256170 467522 256226
rect 467578 256170 498118 256226
rect 498174 256170 498242 256226
rect 498298 256170 528838 256226
rect 528894 256170 528962 256226
rect 529018 256170 559558 256226
rect 559614 256170 559682 256226
rect 559738 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 184518 256102
rect 184574 256046 184642 256102
rect 184698 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 215238 256102
rect 215294 256046 215362 256102
rect 215418 256046 245958 256102
rect 246014 256046 246082 256102
rect 246138 256046 276678 256102
rect 276734 256046 276802 256102
rect 276858 256046 307398 256102
rect 307454 256046 307522 256102
rect 307578 256046 344518 256102
rect 344574 256046 344642 256102
rect 344698 256046 375238 256102
rect 375294 256046 375362 256102
rect 375418 256046 405958 256102
rect 406014 256046 406082 256102
rect 406138 256046 436678 256102
rect 436734 256046 436802 256102
rect 436858 256046 467398 256102
rect 467454 256046 467522 256102
rect 467578 256046 498118 256102
rect 498174 256046 498242 256102
rect 498298 256046 528838 256102
rect 528894 256046 528962 256102
rect 529018 256046 559558 256102
rect 559614 256046 559682 256102
rect 559738 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 184518 255978
rect 184574 255922 184642 255978
rect 184698 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 215238 255978
rect 215294 255922 215362 255978
rect 215418 255922 245958 255978
rect 246014 255922 246082 255978
rect 246138 255922 276678 255978
rect 276734 255922 276802 255978
rect 276858 255922 307398 255978
rect 307454 255922 307522 255978
rect 307578 255922 344518 255978
rect 344574 255922 344642 255978
rect 344698 255922 375238 255978
rect 375294 255922 375362 255978
rect 375418 255922 405958 255978
rect 406014 255922 406082 255978
rect 406138 255922 436678 255978
rect 436734 255922 436802 255978
rect 436858 255922 467398 255978
rect 467454 255922 467522 255978
rect 467578 255922 498118 255978
rect 498174 255922 498242 255978
rect 498298 255922 528838 255978
rect 528894 255922 528962 255978
rect 529018 255922 559558 255978
rect 559614 255922 559682 255978
rect 559738 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect 199260 253738 200804 253754
rect 199260 253682 199276 253738
rect 199332 253682 200732 253738
rect 200788 253682 200804 253738
rect 199260 253666 200804 253682
rect 329180 253738 329828 253754
rect 329180 253682 329196 253738
rect 329252 253682 329756 253738
rect 329812 253682 329828 253738
rect 329180 253666 329828 253682
rect 180556 252298 199348 252314
rect 180556 252242 180572 252298
rect 180628 252242 199276 252298
rect 199332 252242 199348 252298
rect 180556 252226 199348 252242
rect 180668 252118 202708 252134
rect 180668 252062 180684 252118
rect 180740 252062 202636 252118
rect 202692 252062 202708 252118
rect 180668 252046 202708 252062
rect 328620 249598 330500 249614
rect 328620 249542 328636 249598
rect 328692 249542 330428 249598
rect 330484 249542 330500 249598
rect 328620 249526 330500 249542
rect 328732 249418 338900 249434
rect 328732 249362 328748 249418
rect 328804 249362 338828 249418
rect 338884 249362 338900 249418
rect 328732 249346 338900 249362
rect 328284 249238 332740 249254
rect 328284 249182 328300 249238
rect 328356 249182 332668 249238
rect 332724 249182 332740 249238
rect 328284 249166 332740 249182
rect 329068 248518 331060 248534
rect 329068 248462 329084 248518
rect 329140 248462 330988 248518
rect 331044 248462 331060 248518
rect 329068 248446 331060 248462
rect 328620 248338 331284 248354
rect 328620 248282 328636 248338
rect 328692 248282 331212 248338
rect 331268 248282 331284 248338
rect 328620 248266 331284 248282
rect 327388 248158 330948 248174
rect 327388 248102 327404 248158
rect 327460 248102 330876 248158
rect 330932 248102 330948 248158
rect 327388 248086 330948 248102
rect 329180 247978 333636 247994
rect 329180 247922 329196 247978
rect 329252 247922 333564 247978
rect 333620 247922 333636 247978
rect 329180 247906 333636 247922
rect 4604 247078 42884 247094
rect 4604 247022 4620 247078
rect 4676 247022 42812 247078
rect 42868 247022 42884 247078
rect 4604 247006 42884 247022
rect 195900 246898 199460 246914
rect 195900 246842 195916 246898
rect 195972 246842 199388 246898
rect 199444 246842 199460 246898
rect 195900 246826 199460 246842
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 199878 244350
rect 199934 244294 200002 244350
rect 200058 244294 230598 244350
rect 230654 244294 230722 244350
rect 230778 244294 261318 244350
rect 261374 244294 261442 244350
rect 261498 244294 292038 244350
rect 292094 244294 292162 244350
rect 292218 244294 322758 244350
rect 322814 244294 322882 244350
rect 322938 244294 359878 244350
rect 359934 244294 360002 244350
rect 360058 244294 390598 244350
rect 390654 244294 390722 244350
rect 390778 244294 421318 244350
rect 421374 244294 421442 244350
rect 421498 244294 452038 244350
rect 452094 244294 452162 244350
rect 452218 244294 482758 244350
rect 482814 244294 482882 244350
rect 482938 244294 513478 244350
rect 513534 244294 513602 244350
rect 513658 244294 544198 244350
rect 544254 244294 544322 244350
rect 544378 244294 574918 244350
rect 574974 244294 575042 244350
rect 575098 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 199878 244226
rect 199934 244170 200002 244226
rect 200058 244170 230598 244226
rect 230654 244170 230722 244226
rect 230778 244170 261318 244226
rect 261374 244170 261442 244226
rect 261498 244170 292038 244226
rect 292094 244170 292162 244226
rect 292218 244170 322758 244226
rect 322814 244170 322882 244226
rect 322938 244170 359878 244226
rect 359934 244170 360002 244226
rect 360058 244170 390598 244226
rect 390654 244170 390722 244226
rect 390778 244170 421318 244226
rect 421374 244170 421442 244226
rect 421498 244170 452038 244226
rect 452094 244170 452162 244226
rect 452218 244170 482758 244226
rect 482814 244170 482882 244226
rect 482938 244170 513478 244226
rect 513534 244170 513602 244226
rect 513658 244170 544198 244226
rect 544254 244170 544322 244226
rect 544378 244170 574918 244226
rect 574974 244170 575042 244226
rect 575098 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 199878 244102
rect 199934 244046 200002 244102
rect 200058 244046 230598 244102
rect 230654 244046 230722 244102
rect 230778 244046 261318 244102
rect 261374 244046 261442 244102
rect 261498 244046 292038 244102
rect 292094 244046 292162 244102
rect 292218 244046 322758 244102
rect 322814 244046 322882 244102
rect 322938 244046 359878 244102
rect 359934 244046 360002 244102
rect 360058 244046 390598 244102
rect 390654 244046 390722 244102
rect 390778 244046 421318 244102
rect 421374 244046 421442 244102
rect 421498 244046 452038 244102
rect 452094 244046 452162 244102
rect 452218 244046 482758 244102
rect 482814 244046 482882 244102
rect 482938 244046 513478 244102
rect 513534 244046 513602 244102
rect 513658 244046 544198 244102
rect 544254 244046 544322 244102
rect 544378 244046 574918 244102
rect 574974 244046 575042 244102
rect 575098 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 199878 243978
rect 199934 243922 200002 243978
rect 200058 243922 230598 243978
rect 230654 243922 230722 243978
rect 230778 243922 261318 243978
rect 261374 243922 261442 243978
rect 261498 243922 292038 243978
rect 292094 243922 292162 243978
rect 292218 243922 322758 243978
rect 322814 243922 322882 243978
rect 322938 243922 359878 243978
rect 359934 243922 360002 243978
rect 360058 243922 390598 243978
rect 390654 243922 390722 243978
rect 390778 243922 421318 243978
rect 421374 243922 421442 243978
rect 421498 243922 452038 243978
rect 452094 243922 452162 243978
rect 452218 243922 482758 243978
rect 482814 243922 482882 243978
rect 482938 243922 513478 243978
rect 513534 243922 513602 243978
rect 513658 243922 544198 243978
rect 544254 243922 544322 243978
rect 544378 243922 574918 243978
rect 574974 243922 575042 243978
rect 575098 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect 335116 243478 341140 243494
rect 335116 243422 335132 243478
rect 335188 243422 341068 243478
rect 341124 243422 341140 243478
rect 335116 243406 341140 243422
rect 328732 242218 333188 242234
rect 328732 242162 328748 242218
rect 328804 242162 333116 242218
rect 333172 242162 333188 242218
rect 328732 242146 333188 242162
rect 329068 242038 331732 242054
rect 329068 241982 329084 242038
rect 329140 241982 331660 242038
rect 331716 241982 331732 242038
rect 329068 241966 331732 241982
rect 326716 240958 338452 240974
rect 326716 240902 326732 240958
rect 326788 240902 338380 240958
rect 338436 240902 338452 240958
rect 326716 240886 338452 240902
rect 326604 240778 332404 240794
rect 326604 240722 326620 240778
rect 326676 240722 332332 240778
rect 332388 240722 332404 240778
rect 326604 240706 332404 240722
rect 326828 240598 333412 240614
rect 326828 240542 326844 240598
rect 326900 240542 333340 240598
rect 333396 240542 333412 240598
rect 326828 240526 333412 240542
rect 326940 240418 331172 240434
rect 326940 240362 326956 240418
rect 327012 240362 331100 240418
rect 331156 240362 331172 240418
rect 326940 240346 331172 240362
rect 286396 239518 336324 239534
rect 286396 239462 286412 239518
rect 286468 239462 336252 239518
rect 336308 239462 336324 239518
rect 286396 239446 336324 239462
rect 196236 239338 321764 239354
rect 196236 239282 196252 239338
rect 196308 239282 321692 239338
rect 321748 239282 321764 239338
rect 196236 239266 321764 239282
rect 327612 239338 341364 239354
rect 327612 239282 327628 239338
rect 327684 239282 341292 239338
rect 341348 239282 341364 239338
rect 327612 239266 341364 239282
rect 327052 238618 331620 238634
rect 327052 238562 327068 238618
rect 327124 238562 331548 238618
rect 331604 238562 331620 238618
rect 327052 238546 331620 238562
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 344518 238350
rect 344574 238294 344642 238350
rect 344698 238294 375238 238350
rect 375294 238294 375362 238350
rect 375418 238294 405958 238350
rect 406014 238294 406082 238350
rect 406138 238294 436678 238350
rect 436734 238294 436802 238350
rect 436858 238294 467398 238350
rect 467454 238294 467522 238350
rect 467578 238294 498118 238350
rect 498174 238294 498242 238350
rect 498298 238294 528838 238350
rect 528894 238294 528962 238350
rect 529018 238294 559558 238350
rect 559614 238294 559682 238350
rect 559738 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 344518 238226
rect 344574 238170 344642 238226
rect 344698 238170 375238 238226
rect 375294 238170 375362 238226
rect 375418 238170 405958 238226
rect 406014 238170 406082 238226
rect 406138 238170 436678 238226
rect 436734 238170 436802 238226
rect 436858 238170 467398 238226
rect 467454 238170 467522 238226
rect 467578 238170 498118 238226
rect 498174 238170 498242 238226
rect 498298 238170 528838 238226
rect 528894 238170 528962 238226
rect 529018 238170 559558 238226
rect 559614 238170 559682 238226
rect 559738 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 344518 238102
rect 344574 238046 344642 238102
rect 344698 238046 375238 238102
rect 375294 238046 375362 238102
rect 375418 238046 405958 238102
rect 406014 238046 406082 238102
rect 406138 238046 436678 238102
rect 436734 238046 436802 238102
rect 436858 238046 467398 238102
rect 467454 238046 467522 238102
rect 467578 238046 498118 238102
rect 498174 238046 498242 238102
rect 498298 238046 528838 238102
rect 528894 238046 528962 238102
rect 529018 238046 559558 238102
rect 559614 238046 559682 238102
rect 559738 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 344518 237978
rect 344574 237922 344642 237978
rect 344698 237922 375238 237978
rect 375294 237922 375362 237978
rect 375418 237922 405958 237978
rect 406014 237922 406082 237978
rect 406138 237922 436678 237978
rect 436734 237922 436802 237978
rect 436858 237922 467398 237978
rect 467454 237922 467522 237978
rect 467578 237922 498118 237978
rect 498174 237922 498242 237978
rect 498298 237922 528838 237978
rect 528894 237922 528962 237978
rect 529018 237922 559558 237978
rect 559614 237922 559682 237978
rect 559738 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect 67996 237718 91828 237734
rect 67996 237662 68012 237718
rect 68068 237662 91756 237718
rect 91812 237662 91828 237718
rect 67996 237646 91828 237662
rect 71580 237538 91604 237554
rect 71580 237482 71596 237538
rect 71652 237482 91532 237538
rect 91588 237482 91604 237538
rect 71580 237466 91604 237482
rect 235100 237178 267220 237194
rect 235100 237122 235116 237178
rect 235172 237122 267148 237178
rect 267204 237122 267220 237178
rect 235100 237106 267220 237122
rect 234204 236998 267444 237014
rect 234204 236942 234220 236998
rect 234276 236942 267372 236998
rect 267428 236942 267444 236998
rect 234204 236926 267444 236942
rect 323356 236278 329828 236294
rect 323356 236222 323372 236278
rect 323428 236222 329756 236278
rect 329812 236222 329828 236278
rect 323356 236206 329828 236222
rect 279676 236098 341140 236114
rect 279676 236042 279692 236098
rect 279748 236042 341068 236098
rect 341124 236042 341140 236098
rect 279676 236026 341140 236042
rect 176972 234298 294996 234314
rect 176972 234242 176988 234298
rect 177044 234242 294924 234298
rect 294980 234242 294996 234298
rect 176972 234226 294996 234242
rect 187612 231058 281556 231074
rect 187612 231002 187628 231058
rect 187684 231002 281484 231058
rect 281540 231002 281556 231058
rect 187612 230986 281556 231002
rect 288300 231058 333076 231074
rect 288300 231002 288316 231058
rect 288372 231002 333004 231058
rect 333060 231002 333076 231058
rect 288300 230986 333076 231002
rect 35180 229258 333972 229274
rect 35180 229202 35196 229258
rect 35252 229202 333900 229258
rect 333956 229202 333972 229258
rect 35180 229186 333972 229202
rect 201500 227638 332292 227654
rect 201500 227582 201516 227638
rect 201572 227582 332220 227638
rect 332276 227582 332292 227638
rect 201500 227566 332292 227582
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 359878 226350
rect 359934 226294 360002 226350
rect 360058 226294 390598 226350
rect 390654 226294 390722 226350
rect 390778 226294 421318 226350
rect 421374 226294 421442 226350
rect 421498 226294 452038 226350
rect 452094 226294 452162 226350
rect 452218 226294 482758 226350
rect 482814 226294 482882 226350
rect 482938 226294 513478 226350
rect 513534 226294 513602 226350
rect 513658 226294 544198 226350
rect 544254 226294 544322 226350
rect 544378 226294 574918 226350
rect 574974 226294 575042 226350
rect 575098 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 359878 226226
rect 359934 226170 360002 226226
rect 360058 226170 390598 226226
rect 390654 226170 390722 226226
rect 390778 226170 421318 226226
rect 421374 226170 421442 226226
rect 421498 226170 452038 226226
rect 452094 226170 452162 226226
rect 452218 226170 482758 226226
rect 482814 226170 482882 226226
rect 482938 226170 513478 226226
rect 513534 226170 513602 226226
rect 513658 226170 544198 226226
rect 544254 226170 544322 226226
rect 544378 226170 574918 226226
rect 574974 226170 575042 226226
rect 575098 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 359878 226102
rect 359934 226046 360002 226102
rect 360058 226046 390598 226102
rect 390654 226046 390722 226102
rect 390778 226046 421318 226102
rect 421374 226046 421442 226102
rect 421498 226046 452038 226102
rect 452094 226046 452162 226102
rect 452218 226046 482758 226102
rect 482814 226046 482882 226102
rect 482938 226046 513478 226102
rect 513534 226046 513602 226102
rect 513658 226046 544198 226102
rect 544254 226046 544322 226102
rect 544378 226046 574918 226102
rect 574974 226046 575042 226102
rect 575098 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 359878 225978
rect 359934 225922 360002 225978
rect 360058 225922 390598 225978
rect 390654 225922 390722 225978
rect 390778 225922 421318 225978
rect 421374 225922 421442 225978
rect 421498 225922 452038 225978
rect 452094 225922 452162 225978
rect 452218 225922 482758 225978
rect 482814 225922 482882 225978
rect 482938 225922 513478 225978
rect 513534 225922 513602 225978
rect 513658 225922 544198 225978
rect 544254 225922 544322 225978
rect 544378 225922 574918 225978
rect 574974 225922 575042 225978
rect 575098 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect 201276 224218 292420 224234
rect 201276 224162 201292 224218
rect 201348 224162 292348 224218
rect 292404 224162 292420 224218
rect 201276 224146 292420 224162
rect 200828 222598 271476 222614
rect 200828 222542 200844 222598
rect 200900 222542 271404 222598
rect 271460 222542 271476 222598
rect 200828 222526 271476 222542
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 344518 220350
rect 344574 220294 344642 220350
rect 344698 220294 375238 220350
rect 375294 220294 375362 220350
rect 375418 220294 405958 220350
rect 406014 220294 406082 220350
rect 406138 220294 436678 220350
rect 436734 220294 436802 220350
rect 436858 220294 467398 220350
rect 467454 220294 467522 220350
rect 467578 220294 498118 220350
rect 498174 220294 498242 220350
rect 498298 220294 528838 220350
rect 528894 220294 528962 220350
rect 529018 220294 559558 220350
rect 559614 220294 559682 220350
rect 559738 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 344518 220226
rect 344574 220170 344642 220226
rect 344698 220170 375238 220226
rect 375294 220170 375362 220226
rect 375418 220170 405958 220226
rect 406014 220170 406082 220226
rect 406138 220170 436678 220226
rect 436734 220170 436802 220226
rect 436858 220170 467398 220226
rect 467454 220170 467522 220226
rect 467578 220170 498118 220226
rect 498174 220170 498242 220226
rect 498298 220170 528838 220226
rect 528894 220170 528962 220226
rect 529018 220170 559558 220226
rect 559614 220170 559682 220226
rect 559738 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 344518 220102
rect 344574 220046 344642 220102
rect 344698 220046 375238 220102
rect 375294 220046 375362 220102
rect 375418 220046 405958 220102
rect 406014 220046 406082 220102
rect 406138 220046 436678 220102
rect 436734 220046 436802 220102
rect 436858 220046 467398 220102
rect 467454 220046 467522 220102
rect 467578 220046 498118 220102
rect 498174 220046 498242 220102
rect 498298 220046 528838 220102
rect 528894 220046 528962 220102
rect 529018 220046 559558 220102
rect 559614 220046 559682 220102
rect 559738 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 344518 219978
rect 344574 219922 344642 219978
rect 344698 219922 375238 219978
rect 375294 219922 375362 219978
rect 375418 219922 405958 219978
rect 406014 219922 406082 219978
rect 406138 219922 436678 219978
rect 436734 219922 436802 219978
rect 436858 219922 467398 219978
rect 467454 219922 467522 219978
rect 467578 219922 498118 219978
rect 498174 219922 498242 219978
rect 498298 219922 528838 219978
rect 528894 219922 528962 219978
rect 529018 219922 559558 219978
rect 559614 219922 559682 219978
rect 559738 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect 192652 219178 285252 219194
rect 192652 219122 192668 219178
rect 192724 219122 285180 219178
rect 285236 219122 285252 219178
rect 192652 219106 285252 219122
rect 199596 217558 333524 217574
rect 199596 217502 199612 217558
rect 199668 217502 333452 217558
rect 333508 217502 333524 217558
rect 199596 217486 333524 217502
rect 192092 215938 283236 215954
rect 192092 215882 192108 215938
rect 192164 215882 283164 215938
rect 283220 215882 283236 215938
rect 192092 215866 283236 215882
rect 201388 214138 295108 214154
rect 201388 214082 201404 214138
rect 201460 214082 295036 214138
rect 295092 214082 295108 214138
rect 201388 214066 295108 214082
rect 191308 212518 274836 212534
rect 191308 212462 191324 212518
rect 191380 212462 274764 212518
rect 274820 212462 274836 212518
rect 191308 212446 274836 212462
rect 177532 211798 276404 211814
rect 177532 211742 177548 211798
rect 177604 211742 276332 211798
rect 276388 211742 276404 211798
rect 177532 211726 276404 211742
rect 190748 211078 274724 211094
rect 190748 211022 190764 211078
rect 190820 211022 274652 211078
rect 274708 211022 274724 211078
rect 190748 211006 274724 211022
rect 41788 210898 325348 210914
rect 41788 210842 41804 210898
rect 41860 210842 325276 210898
rect 325332 210842 325348 210898
rect 41788 210826 325348 210842
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 359878 208350
rect 359934 208294 360002 208350
rect 360058 208294 390598 208350
rect 390654 208294 390722 208350
rect 390778 208294 421318 208350
rect 421374 208294 421442 208350
rect 421498 208294 452038 208350
rect 452094 208294 452162 208350
rect 452218 208294 482758 208350
rect 482814 208294 482882 208350
rect 482938 208294 513478 208350
rect 513534 208294 513602 208350
rect 513658 208294 544198 208350
rect 544254 208294 544322 208350
rect 544378 208294 574918 208350
rect 574974 208294 575042 208350
rect 575098 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 359878 208226
rect 359934 208170 360002 208226
rect 360058 208170 390598 208226
rect 390654 208170 390722 208226
rect 390778 208170 421318 208226
rect 421374 208170 421442 208226
rect 421498 208170 452038 208226
rect 452094 208170 452162 208226
rect 452218 208170 482758 208226
rect 482814 208170 482882 208226
rect 482938 208170 513478 208226
rect 513534 208170 513602 208226
rect 513658 208170 544198 208226
rect 544254 208170 544322 208226
rect 544378 208170 574918 208226
rect 574974 208170 575042 208226
rect 575098 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 359878 208102
rect 359934 208046 360002 208102
rect 360058 208046 390598 208102
rect 390654 208046 390722 208102
rect 390778 208046 421318 208102
rect 421374 208046 421442 208102
rect 421498 208046 452038 208102
rect 452094 208046 452162 208102
rect 452218 208046 482758 208102
rect 482814 208046 482882 208102
rect 482938 208046 513478 208102
rect 513534 208046 513602 208102
rect 513658 208046 544198 208102
rect 544254 208046 544322 208102
rect 544378 208046 574918 208102
rect 574974 208046 575042 208102
rect 575098 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 359878 207978
rect 359934 207922 360002 207978
rect 360058 207922 390598 207978
rect 390654 207922 390722 207978
rect 390778 207922 421318 207978
rect 421374 207922 421442 207978
rect 421498 207922 452038 207978
rect 452094 207922 452162 207978
rect 452218 207922 482758 207978
rect 482814 207922 482882 207978
rect 482938 207922 513478 207978
rect 513534 207922 513602 207978
rect 513658 207922 544198 207978
rect 544254 207922 544322 207978
rect 544378 207922 574918 207978
rect 574974 207922 575042 207978
rect 575098 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect 233420 207478 273156 207494
rect 233420 207422 233436 207478
rect 233492 207422 273084 207478
rect 273140 207422 273156 207478
rect 233420 207406 273156 207422
rect 4044 206578 196604 206594
rect 4044 206522 4060 206578
rect 4116 206522 196476 206578
rect 196532 206522 196604 206578
rect 4044 206506 196604 206522
rect 231740 206578 262124 206594
rect 231740 206522 231756 206578
rect 231812 206522 262124 206578
rect 231740 206506 262124 206522
rect 265228 206578 269796 206594
rect 265228 206522 265244 206578
rect 265300 206522 269724 206578
rect 269780 206522 269796 206578
rect 265228 206506 269796 206522
rect 196516 206054 196604 206506
rect 262036 206414 262124 206506
rect 262036 206398 273044 206414
rect 262036 206342 272972 206398
rect 273028 206342 273044 206398
rect 262036 206326 273044 206342
rect 266796 206218 271700 206234
rect 266796 206162 266812 206218
rect 266868 206162 271628 206218
rect 271684 206162 271700 206218
rect 266796 206146 271700 206162
rect 196516 206038 271924 206054
rect 196516 205982 271852 206038
rect 271908 205982 271924 206038
rect 196516 205966 271924 205982
rect 39436 205858 268004 205874
rect 39436 205802 39452 205858
rect 39508 205802 203084 205858
rect 203140 205802 267932 205858
rect 267988 205802 268004 205858
rect 39436 205786 268004 205802
rect 267020 204958 269908 204974
rect 267020 204902 267036 204958
rect 267092 204902 269836 204958
rect 269892 204902 269908 204958
rect 267020 204886 269908 204902
rect 265340 204418 274948 204434
rect 265340 204362 265356 204418
rect 265412 204362 274876 204418
rect 274932 204362 274948 204418
rect 265340 204346 274948 204362
rect 254476 204238 272372 204254
rect 254476 204182 254492 204238
rect 254548 204182 272300 204238
rect 272356 204182 272372 204238
rect 254476 204166 272372 204182
rect 226700 204058 267668 204074
rect 226700 204002 226716 204058
rect 226772 204002 267596 204058
rect 267652 204002 267668 204058
rect 226700 203986 267668 204002
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 344518 202350
rect 344574 202294 344642 202350
rect 344698 202294 375238 202350
rect 375294 202294 375362 202350
rect 375418 202294 405958 202350
rect 406014 202294 406082 202350
rect 406138 202294 436678 202350
rect 436734 202294 436802 202350
rect 436858 202294 467398 202350
rect 467454 202294 467522 202350
rect 467578 202294 498118 202350
rect 498174 202294 498242 202350
rect 498298 202294 528838 202350
rect 528894 202294 528962 202350
rect 529018 202294 559558 202350
rect 559614 202294 559682 202350
rect 559738 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 344518 202226
rect 344574 202170 344642 202226
rect 344698 202170 375238 202226
rect 375294 202170 375362 202226
rect 375418 202170 405958 202226
rect 406014 202170 406082 202226
rect 406138 202170 436678 202226
rect 436734 202170 436802 202226
rect 436858 202170 467398 202226
rect 467454 202170 467522 202226
rect 467578 202170 498118 202226
rect 498174 202170 498242 202226
rect 498298 202170 528838 202226
rect 528894 202170 528962 202226
rect 529018 202170 559558 202226
rect 559614 202170 559682 202226
rect 559738 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 344518 202102
rect 344574 202046 344642 202102
rect 344698 202046 375238 202102
rect 375294 202046 375362 202102
rect 375418 202046 405958 202102
rect 406014 202046 406082 202102
rect 406138 202046 436678 202102
rect 436734 202046 436802 202102
rect 436858 202046 467398 202102
rect 467454 202046 467522 202102
rect 467578 202046 498118 202102
rect 498174 202046 498242 202102
rect 498298 202046 528838 202102
rect 528894 202046 528962 202102
rect 529018 202046 559558 202102
rect 559614 202046 559682 202102
rect 559738 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 344518 201978
rect 344574 201922 344642 201978
rect 344698 201922 375238 201978
rect 375294 201922 375362 201978
rect 375418 201922 405958 201978
rect 406014 201922 406082 201978
rect 406138 201922 436678 201978
rect 436734 201922 436802 201978
rect 436858 201922 467398 201978
rect 467454 201922 467522 201978
rect 467578 201922 498118 201978
rect 498174 201922 498242 201978
rect 498298 201922 528838 201978
rect 528894 201922 528962 201978
rect 529018 201922 559558 201978
rect 559614 201922 559682 201978
rect 559738 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect 268028 201538 269684 201554
rect 268028 201482 268044 201538
rect 268100 201482 269612 201538
rect 269668 201482 269684 201538
rect 268028 201466 269684 201482
rect 298940 199018 326916 199034
rect 298940 198962 298956 199018
rect 299012 198962 326844 199018
rect 326900 198962 326916 199018
rect 298940 198946 326916 198962
rect 321676 197398 337108 197414
rect 321676 197342 321692 197398
rect 321748 197342 337036 197398
rect 337092 197342 337108 197398
rect 321676 197326 337108 197342
rect 323132 191458 336100 191474
rect 323132 191402 323148 191458
rect 323204 191402 336028 191458
rect 336084 191402 336100 191458
rect 323132 191386 336100 191402
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 295578 190350
rect 295634 190294 295702 190350
rect 295758 190294 304902 190350
rect 304958 190294 305026 190350
rect 305082 190294 314226 190350
rect 314282 190294 314350 190350
rect 314406 190294 323550 190350
rect 323606 190294 323674 190350
rect 323730 190294 359878 190350
rect 359934 190294 360002 190350
rect 360058 190294 390598 190350
rect 390654 190294 390722 190350
rect 390778 190294 421318 190350
rect 421374 190294 421442 190350
rect 421498 190294 452038 190350
rect 452094 190294 452162 190350
rect 452218 190294 482758 190350
rect 482814 190294 482882 190350
rect 482938 190294 513478 190350
rect 513534 190294 513602 190350
rect 513658 190294 544198 190350
rect 544254 190294 544322 190350
rect 544378 190294 574918 190350
rect 574974 190294 575042 190350
rect 575098 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 295578 190226
rect 295634 190170 295702 190226
rect 295758 190170 304902 190226
rect 304958 190170 305026 190226
rect 305082 190170 314226 190226
rect 314282 190170 314350 190226
rect 314406 190170 323550 190226
rect 323606 190170 323674 190226
rect 323730 190170 359878 190226
rect 359934 190170 360002 190226
rect 360058 190170 390598 190226
rect 390654 190170 390722 190226
rect 390778 190170 421318 190226
rect 421374 190170 421442 190226
rect 421498 190170 452038 190226
rect 452094 190170 452162 190226
rect 452218 190170 482758 190226
rect 482814 190170 482882 190226
rect 482938 190170 513478 190226
rect 513534 190170 513602 190226
rect 513658 190170 544198 190226
rect 544254 190170 544322 190226
rect 544378 190170 574918 190226
rect 574974 190170 575042 190226
rect 575098 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 295578 190102
rect 295634 190046 295702 190102
rect 295758 190046 304902 190102
rect 304958 190046 305026 190102
rect 305082 190046 314226 190102
rect 314282 190046 314350 190102
rect 314406 190046 323550 190102
rect 323606 190046 323674 190102
rect 323730 190046 359878 190102
rect 359934 190046 360002 190102
rect 360058 190046 390598 190102
rect 390654 190046 390722 190102
rect 390778 190046 421318 190102
rect 421374 190046 421442 190102
rect 421498 190046 452038 190102
rect 452094 190046 452162 190102
rect 452218 190046 482758 190102
rect 482814 190046 482882 190102
rect 482938 190046 513478 190102
rect 513534 190046 513602 190102
rect 513658 190046 544198 190102
rect 544254 190046 544322 190102
rect 544378 190046 574918 190102
rect 574974 190046 575042 190102
rect 575098 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 295578 189978
rect 295634 189922 295702 189978
rect 295758 189922 304902 189978
rect 304958 189922 305026 189978
rect 305082 189922 314226 189978
rect 314282 189922 314350 189978
rect 314406 189922 323550 189978
rect 323606 189922 323674 189978
rect 323730 189922 359878 189978
rect 359934 189922 360002 189978
rect 360058 189922 390598 189978
rect 390654 189922 390722 189978
rect 390778 189922 421318 189978
rect 421374 189922 421442 189978
rect 421498 189922 452038 189978
rect 452094 189922 452162 189978
rect 452218 189922 482758 189978
rect 482814 189922 482882 189978
rect 482938 189922 513478 189978
rect 513534 189922 513602 189978
rect 513658 189922 544198 189978
rect 544254 189922 544322 189978
rect 544378 189922 574918 189978
rect 574974 189922 575042 189978
rect 575098 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 290916 184350
rect 290972 184294 291040 184350
rect 291096 184294 300240 184350
rect 300296 184294 300364 184350
rect 300420 184294 309564 184350
rect 309620 184294 309688 184350
rect 309744 184294 318888 184350
rect 318944 184294 319012 184350
rect 319068 184294 344518 184350
rect 344574 184294 344642 184350
rect 344698 184294 375238 184350
rect 375294 184294 375362 184350
rect 375418 184294 405958 184350
rect 406014 184294 406082 184350
rect 406138 184294 436678 184350
rect 436734 184294 436802 184350
rect 436858 184294 467398 184350
rect 467454 184294 467522 184350
rect 467578 184294 498118 184350
rect 498174 184294 498242 184350
rect 498298 184294 528838 184350
rect 528894 184294 528962 184350
rect 529018 184294 559558 184350
rect 559614 184294 559682 184350
rect 559738 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 290916 184226
rect 290972 184170 291040 184226
rect 291096 184170 300240 184226
rect 300296 184170 300364 184226
rect 300420 184170 309564 184226
rect 309620 184170 309688 184226
rect 309744 184170 318888 184226
rect 318944 184170 319012 184226
rect 319068 184170 344518 184226
rect 344574 184170 344642 184226
rect 344698 184170 375238 184226
rect 375294 184170 375362 184226
rect 375418 184170 405958 184226
rect 406014 184170 406082 184226
rect 406138 184170 436678 184226
rect 436734 184170 436802 184226
rect 436858 184170 467398 184226
rect 467454 184170 467522 184226
rect 467578 184170 498118 184226
rect 498174 184170 498242 184226
rect 498298 184170 528838 184226
rect 528894 184170 528962 184226
rect 529018 184170 559558 184226
rect 559614 184170 559682 184226
rect 559738 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 290916 184102
rect 290972 184046 291040 184102
rect 291096 184046 300240 184102
rect 300296 184046 300364 184102
rect 300420 184046 309564 184102
rect 309620 184046 309688 184102
rect 309744 184046 318888 184102
rect 318944 184046 319012 184102
rect 319068 184046 344518 184102
rect 344574 184046 344642 184102
rect 344698 184046 375238 184102
rect 375294 184046 375362 184102
rect 375418 184046 405958 184102
rect 406014 184046 406082 184102
rect 406138 184046 436678 184102
rect 436734 184046 436802 184102
rect 436858 184046 467398 184102
rect 467454 184046 467522 184102
rect 467578 184046 498118 184102
rect 498174 184046 498242 184102
rect 498298 184046 528838 184102
rect 528894 184046 528962 184102
rect 529018 184046 559558 184102
rect 559614 184046 559682 184102
rect 559738 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 290916 183978
rect 290972 183922 291040 183978
rect 291096 183922 300240 183978
rect 300296 183922 300364 183978
rect 300420 183922 309564 183978
rect 309620 183922 309688 183978
rect 309744 183922 318888 183978
rect 318944 183922 319012 183978
rect 319068 183922 344518 183978
rect 344574 183922 344642 183978
rect 344698 183922 375238 183978
rect 375294 183922 375362 183978
rect 375418 183922 405958 183978
rect 406014 183922 406082 183978
rect 406138 183922 436678 183978
rect 436734 183922 436802 183978
rect 436858 183922 467398 183978
rect 467454 183922 467522 183978
rect 467578 183922 498118 183978
rect 498174 183922 498242 183978
rect 498298 183922 528838 183978
rect 528894 183922 528962 183978
rect 529018 183922 559558 183978
rect 559614 183922 559682 183978
rect 559738 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect 336012 173098 341476 173114
rect 336012 173042 336028 173098
rect 336084 173042 341404 173098
rect 341460 173042 341476 173098
rect 336012 173026 341476 173042
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 295578 172350
rect 295634 172294 295702 172350
rect 295758 172294 304902 172350
rect 304958 172294 305026 172350
rect 305082 172294 314226 172350
rect 314282 172294 314350 172350
rect 314406 172294 323550 172350
rect 323606 172294 323674 172350
rect 323730 172294 359878 172350
rect 359934 172294 360002 172350
rect 360058 172294 390598 172350
rect 390654 172294 390722 172350
rect 390778 172294 421318 172350
rect 421374 172294 421442 172350
rect 421498 172294 452038 172350
rect 452094 172294 452162 172350
rect 452218 172294 482758 172350
rect 482814 172294 482882 172350
rect 482938 172294 513478 172350
rect 513534 172294 513602 172350
rect 513658 172294 544198 172350
rect 544254 172294 544322 172350
rect 544378 172294 574918 172350
rect 574974 172294 575042 172350
rect 575098 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 295578 172226
rect 295634 172170 295702 172226
rect 295758 172170 304902 172226
rect 304958 172170 305026 172226
rect 305082 172170 314226 172226
rect 314282 172170 314350 172226
rect 314406 172170 323550 172226
rect 323606 172170 323674 172226
rect 323730 172170 359878 172226
rect 359934 172170 360002 172226
rect 360058 172170 390598 172226
rect 390654 172170 390722 172226
rect 390778 172170 421318 172226
rect 421374 172170 421442 172226
rect 421498 172170 452038 172226
rect 452094 172170 452162 172226
rect 452218 172170 482758 172226
rect 482814 172170 482882 172226
rect 482938 172170 513478 172226
rect 513534 172170 513602 172226
rect 513658 172170 544198 172226
rect 544254 172170 544322 172226
rect 544378 172170 574918 172226
rect 574974 172170 575042 172226
rect 575098 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 295578 172102
rect 295634 172046 295702 172102
rect 295758 172046 304902 172102
rect 304958 172046 305026 172102
rect 305082 172046 314226 172102
rect 314282 172046 314350 172102
rect 314406 172046 323550 172102
rect 323606 172046 323674 172102
rect 323730 172046 359878 172102
rect 359934 172046 360002 172102
rect 360058 172046 390598 172102
rect 390654 172046 390722 172102
rect 390778 172046 421318 172102
rect 421374 172046 421442 172102
rect 421498 172046 452038 172102
rect 452094 172046 452162 172102
rect 452218 172046 482758 172102
rect 482814 172046 482882 172102
rect 482938 172046 513478 172102
rect 513534 172046 513602 172102
rect 513658 172046 544198 172102
rect 544254 172046 544322 172102
rect 544378 172046 574918 172102
rect 574974 172046 575042 172102
rect 575098 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 295578 171978
rect 295634 171922 295702 171978
rect 295758 171922 304902 171978
rect 304958 171922 305026 171978
rect 305082 171922 314226 171978
rect 314282 171922 314350 171978
rect 314406 171922 323550 171978
rect 323606 171922 323674 171978
rect 323730 171922 359878 171978
rect 359934 171922 360002 171978
rect 360058 171922 390598 171978
rect 390654 171922 390722 171978
rect 390778 171922 421318 171978
rect 421374 171922 421442 171978
rect 421498 171922 452038 171978
rect 452094 171922 452162 171978
rect 452218 171922 482758 171978
rect 482814 171922 482882 171978
rect 482938 171922 513478 171978
rect 513534 171922 513602 171978
rect 513658 171922 544198 171978
rect 544254 171922 544322 171978
rect 544378 171922 574918 171978
rect 574974 171922 575042 171978
rect 575098 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect 295244 170578 297572 170594
rect 295244 170522 295260 170578
rect 295316 170522 297500 170578
rect 297556 170522 297572 170578
rect 295244 170506 297572 170522
rect 293340 169858 297460 169874
rect 293340 169802 293356 169858
rect 293412 169802 297388 169858
rect 297444 169802 297460 169858
rect 293340 169786 297460 169802
rect 336012 168058 341364 168074
rect 336012 168002 336028 168058
rect 336084 168002 341292 168058
rect 341348 168002 341364 168058
rect 336012 167986 341364 168002
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 290916 166350
rect 290972 166294 291040 166350
rect 291096 166294 300240 166350
rect 300296 166294 300364 166350
rect 300420 166294 309564 166350
rect 309620 166294 309688 166350
rect 309744 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 318888 166350
rect 318944 166294 319012 166350
rect 319068 166294 344518 166350
rect 344574 166294 344642 166350
rect 344698 166294 375238 166350
rect 375294 166294 375362 166350
rect 375418 166294 405958 166350
rect 406014 166294 406082 166350
rect 406138 166294 436678 166350
rect 436734 166294 436802 166350
rect 436858 166294 467398 166350
rect 467454 166294 467522 166350
rect 467578 166294 498118 166350
rect 498174 166294 498242 166350
rect 498298 166294 528838 166350
rect 528894 166294 528962 166350
rect 529018 166294 559558 166350
rect 559614 166294 559682 166350
rect 559738 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 290916 166226
rect 290972 166170 291040 166226
rect 291096 166170 300240 166226
rect 300296 166170 300364 166226
rect 300420 166170 309564 166226
rect 309620 166170 309688 166226
rect 309744 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 318888 166226
rect 318944 166170 319012 166226
rect 319068 166170 344518 166226
rect 344574 166170 344642 166226
rect 344698 166170 375238 166226
rect 375294 166170 375362 166226
rect 375418 166170 405958 166226
rect 406014 166170 406082 166226
rect 406138 166170 436678 166226
rect 436734 166170 436802 166226
rect 436858 166170 467398 166226
rect 467454 166170 467522 166226
rect 467578 166170 498118 166226
rect 498174 166170 498242 166226
rect 498298 166170 528838 166226
rect 528894 166170 528962 166226
rect 529018 166170 559558 166226
rect 559614 166170 559682 166226
rect 559738 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 290916 166102
rect 290972 166046 291040 166102
rect 291096 166046 300240 166102
rect 300296 166046 300364 166102
rect 300420 166046 309564 166102
rect 309620 166046 309688 166102
rect 309744 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 318888 166102
rect 318944 166046 319012 166102
rect 319068 166046 344518 166102
rect 344574 166046 344642 166102
rect 344698 166046 375238 166102
rect 375294 166046 375362 166102
rect 375418 166046 405958 166102
rect 406014 166046 406082 166102
rect 406138 166046 436678 166102
rect 436734 166046 436802 166102
rect 436858 166046 467398 166102
rect 467454 166046 467522 166102
rect 467578 166046 498118 166102
rect 498174 166046 498242 166102
rect 498298 166046 528838 166102
rect 528894 166046 528962 166102
rect 529018 166046 559558 166102
rect 559614 166046 559682 166102
rect 559738 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 290916 165978
rect 290972 165922 291040 165978
rect 291096 165922 300240 165978
rect 300296 165922 300364 165978
rect 300420 165922 309564 165978
rect 309620 165922 309688 165978
rect 309744 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 318888 165978
rect 318944 165922 319012 165978
rect 319068 165922 344518 165978
rect 344574 165922 344642 165978
rect 344698 165922 375238 165978
rect 375294 165922 375362 165978
rect 375418 165922 405958 165978
rect 406014 165922 406082 165978
rect 406138 165922 436678 165978
rect 436734 165922 436802 165978
rect 436858 165922 467398 165978
rect 467454 165922 467522 165978
rect 467578 165922 498118 165978
rect 498174 165922 498242 165978
rect 498298 165922 528838 165978
rect 528894 165922 528962 165978
rect 529018 165922 559558 165978
rect 559614 165922 559682 165978
rect 559738 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect 336124 162298 341252 162314
rect 336124 162242 336140 162298
rect 336196 162242 341180 162298
rect 341236 162242 341252 162298
rect 336124 162226 341252 162242
rect 326604 162118 341588 162134
rect 326604 162062 326620 162118
rect 326676 162062 341516 162118
rect 341572 162062 341588 162118
rect 326604 162046 341588 162062
rect 274972 161218 591348 161234
rect 274972 161162 274988 161218
rect 275044 161162 591276 161218
rect 591332 161162 591348 161218
rect 274972 161146 591348 161162
rect 276540 161038 590564 161054
rect 276540 160982 276556 161038
rect 276612 160982 590492 161038
rect 590548 160982 590564 161038
rect 276540 160966 590564 160982
rect 340044 160858 590900 160874
rect 340044 160802 340060 160858
rect 340116 160802 590828 160858
rect 590884 160802 590900 160858
rect 340044 160786 590900 160802
rect 281692 159598 357940 159614
rect 281692 159542 281708 159598
rect 281764 159542 357868 159598
rect 357924 159542 357940 159598
rect 281692 159526 357940 159542
rect 328956 158698 576340 158714
rect 328956 158642 328972 158698
rect 329028 158642 576268 158698
rect 576324 158642 576340 158698
rect 328956 158626 576340 158642
rect 325148 157798 591124 157814
rect 325148 157742 325164 157798
rect 325220 157742 591052 157798
rect 591108 157742 591124 157798
rect 325148 157726 591124 157742
rect 340492 157618 558532 157634
rect 340492 157562 340508 157618
rect 340564 157562 558460 157618
rect 558516 157562 558532 157618
rect 340492 157546 558532 157562
rect 340828 157438 514180 157454
rect 340828 157382 340844 157438
rect 340900 157382 514108 157438
rect 514164 157382 514180 157438
rect 340828 157366 514180 157382
rect 333772 155638 574884 155654
rect 333772 155582 333788 155638
rect 333844 155582 574812 155638
rect 574868 155582 574884 155638
rect 333772 155566 574884 155582
rect 327164 155458 578132 155474
rect 327164 155402 327180 155458
rect 327236 155402 578060 155458
rect 578116 155402 578132 155458
rect 327164 155386 578132 155402
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect 294908 152758 590116 152774
rect 294908 152702 294924 152758
rect 294980 152702 590044 152758
rect 590100 152702 590116 152758
rect 294908 152686 590116 152702
rect 285276 152038 590676 152054
rect 285276 151982 285292 152038
rect 285348 151982 590604 152038
rect 590660 151982 590676 152038
rect 285276 151966 590676 151982
rect 283148 150418 590564 150434
rect 283148 150362 283164 150418
rect 283220 150362 590492 150418
rect 590548 150362 590564 150418
rect 283148 150346 590564 150362
rect 457980 149698 576452 149714
rect 457980 149642 457996 149698
rect 458052 149642 576380 149698
rect 576436 149642 576452 149698
rect 457980 149626 576452 149642
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect 332316 146998 574996 147014
rect 332316 146942 332332 146998
rect 332388 146942 574924 146998
rect 574980 146942 574996 146998
rect 332316 146926 574996 146942
rect 338700 145378 574660 145394
rect 338700 145322 338716 145378
rect 338772 145322 574588 145378
rect 574644 145322 574660 145378
rect 338700 145306 574660 145322
rect 466716 144838 490100 144854
rect 466716 144782 466732 144838
rect 466788 144782 490028 144838
rect 490084 144782 490100 144838
rect 466716 144766 490100 144782
rect 463132 144658 497940 144674
rect 463132 144602 463148 144658
rect 463204 144602 497868 144658
rect 497924 144602 497940 144658
rect 463132 144586 497940 144602
rect 290596 144478 505780 144494
rect 290596 144422 290668 144478
rect 290724 144422 505708 144478
rect 505764 144422 505780 144478
rect 290596 144406 505780 144422
rect 290596 143954 290684 144406
rect 272956 143938 290684 143954
rect 272956 143882 272972 143938
rect 273028 143882 290684 143938
rect 272956 143866 290684 143882
rect 336124 143938 513620 143954
rect 336124 143882 336140 143938
rect 336196 143882 337148 143938
rect 337204 143882 513548 143938
rect 513604 143882 513620 143938
rect 336124 143866 513620 143882
rect 280124 143758 507348 143774
rect 280124 143702 280140 143758
rect 280196 143702 507276 143758
rect 507332 143702 507348 143758
rect 280124 143686 507348 143702
rect 273180 143578 508916 143594
rect 273180 143522 273196 143578
rect 273252 143522 273756 143578
rect 273812 143522 508844 143578
rect 508900 143522 508916 143578
rect 273180 143506 508916 143522
rect 267916 143398 272260 143414
rect 267916 143342 267932 143398
rect 267988 143342 272188 143398
rect 272244 143342 272260 143398
rect 267916 143326 272260 143342
rect 272172 142858 512052 142874
rect 272172 142802 272188 142858
rect 272244 142802 511980 142858
rect 512036 142802 512052 142858
rect 272172 142786 512052 142802
rect 331980 142678 472964 142694
rect 331980 142622 331996 142678
rect 332052 142622 472892 142678
rect 472948 142622 472964 142678
rect 331980 142606 472964 142622
rect 338588 142498 468708 142514
rect 338588 142442 338604 142498
rect 338660 142442 468636 142498
rect 468692 142442 468708 142498
rect 338588 142426 468708 142442
rect 332428 141958 578020 141974
rect 332428 141902 332444 141958
rect 332500 141902 577948 141958
rect 578004 141902 578020 141958
rect 332428 141886 578020 141902
rect 463244 141238 590788 141254
rect 463244 141182 463260 141238
rect 463316 141182 590716 141238
rect 590772 141182 590788 141238
rect 463244 141166 590788 141182
rect 326828 140338 578916 140354
rect 326828 140282 326844 140338
rect 326900 140282 578844 140338
rect 578900 140282 578916 140338
rect 326828 140266 578916 140282
rect 465372 139798 480692 139814
rect 465372 139742 465388 139798
rect 465444 139742 480620 139798
rect 480676 139742 480692 139798
rect 465372 139726 480692 139742
rect 465484 139618 482260 139634
rect 465484 139562 465500 139618
rect 465556 139562 482188 139618
rect 482244 139562 482260 139618
rect 465484 139546 482260 139562
rect 278220 139438 590228 139454
rect 278220 139382 278236 139438
rect 278292 139382 590156 139438
rect 590212 139382 590228 139438
rect 278220 139366 590228 139382
rect 340940 138538 574324 138554
rect 340940 138482 340956 138538
rect 341012 138482 574252 138538
rect 574308 138482 574324 138538
rect 340940 138466 574324 138482
rect 335004 137638 466804 137654
rect 335004 137582 335020 137638
rect 335076 137582 466732 137638
rect 466788 137582 466804 137638
rect 335004 137566 466804 137582
rect 337636 137458 462996 137474
rect 337636 137402 462924 137458
rect 462980 137402 462996 137458
rect 337636 137386 462996 137402
rect 337636 136934 337724 137386
rect 306556 136918 337724 136934
rect 306556 136862 306572 136918
rect 306628 136862 336812 136918
rect 336868 136862 337724 136918
rect 306556 136846 337724 136862
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 572038 136350
rect 572094 136294 572162 136350
rect 572218 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 572038 136226
rect 572094 136170 572162 136226
rect 572218 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 572038 136102
rect 572094 136046 572162 136102
rect 572218 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 572038 135978
rect 572094 135922 572162 135978
rect 572218 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect 297372 135658 463220 135674
rect 297372 135602 297388 135658
rect 297444 135602 463148 135658
rect 463204 135602 463220 135658
rect 297372 135586 463220 135602
rect 367036 135478 466468 135494
rect 367036 135422 367052 135478
rect 367108 135422 466396 135478
rect 466452 135422 466468 135478
rect 367036 135406 466468 135422
rect 333324 135298 465460 135314
rect 333324 135242 333340 135298
rect 333396 135242 465388 135298
rect 465444 135242 465460 135298
rect 333324 135226 465460 135242
rect 293116 134578 297460 134594
rect 293116 134522 293132 134578
rect 293188 134522 297388 134578
rect 297444 134522 297460 134578
rect 293116 134506 297460 134522
rect 285164 134398 463332 134414
rect 285164 134342 285180 134398
rect 285236 134342 463260 134398
rect 463316 134342 463332 134398
rect 285164 134326 463332 134342
rect 336012 134218 467140 134234
rect 336012 134162 336028 134218
rect 336084 134162 336812 134218
rect 336868 134162 467068 134218
rect 467124 134162 467140 134218
rect 336012 134146 467140 134162
rect 335900 134038 466692 134054
rect 335900 133982 335916 134038
rect 335972 133982 466620 134038
rect 466676 133982 466692 134038
rect 335900 133966 466692 133982
rect 304876 132778 336100 132794
rect 304876 132722 304892 132778
rect 304948 132722 336028 132778
rect 336084 132722 336100 132778
rect 304876 132706 336100 132722
rect 274972 132598 463108 132614
rect 274972 132542 274988 132598
rect 275044 132542 282604 132598
rect 282660 132542 463036 132598
rect 463092 132542 463108 132598
rect 274972 132526 463108 132542
rect 290596 132418 462884 132434
rect 290596 132362 292348 132418
rect 292404 132362 462812 132418
rect 462868 132362 462884 132418
rect 290596 132346 462884 132362
rect 290596 131894 290684 132346
rect 336796 132238 465572 132254
rect 336796 132182 336812 132238
rect 336868 132182 337708 132238
rect 337764 132182 465500 132238
rect 465556 132182 465572 132238
rect 336796 132166 465572 132182
rect 280236 131878 290684 131894
rect 280236 131822 280252 131878
rect 280308 131822 290684 131878
rect 280236 131806 290684 131822
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 556678 130350
rect 556734 130294 556802 130350
rect 556858 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 556678 130226
rect 556734 130170 556802 130226
rect 556858 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 556678 130102
rect 556734 130046 556802 130102
rect 556858 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 556678 129978
rect 556734 129922 556802 129978
rect 556858 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect 333884 127558 466356 127574
rect 333884 127502 333900 127558
rect 333956 127502 337148 127558
rect 337204 127502 466284 127558
rect 466340 127502 466356 127558
rect 333884 127486 466356 127502
rect 423260 122518 466244 122534
rect 423260 122462 423276 122518
rect 423332 122462 466172 122518
rect 466228 122462 466244 122518
rect 423260 122446 466244 122462
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 572038 118350
rect 572094 118294 572162 118350
rect 572218 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 572038 118226
rect 572094 118170 572162 118226
rect 572218 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 572038 118102
rect 572094 118046 572162 118102
rect 572218 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 572038 117978
rect 572094 117922 572162 117978
rect 572218 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect 268700 115318 413380 115334
rect 268700 115262 268716 115318
rect 268772 115262 413308 115318
rect 413364 115262 413380 115318
rect 268700 115246 413380 115262
rect 268588 115138 415060 115154
rect 268588 115082 268604 115138
rect 268660 115082 414988 115138
rect 415044 115082 415060 115138
rect 268588 115066 415060 115082
rect 574124 113878 575220 113894
rect 574124 113822 574140 113878
rect 574196 113822 575148 113878
rect 575204 113822 575220 113878
rect 574124 113806 575220 113822
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 556678 112350
rect 556734 112294 556802 112350
rect 556858 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 556678 112226
rect 556734 112170 556802 112226
rect 556858 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 556678 112102
rect 556734 112046 556802 112102
rect 556858 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 556678 111978
rect 556734 111922 556802 111978
rect 556858 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect 281356 104158 406772 104174
rect 281356 104102 281372 104158
rect 281428 104102 406700 104158
rect 406756 104102 406772 104158
rect 281356 104086 406772 104102
rect 283036 103978 403300 103994
rect 283036 103922 283052 103978
rect 283108 103922 403228 103978
rect 403284 103922 403300 103978
rect 283036 103906 403300 103922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 572038 100350
rect 572094 100294 572162 100350
rect 572218 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 572038 100226
rect 572094 100170 572162 100226
rect 572218 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 572038 100102
rect 572094 100046 572162 100102
rect 572218 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 572038 99978
rect 572094 99922 572162 99978
rect 572218 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 374518 94350
rect 374574 94294 374642 94350
rect 374698 94294 405238 94350
rect 405294 94294 405362 94350
rect 405418 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 556678 94350
rect 556734 94294 556802 94350
rect 556858 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 374518 94226
rect 374574 94170 374642 94226
rect 374698 94170 405238 94226
rect 405294 94170 405362 94226
rect 405418 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 556678 94226
rect 556734 94170 556802 94226
rect 556858 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 374518 94102
rect 374574 94046 374642 94102
rect 374698 94046 405238 94102
rect 405294 94046 405362 94102
rect 405418 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 556678 94102
rect 556734 94046 556802 94102
rect 556858 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 374518 93978
rect 374574 93922 374642 93978
rect 374698 93922 405238 93978
rect 405294 93922 405362 93978
rect 405418 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 556678 93978
rect 556734 93922 556802 93978
rect 556858 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 389878 82350
rect 389934 82294 390002 82350
rect 390058 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 572038 82350
rect 572094 82294 572162 82350
rect 572218 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 389878 82226
rect 389934 82170 390002 82226
rect 390058 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 572038 82226
rect 572094 82170 572162 82226
rect 572218 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82147 597980 82170
rect -1916 82102 299528 82147
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82091 299528 82102
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82102 597980 82147
rect 324740 82091 347154 82102
rect 286142 82046 347154 82091
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 389878 82102
rect 389934 82046 390002 82102
rect 390058 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 572038 82102
rect 572094 82046 572162 82102
rect 572218 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 82043 597980 82046
rect -1916 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 597980 82043
rect -1916 81978 597980 81987
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81939 347154 81978
rect 286142 81922 299528 81939
rect -1916 81883 299528 81922
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81922 347154 81939
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 389878 81978
rect 389934 81922 390002 81978
rect 390058 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 572038 81978
rect 572094 81922 572162 81978
rect 572218 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 324740 81883 597980 81922
rect -1916 81826 597980 81883
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 374518 76350
rect 374574 76294 374642 76350
rect 374698 76294 405238 76350
rect 405294 76294 405362 76350
rect 405418 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 556678 76350
rect 556734 76294 556802 76350
rect 556858 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 374518 76226
rect 374574 76170 374642 76226
rect 374698 76170 405238 76226
rect 405294 76170 405362 76226
rect 405418 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 556678 76226
rect 556734 76170 556802 76226
rect 556858 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 374518 76102
rect 374574 76046 374642 76102
rect 374698 76046 405238 76102
rect 405294 76046 405362 76102
rect 405418 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 556678 76102
rect 556734 76046 556802 76102
rect 556858 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 374518 75978
rect 374574 75922 374642 75978
rect 374698 75922 405238 75978
rect 405294 75922 405362 75978
rect 405418 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 556678 75978
rect 556734 75922 556802 75978
rect 556858 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 389878 64350
rect 389934 64294 390002 64350
rect 390058 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 572038 64350
rect 572094 64294 572162 64350
rect 572218 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 389878 64226
rect 389934 64170 390002 64226
rect 390058 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 572038 64226
rect 572094 64170 572162 64226
rect 572218 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 389878 64102
rect 389934 64046 390002 64102
rect 390058 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 572038 64102
rect 572094 64046 572162 64102
rect 572218 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 389878 63978
rect 389934 63922 390002 63978
rect 390058 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 572038 63978
rect 572094 63922 572162 63978
rect 572218 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 374518 58350
rect 374574 58294 374642 58350
rect 374698 58294 405238 58350
rect 405294 58294 405362 58350
rect 405418 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 556678 58350
rect 556734 58294 556802 58350
rect 556858 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 374518 58226
rect 374574 58170 374642 58226
rect 374698 58170 405238 58226
rect 405294 58170 405362 58226
rect 405418 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 556678 58226
rect 556734 58170 556802 58226
rect 556858 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 374518 58102
rect 374574 58046 374642 58102
rect 374698 58046 405238 58102
rect 405294 58046 405362 58102
rect 405418 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 556678 58102
rect 556734 58046 556802 58102
rect 556858 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 374518 57978
rect 374574 57922 374642 57978
rect 374698 57922 405238 57978
rect 405294 57922 405362 57978
rect 405418 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 556678 57978
rect 556734 57922 556802 57978
rect 556858 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 4268 55378 270692 55394
rect 4268 55322 4284 55378
rect 4340 55322 270620 55378
rect 270676 55322 270692 55378
rect 4268 55306 270692 55322
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 479878 46350
rect 479934 46294 480002 46350
rect 480058 46294 510598 46350
rect 510654 46294 510722 46350
rect 510778 46294 541318 46350
rect 541374 46294 541442 46350
rect 541498 46294 572038 46350
rect 572094 46294 572162 46350
rect 572218 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 479878 46226
rect 479934 46170 480002 46226
rect 480058 46170 510598 46226
rect 510654 46170 510722 46226
rect 510778 46170 541318 46226
rect 541374 46170 541442 46226
rect 541498 46170 572038 46226
rect 572094 46170 572162 46226
rect 572218 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 479878 46102
rect 479934 46046 480002 46102
rect 480058 46046 510598 46102
rect 510654 46046 510722 46102
rect 510778 46046 541318 46102
rect 541374 46046 541442 46102
rect 541498 46046 572038 46102
rect 572094 46046 572162 46102
rect 572218 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 479878 45978
rect 479934 45922 480002 45978
rect 480058 45922 510598 45978
rect 510654 45922 510722 45978
rect 510778 45922 541318 45978
rect 541374 45922 541442 45978
rect 541498 45922 572038 45978
rect 572094 45922 572162 45978
rect 572218 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 464518 40350
rect 464574 40294 464642 40350
rect 464698 40294 495238 40350
rect 495294 40294 495362 40350
rect 495418 40294 525958 40350
rect 526014 40294 526082 40350
rect 526138 40294 556678 40350
rect 556734 40294 556802 40350
rect 556858 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 464518 40226
rect 464574 40170 464642 40226
rect 464698 40170 495238 40226
rect 495294 40170 495362 40226
rect 495418 40170 525958 40226
rect 526014 40170 526082 40226
rect 526138 40170 556678 40226
rect 556734 40170 556802 40226
rect 556858 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 464518 40102
rect 464574 40046 464642 40102
rect 464698 40046 495238 40102
rect 495294 40046 495362 40102
rect 495418 40046 525958 40102
rect 526014 40046 526082 40102
rect 526138 40046 556678 40102
rect 556734 40046 556802 40102
rect 556858 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 464518 39978
rect 464574 39922 464642 39978
rect 464698 39922 495238 39978
rect 495294 39922 495362 39978
rect 495418 39922 525958 39978
rect 526014 39922 526082 39978
rect 526138 39922 556678 39978
rect 556734 39922 556802 39978
rect 556858 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect 276316 35218 590004 35234
rect 276316 35162 276332 35218
rect 276388 35162 589932 35218
rect 589988 35162 590004 35218
rect 276316 35146 590004 35162
rect 334220 33598 578244 33614
rect 334220 33542 334236 33598
rect 334292 33542 578172 33598
rect 578228 33542 578244 33598
rect 334220 33526 578244 33542
rect 330748 31798 578020 31814
rect 330748 31742 330764 31798
rect 330820 31742 577948 31798
rect 578004 31742 578020 31798
rect 330748 31726 578020 31742
rect 339260 30178 574660 30194
rect 339260 30122 339276 30178
rect 339332 30122 574588 30178
rect 574644 30122 574660 30178
rect 339260 30106 574660 30122
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 479878 28350
rect 479934 28294 480002 28350
rect 480058 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 510598 28350
rect 510654 28294 510722 28350
rect 510778 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 541318 28350
rect 541374 28294 541442 28350
rect 541498 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 572038 28350
rect 572094 28294 572162 28350
rect 572218 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 479878 28226
rect 479934 28170 480002 28226
rect 480058 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 510598 28226
rect 510654 28170 510722 28226
rect 510778 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 541318 28226
rect 541374 28170 541442 28226
rect 541498 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 572038 28226
rect 572094 28170 572162 28226
rect 572218 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 479878 28102
rect 479934 28046 480002 28102
rect 480058 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 510598 28102
rect 510654 28046 510722 28102
rect 510778 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 541318 28102
rect 541374 28046 541442 28102
rect 541498 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 572038 28102
rect 572094 28046 572162 28102
rect 572218 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 479878 27978
rect 479934 27922 480002 27978
rect 480058 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 510598 27978
rect 510654 27922 510722 27978
rect 510778 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 541318 27978
rect 541374 27922 541442 27978
rect 541498 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 572038 27978
rect 572094 27922 572162 27978
rect 572218 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use avali_logo  avali_logo
timestamp 0
transform 1 0 60000 0 1 475000
box 0 0 90000 105660
use wrapped_ay8913  ay8913
timestamp 0
transform 1 0 40000 0 1 240000
box 1120 0 51000 51000
use blinker  blinker
timestamp 0
transform 1 0 290000 0 1 50000
box 1258 0 34768 32230
use diceroll  diceroll
timestamp 0
transform 1 0 45000 0 1 315000
box 1258 3050 44662 46000
use hellorld  hellorld
timestamp 0
transform 1 0 135000 0 1 260000
box 1258 1792 26000 26000
use wrapped_mc14500  mc14500
timestamp 0
transform 1 0 285000 0 1 160000
box 1120 0 40000 40000
use multiplexer  multiplexer
timestamp 0
transform 1 0 180000 0 1 240000
box 0 0 150000 140000
use wrapped_sid  sid
timestamp 0
transform 1 0 40000 0 1 50000
box 1258 0 230000 160000
use tholin_avalonsemi_tbb1143  tbb1143
timestamp 0
transform 1 0 115000 0 1 320000
box 1258 2688 46000 43120
use ue1  ue1
timestamp 0
transform 1 0 60000 0 1 390000
box 1258 1568 24000 24000
use wrapped_pdp11  wrapped_pdp11
timestamp 0
transform 1 0 190000 0 1 410000
box 0 0 340000 156886
use wrapped_qcpu  wrapped_qcpu
timestamp 0
transform 1 0 460000 0 1 20000
box 0 3050 115000 120000
use wrapped_sn76489  wrapped_sn76489
timestamp 0
transform 1 0 370000 0 1 50000
box 0 2688 50000 50000
use wrapped_tholin_riscv  wrapped_tholin_riscv
timestamp 0
transform 1 0 340000 0 1 160000
box 0 0 243686 245000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal output
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal output
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal output
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal output
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal output
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal output
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal output
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal output
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal output
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal output
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal output
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal output
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal output
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal output
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal output
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal output
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal output
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal output
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal output
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal output
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal output
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal output
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal output
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal output
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal output
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal output
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal output
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal output
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal output
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal output
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal output
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal output
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal output
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal output
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal output
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal output
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal output
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal output
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal output
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal output
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal output
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal output
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal output
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal output
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal output
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal output
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal output
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal output
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal output
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal output
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal output
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal output
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal output
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal output
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal output
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal output
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal output
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal output
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal output
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal output
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal output
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal output
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal output
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal output
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal output
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal output
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal output
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal output
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal output
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal output
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal output
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal output
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal output
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal output
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal output
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal output
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal output
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal output
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal output
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal output
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal output
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal output
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal output
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal output
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal output
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal output
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal output
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal output
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal output
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal output
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal output
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal output
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal output
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal output
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal output
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal output
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal output
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal output
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal output
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal output
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal output
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal output
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal output
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal output
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal output
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal output
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal output
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal output
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal output
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal output
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal output
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal output
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal output
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal output
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal output
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal output
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal output
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal output
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal output
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal output
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal output
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal output
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal output
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal output
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal output
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal output
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal output
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal output
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal output
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal output
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal output
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal output
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal output
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal output
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal output
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal output
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal output
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal output
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal output
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal output
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal output
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal output
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal output
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 53002 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 205590 67478 241770 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 289526 67478 337490 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 351422 67478 390964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 412556 67478 486928 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 535792 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 53002 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 205590 98198 472944 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 549832 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 53002 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 205590 128918 488604 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 53002 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 205590 159638 260964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 284908 159638 322218 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 359670 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 53002 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 205590 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 53002 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 205590 221078 239082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 379126 221078 409194 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 568502 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 53002 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 205590 251798 239082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 379126 251798 409194 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 568502 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 239082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 379126 282518 409194 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 568502 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 53674 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 77350 313238 170618 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 197430 313238 239082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 379126 313238 409194 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 568502 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 159418 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 568502 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 50964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 98428 374678 159418 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 568502 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 50964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 98428 405398 159418 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 568502 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 159418 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 568502 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 34090 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 568502 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 34090 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 402950 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 34090 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 402950 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 34090 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 402950 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 53002 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 205590 71198 241770 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 289526 71198 337490 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 351422 71198 400170 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 405142 71198 482968 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 539752 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 53002 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 205590 101918 473124 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 549472 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 53002 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 205590 132638 322218 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 359670 132638 490764 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 578452 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 53002 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 205590 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 53002 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 205590 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 53002 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 205590 224798 239082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 379126 224798 409194 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 568502 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 53002 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 205590 255518 239082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 379126 255518 409194 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 568502 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 239082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 379126 286238 409194 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 568502 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 50964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 84316 316958 170618 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 197430 316958 239082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 379126 316958 409194 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 568502 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 159418 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 568502 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 51210 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 97622 378398 159418 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 568502 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 -1644 409118 51210 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 97622 409118 159418 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 568502 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 159418 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 568502 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 34090 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 568502 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 34090 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 402950 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 34090 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 402950 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 34090 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 402950 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal output
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal output
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal output
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal output
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal output
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal output
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal output
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal output
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal output
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal output
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal output
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal output
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal output
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal output
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal output
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal output
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal output
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal output
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal output
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal output
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal output
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal output
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal output
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal output
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal output
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal output
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal output
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal output
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal output
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal output
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal output
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal output
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal output
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 559710 400322 559710 400322 0 vdd
rlabel via4 575070 388322 575070 388322 0 vss
rlabel metal2 40810 240744 40810 240744 0 ay8913_do\[0\]
rlabel metal2 59080 238994 59080 238994 0 ay8913_do\[10\]
rlabel metal3 129136 240520 129136 240520 0 ay8913_do\[11\]
rlabel metal2 62664 236698 62664 236698 0 ay8913_do\[12\]
rlabel metal2 77336 238896 77336 238896 0 ay8913_do\[13\]
rlabel metal3 122584 240072 122584 240072 0 ay8913_do\[14\]
rlabel via4 68040 237705 68040 237705 0 ay8913_do\[15\]
rlabel metal2 69832 238938 69832 238938 0 ay8913_do\[16\]
rlabel metal4 71624 237559 71624 237559 0 ay8913_do\[17\]
rlabel metal2 73416 238994 73416 238994 0 ay8913_do\[18\]
rlabel metal2 75208 239106 75208 239106 0 ay8913_do\[19\]
rlabel metal2 42952 239274 42952 239274 0 ay8913_do\[1\]
rlabel metal2 77000 238826 77000 238826 0 ay8913_do\[20\]
rlabel metal2 78792 239050 78792 239050 0 ay8913_do\[21\]
rlabel metal2 95144 313544 95144 313544 0 ay8913_do\[22\]
rlabel metal2 234696 382550 234696 382550 0 ay8913_do\[23\]
rlabel metal2 94920 313432 94920 313432 0 ay8913_do\[24\]
rlabel metal2 236040 381038 236040 381038 0 ay8913_do\[25\]
rlabel metal2 99960 314328 99960 314328 0 ay8913_do\[26\]
rlabel metal2 237384 385798 237384 385798 0 ay8913_do\[27\]
rlabel metal3 79072 240408 79072 240408 0 ay8913_do\[2\]
rlabel metal2 46536 239218 46536 239218 0 ay8913_do\[3\]
rlabel metal2 118440 311248 118440 311248 0 ay8913_do\[4\]
rlabel metal3 105280 240184 105280 240184 0 ay8913_do\[5\]
rlabel metal2 51912 239162 51912 239162 0 ay8913_do\[6\]
rlabel metal2 116760 311024 116760 311024 0 ay8913_do\[7\]
rlabel metal2 55496 239106 55496 239106 0 ay8913_do\[8\]
rlabel metal2 57288 239946 57288 239946 0 ay8913_do\[9\]
rlabel metal2 307944 49266 307944 49266 0 blinker_do\[0\]
rlabel metal4 285096 131432 285096 131432 0 blinker_do\[1\]
rlabel metal4 288680 132328 288680 132328 0 blinker_do\[2\]
rlabel metal3 189602 428904 189602 428904 0 custom_settings\[0\]
rlabel metal4 191576 236544 191576 236544 0 custom_settings\[10\]
rlabel metal3 333494 288008 333494 288008 0 custom_settings\[11\]
rlabel metal3 331310 288904 331310 288904 0 custom_settings\[12\]
rlabel metal3 188258 522088 188258 522088 0 custom_settings\[13\]
rlabel metal3 332976 308056 332976 308056 0 custom_settings\[14\]
rlabel metal3 331478 291592 331478 291592 0 custom_settings\[15\]
rlabel metal4 330344 249312 330344 249312 0 custom_settings\[16\]
rlabel metal4 332472 248640 332472 248640 0 custom_settings\[17\]
rlabel metal3 188874 557928 188874 557928 0 custom_settings\[18\]
rlabel metal3 188986 565096 188986 565096 0 custom_settings\[19\]
rlabel metal3 92302 280392 92302 280392 0 custom_settings\[1\]
rlabel metal4 330120 257628 330120 257628 0 custom_settings\[20\]
rlabel metal3 459368 101836 459368 101836 0 custom_settings\[21\]
rlabel metal3 331464 264264 331464 264264 0 custom_settings\[22\]
rlabel metal4 327432 237510 327432 237510 0 custom_settings\[23\]
rlabel metal3 330960 264040 330960 264040 0 custom_settings\[24\]
rlabel metal3 330862 300552 330862 300552 0 custom_settings\[25\]
rlabel metal3 330918 301448 330918 301448 0 custom_settings\[26\]
rlabel metal3 331590 302344 331590 302344 0 custom_settings\[27\]
rlabel metal3 332150 303240 332150 303240 0 custom_settings\[28\]
rlabel metal3 332710 304136 332710 304136 0 custom_settings\[29\]
rlabel metal4 161896 282576 161896 282576 0 custom_settings\[2\]
rlabel metal3 332640 282184 332640 282184 0 custom_settings\[30\]
rlabel metal3 332486 305928 332486 305928 0 custom_settings\[31\]
rlabel metal3 163016 282184 163016 282184 0 custom_settings\[3\]
rlabel metal3 332206 281736 332206 281736 0 custom_settings\[4\]
rlabel metal4 187320 283410 187320 283410 0 custom_settings\[5\]
rlabel metal3 189042 471912 189042 471912 0 custom_settings\[6\]
rlabel metal4 188104 285210 188104 285210 0 custom_settings\[7\]
rlabel metal4 195944 284400 195944 284400 0 custom_settings\[8\]
rlabel metal3 188706 493416 188706 493416 0 custom_settings\[9\]
rlabel metal2 58296 370342 58296 370342 0 diceroll_do\[0\]
rlabel metal2 306600 381710 306600 381710 0 diceroll_do\[1\]
rlabel metal2 307272 381654 307272 381654 0 diceroll_do\[2\]
rlabel metal2 69720 374598 69720 374598 0 diceroll_do\[3\]
rlabel metal2 73528 373702 73528 373702 0 diceroll_do\[4\]
rlabel metal2 77336 362446 77336 362446 0 diceroll_do\[5\]
rlabel metal2 81144 370398 81144 370398 0 diceroll_do\[6\]
rlabel metal3 197792 379400 197792 379400 0 diceroll_do\[7\]
rlabel metal2 311304 383446 311304 383446 0 diceroll_do\[8\]
rlabel metal2 165704 326144 165704 326144 0 hellorld_do
rlabel metal2 190582 379512 190582 379512 0 io_in[0]
rlabel metal3 92190 263368 92190 263368 0 io_in[10]
rlabel metal3 327096 117544 327096 117544 0 io_in[11]
rlabel metal2 287336 238280 287336 238280 0 io_in[12]
rlabel metal4 232344 406999 232344 406999 0 io_in[13]
rlabel metal3 332584 261408 332584 261408 0 io_in[14]
rlabel metal2 331912 260960 331912 260960 0 io_in[15]
rlabel metal3 337232 262920 337232 262920 0 io_in[16]
rlabel metal3 332416 237272 332416 237272 0 io_in[17]
rlabel metal2 259448 409682 259448 409682 0 io_in[18]
rlabel metal2 282184 93744 282184 93744 0 io_in[19]
rlabel metal3 332864 289016 332864 289016 0 io_in[20]
rlabel metal3 188384 590184 188384 590184 0 io_in[21]
rlabel metal2 493192 143094 493192 143094 0 io_in[22]
rlabel metal4 336056 145208 336056 145208 0 io_in[23]
rlabel metal3 2702 587160 2702 587160 0 io_in[24]
rlabel metal3 2310 544824 2310 544824 0 io_in[25]
rlabel metal4 4368 420000 4368 420000 0 io_in[26]
rlabel metal3 306320 406616 306320 406616 0 io_in[27]
rlabel metal2 468552 141512 468552 141512 0 io_in[28]
rlabel metal3 2310 375704 2310 375704 0 io_in[29]
rlabel metal3 2310 333368 2310 333368 0 io_in[30]
rlabel metal5 331912 360810 331912 360810 0 io_in[31]
rlabel metal4 4648 247761 4648 247761 0 io_in[32]
rlabel metal3 2254 206360 2254 206360 0 io_in[33]
rlabel metal3 336448 383544 336448 383544 0 io_in[34]
rlabel metal4 336168 141983 336168 141983 0 io_in[35]
rlabel metal3 329784 236432 329784 236432 0 io_in[36]
rlabel metal4 336168 401856 336168 401856 0 io_in[37]
rlabel metal3 92904 241976 92904 241976 0 io_in[5]
rlabel metal2 467978 139944 467978 139944 0 io_in[6]
rlabel metal3 171808 374584 171808 374584 0 io_in[7]
rlabel metal4 374584 403760 374584 403760 0 io_in[8]
rlabel metal2 163688 405608 163688 405608 0 io_in[9]
rlabel metal4 589960 34479 589960 34479 0 io_oeb[0]
rlabel metal3 593474 430136 593474 430136 0 io_oeb[10]
rlabel metal3 593082 469896 593082 469896 0 io_oeb[11]
rlabel metal3 593194 509544 593194 509544 0 io_oeb[12]
rlabel metal3 593250 549192 593250 549192 0 io_oeb[13]
rlabel metal3 593082 588616 593082 588616 0 io_oeb[14]
rlabel metal2 172872 422464 172872 422464 0 io_oeb[15]
rlabel metal2 172984 423864 172984 423864 0 io_oeb[16]
rlabel metal2 408296 592242 408296 592242 0 io_oeb[17]
rlabel metal5 260400 571950 260400 571950 0 io_oeb[18]
rlabel metal3 227696 570472 227696 570472 0 io_oeb[19]
rlabel metal3 593138 73416 593138 73416 0 io_oeb[1]
rlabel metal2 209608 589722 209608 589722 0 io_oeb[20]
rlabel metal2 143416 589778 143416 589778 0 io_oeb[21]
rlabel metal2 77448 592242 77448 592242 0 io_oeb[22]
rlabel metal2 168840 286664 168840 286664 0 io_oeb[23]
rlabel metal3 2422 558936 2422 558936 0 io_oeb[24]
rlabel metal3 2478 516600 2478 516600 0 io_oeb[25]
rlabel metal3 2534 474264 2534 474264 0 io_oeb[26]
rlabel metal4 162120 356608 162120 356608 0 io_oeb[27]
rlabel metal3 2366 389592 2366 389592 0 io_oeb[28]
rlabel metal3 2366 347256 2366 347256 0 io_oeb[29]
rlabel metal4 281624 183176 281624 183176 0 io_oeb[2]
rlabel metal3 77910 304920 77910 304920 0 io_oeb[30]
rlabel metal3 2366 262808 2366 262808 0 io_oeb[31]
rlabel metal3 144186 286888 144186 286888 0 io_oeb[32]
rlabel metal3 2366 178024 2366 178024 0 io_oeb[33]
rlabel metal4 29400 212352 29400 212352 0 io_oeb[34]
rlabel metal3 5670 93464 5670 93464 0 io_oeb[35]
rlabel metal4 27720 171136 27720 171136 0 io_oeb[36]
rlabel metal3 2310 8792 2310 8792 0 io_oeb[37]
rlabel via4 590072 152721 590072 152721 0 io_oeb[3]
rlabel metal3 593026 192136 593026 192136 0 io_oeb[4]
rlabel metal3 593418 231896 593418 231896 0 io_oeb[5]
rlabel metal4 195832 237737 195832 237737 0 io_oeb[6]
rlabel metal3 593194 311080 593194 311080 0 io_oeb[7]
rlabel metal3 593138 350728 593138 350728 0 io_oeb[8]
rlabel metal4 187432 248845 187432 248845 0 io_oeb[9]
rlabel metal2 191198 379512 191198 379512 0 io_out[0]
rlabel metal3 593082 417032 593082 417032 0 io_out[10]
rlabel metal3 593194 456680 593194 456680 0 io_out[11]
rlabel metal3 593138 496328 593138 496328 0 io_out[12]
rlabel metal4 189560 475384 189560 475384 0 io_out[13]
rlabel metal4 189224 489795 189224 489795 0 io_out[14]
rlabel metal2 562632 593082 562632 593082 0 io_out[15]
rlabel metal2 496440 593194 496440 593194 0 io_out[16]
rlabel metal2 430248 593306 430248 593306 0 io_out[17]
rlabel metal2 189672 498400 189672 498400 0 io_out[18]
rlabel metal2 189560 500920 189560 500920 0 io_out[19]
rlabel metal2 191926 379512 191926 379512 0 io_out[1]
rlabel metal2 189784 497112 189784 497112 0 io_out[20]
rlabel metal2 165704 593082 165704 593082 0 io_out[21]
rlabel metal2 99512 593138 99512 593138 0 io_out[22]
rlabel metal2 33320 593082 33320 593082 0 io_out[23]
rlabel metal2 52920 481824 52920 481824 0 io_out[24]
rlabel metal5 132328 404010 132328 404010 0 io_out[25]
rlabel metal5 110488 402390 110488 402390 0 io_out[26]
rlabel metal2 94920 421736 94920 421736 0 io_out[27]
rlabel metal3 30030 403704 30030 403704 0 io_out[28]
rlabel metal3 56966 361368 56966 361368 0 io_out[29]
rlabel metal2 192542 379512 192542 379512 0 io_out[2]
rlabel metal2 44520 349328 44520 349328 0 io_out[30]
rlabel metal3 17430 276696 17430 276696 0 io_out[31]
rlabel metal2 24360 309232 24360 309232 0 io_out[32]
rlabel metal4 213192 379229 213192 379229 0 io_out[33]
rlabel metal4 213864 379049 213864 379049 0 io_out[34]
rlabel metal3 7350 107352 7350 107352 0 io_out[35]
rlabel metal4 215208 379139 215208 379139 0 io_out[36]
rlabel metal3 2310 22904 2310 22904 0 io_out[37]
rlabel via4 590184 139397 590184 139397 0 io_out[3]
rlabel metal2 193522 379512 193522 379512 0 io_out[4]
rlabel metal2 194558 379512 194558 379512 0 io_out[5]
rlabel metal3 195608 379288 195608 379288 0 io_out[6]
rlabel metal5 192304 288990 192304 288990 0 io_out[7]
rlabel metal5 376264 403110 376264 403110 0 io_out[8]
rlabel metal3 591402 377384 591402 377384 0 io_out[9]
rlabel metal2 288232 214102 288232 214102 0 mc14500_do\[0\]
rlabel metal3 177338 332808 177338 332808 0 mc14500_do\[10\]
rlabel metal2 172648 279384 172648 279384 0 mc14500_do\[11\]
rlabel metal2 172312 284032 172312 284032 0 mc14500_do\[12\]
rlabel metal2 302792 214774 302792 214774 0 mc14500_do\[13\]
rlabel metal2 171080 280224 171080 280224 0 mc14500_do\[14\]
rlabel metal2 305032 215670 305032 215670 0 mc14500_do\[15\]
rlabel metal2 170968 283808 170968 283808 0 mc14500_do\[16\]
rlabel metal2 172424 287672 172424 287672 0 mc14500_do\[17\]
rlabel metal2 169512 278880 169512 278880 0 mc14500_do\[18\]
rlabel metal2 169400 280336 169400 280336 0 mc14500_do\[19\]
rlabel metal2 289352 209846 289352 209846 0 mc14500_do\[1\]
rlabel metal2 171192 284312 171192 284312 0 mc14500_do\[20\]
rlabel metal2 167720 284088 167720 284088 0 mc14500_do\[21\]
rlabel metal2 169624 281064 169624 281064 0 mc14500_do\[22\]
rlabel metal2 167944 284144 167944 284144 0 mc14500_do\[23\]
rlabel metal2 172760 290696 172760 290696 0 mc14500_do\[24\]
rlabel metal3 179746 349608 179746 349608 0 mc14500_do\[25\]
rlabel metal3 178178 350728 178178 350728 0 mc14500_do\[26\]
rlabel metal3 180152 351554 180152 351554 0 mc14500_do\[27\]
rlabel metal2 171304 292096 171304 292096 0 mc14500_do\[28\]
rlabel metal2 167832 291032 167832 291032 0 mc14500_do\[29\]
rlabel metal2 169288 279328 169288 279328 0 mc14500_do\[2\]
rlabel metal2 166264 289856 166264 289856 0 mc14500_do\[30\]
rlabel metal2 166040 277368 166040 277368 0 mc14500_do\[3\]
rlabel metal3 177226 326088 177226 326088 0 mc14500_do\[4\]
rlabel metal2 167608 280168 167608 280168 0 mc14500_do\[5\]
rlabel metal2 166152 279832 166152 279832 0 mc14500_do\[6\]
rlabel metal2 172536 276360 172536 276360 0 mc14500_do\[7\]
rlabel metal2 170856 278376 170856 278376 0 mc14500_do\[8\]
rlabel metal3 179690 331688 179690 331688 0 mc14500_do\[9\]
rlabel metal3 285600 160552 285600 160552 0 mc14500_sram_addr\[0\]
rlabel metal2 313096 237090 313096 237090 0 mc14500_sram_addr\[1\]
rlabel metal2 313992 237146 313992 237146 0 mc14500_sram_addr\[2\]
rlabel metal2 284648 178808 284648 178808 0 mc14500_sram_addr\[3\]
rlabel metal2 283640 178696 283640 178696 0 mc14500_sram_addr\[4\]
rlabel metal2 283752 178416 283752 178416 0 mc14500_sram_addr\[5\]
rlabel metal2 324240 236936 324240 236936 0 mc14500_sram_gwe
rlabel metal2 283416 178472 283416 178472 0 mc14500_sram_in\[0\]
rlabel metal5 296408 170550 296408 170550 0 mc14500_sram_in\[1\]
rlabel metal2 300552 158634 300552 158634 0 mc14500_sram_in\[2\]
rlabel metal2 302344 158914 302344 158914 0 mc14500_sram_in\[3\]
rlabel metal2 321160 238826 321160 238826 0 mc14500_sram_in\[4\]
rlabel metal2 305928 158858 305928 158858 0 mc14500_sram_in\[5\]
rlabel metal2 322952 238770 322952 238770 0 mc14500_sram_in\[6\]
rlabel metal2 309512 158970 309512 158970 0 mc14500_sram_in\[7\]
rlabel metal2 238056 395038 238056 395038 0 pdp11_do\[0\]
rlabel metal4 193144 482328 193144 482328 0 pdp11_do\[10\]
rlabel metal3 295260 406728 295260 406728 0 pdp11_do\[11\]
rlabel metal3 189392 566104 189392 566104 0 pdp11_do\[12\]
rlabel metal2 255528 392350 255528 392350 0 pdp11_do\[13\]
rlabel metal4 383208 403592 383208 403592 0 pdp11_do\[14\]
rlabel metal2 258216 386358 258216 386358 0 pdp11_do\[15\]
rlabel metal2 259560 392294 259560 392294 0 pdp11_do\[16\]
rlabel metal2 260904 380814 260904 380814 0 pdp11_do\[17\]
rlabel metal2 262248 380982 262248 380982 0 pdp11_do\[18\]
rlabel metal2 263592 381262 263592 381262 0 pdp11_do\[19\]
rlabel metal2 239400 381150 239400 381150 0 pdp11_do\[1\]
rlabel metal2 264936 394534 264936 394534 0 pdp11_do\[20\]
rlabel metal2 266280 381990 266280 381990 0 pdp11_do\[21\]
rlabel metal4 403256 404656 403256 404656 0 pdp11_do\[22\]
rlabel metal4 192584 488544 192584 488544 0 pdp11_do\[23\]
rlabel metal2 270312 381206 270312 381206 0 pdp11_do\[24\]
rlabel metal2 491288 407890 491288 407890 0 pdp11_do\[25\]
rlabel metal4 356664 405771 356664 405771 0 pdp11_do\[26\]
rlabel metal4 356216 404320 356216 404320 0 pdp11_do\[27\]
rlabel metal2 275688 387982 275688 387982 0 pdp11_do\[28\]
rlabel metal2 277032 381262 277032 381262 0 pdp11_do\[29\]
rlabel metal2 240744 391174 240744 391174 0 pdp11_do\[2\]
rlabel metal4 517048 404503 517048 404503 0 pdp11_do\[30\]
rlabel metal4 522200 405403 522200 405403 0 pdp11_do\[31\]
rlabel metal2 281064 388038 281064 388038 0 pdp11_do\[32\]
rlabel metal2 242088 392238 242088 392238 0 pdp11_do\[3\]
rlabel metal2 243432 381934 243432 381934 0 pdp11_do\[4\]
rlabel metal2 358344 408912 358344 408912 0 pdp11_do\[5\]
rlabel metal3 192640 567112 192640 567112 0 pdp11_do\[6\]
rlabel metal2 378840 409976 378840 409976 0 pdp11_do\[7\]
rlabel metal5 355656 401490 355656 401490 0 pdp11_do\[8\]
rlabel metal2 250152 387926 250152 387926 0 pdp11_do\[9\]
rlabel metal2 238728 394590 238728 394590 0 pdp11_oeb\[0\]
rlabel metal4 192808 486472 192808 486472 0 pdp11_oeb\[10\]
rlabel metal3 225568 407512 225568 407512 0 pdp11_oeb\[11\]
rlabel metal3 227136 407736 227136 407736 0 pdp11_oeb\[12\]
rlabel metal4 196168 486472 196168 486472 0 pdp11_oeb\[13\]
rlabel metal2 189224 485296 189224 485296 0 pdp11_oeb\[14\]
rlabel metal2 189448 487200 189448 487200 0 pdp11_oeb\[15\]
rlabel metal2 189336 489608 189336 489608 0 pdp11_oeb\[16\]
rlabel metal4 195944 488152 195944 488152 0 pdp11_oeb\[17\]
rlabel metal4 196280 488600 196280 488600 0 pdp11_oeb\[18\]
rlabel metal2 264264 392406 264264 392406 0 pdp11_oeb\[19\]
rlabel metal2 188104 483784 188104 483784 0 pdp11_oeb\[1\]
rlabel metal4 192920 487032 192920 487032 0 pdp11_oeb\[20\]
rlabel metal2 266952 387982 266952 387982 0 pdp11_oeb\[21\]
rlabel metal2 268296 381206 268296 381206 0 pdp11_oeb\[22\]
rlabel metal3 233688 404376 233688 404376 0 pdp11_oeb\[23\]
rlabel metal3 234416 399336 234416 399336 0 pdp11_oeb\[24\]
rlabel metal3 201936 398104 201936 398104 0 pdp11_oeb\[25\]
rlabel metal3 236600 404152 236600 404152 0 pdp11_oeb\[26\]
rlabel metal3 238784 404264 238784 404264 0 pdp11_oeb\[27\]
rlabel metal3 238840 397656 238840 397656 0 pdp11_oeb\[28\]
rlabel metal3 240184 400680 240184 400680 0 pdp11_oeb\[29\]
rlabel metal3 190008 567112 190008 567112 0 pdp11_oeb\[2\]
rlabel metal2 279048 388766 279048 388766 0 pdp11_oeb\[30\]
rlabel metal4 189448 487816 189448 487816 0 pdp11_oeb\[31\]
rlabel metal4 189336 488712 189336 488712 0 pdp11_oeb\[32\]
rlabel metal2 242760 380982 242760 380982 0 pdp11_oeb\[3\]
rlabel metal4 191352 485576 191352 485576 0 pdp11_oeb\[4\]
rlabel metal4 193032 484680 193032 484680 0 pdp11_oeb\[5\]
rlabel metal3 190904 567336 190904 567336 0 pdp11_oeb\[6\]
rlabel metal3 216440 402808 216440 402808 0 pdp11_oeb\[7\]
rlabel metal4 196392 485408 196392 485408 0 pdp11_oeb\[8\]
rlabel metal2 187992 487984 187992 487984 0 pdp11_oeb\[9\]
rlabel metal2 518280 141078 518280 141078 0 qcpu_do\[0\]
rlabel metal2 514920 149800 514920 149800 0 qcpu_do\[10\]
rlabel metal2 279048 191394 279048 191394 0 qcpu_do\[11\]
rlabel metal2 279944 200186 279944 200186 0 qcpu_do\[12\]
rlabel metal2 538664 142870 538664 142870 0 qcpu_do\[13\]
rlabel metal2 540232 142814 540232 142814 0 qcpu_do\[14\]
rlabel metal2 541800 142758 541800 142758 0 qcpu_do\[15\]
rlabel metal2 543368 142702 543368 142702 0 qcpu_do\[16\]
rlabel metal3 519960 143696 519960 143696 0 qcpu_do\[17\]
rlabel metal3 518560 143976 518560 143976 0 qcpu_do\[18\]
rlabel metal2 285544 237608 285544 237608 0 qcpu_do\[19\]
rlabel metal2 519848 142534 519848 142534 0 qcpu_do\[1\]
rlabel metal3 284648 237048 284648 237048 0 qcpu_do\[20\]
rlabel metal3 284256 237160 284256 237160 0 qcpu_do\[21\]
rlabel metal3 286384 236936 286384 236936 0 qcpu_do\[22\]
rlabel metal3 290528 236936 290528 236936 0 qcpu_do\[23\]
rlabel metal2 285544 192304 285544 192304 0 qcpu_do\[24\]
rlabel metal2 280392 192472 280392 192472 0 qcpu_do\[25\]
rlabel metal4 288904 192528 288904 192528 0 qcpu_do\[26\]
rlabel metal2 293832 238504 293832 238504 0 qcpu_do\[27\]
rlabel metal2 562184 146118 562184 146118 0 qcpu_do\[28\]
rlabel metal2 563752 141750 563752 141750 0 qcpu_do\[29\]
rlabel metal2 521416 142254 521416 142254 0 qcpu_do\[2\]
rlabel metal2 565320 145502 565320 145502 0 qcpu_do\[30\]
rlabel metal2 566888 142646 566888 142646 0 qcpu_do\[31\]
rlabel metal2 568456 144326 568456 144326 0 qcpu_do\[32\]
rlabel metal2 522984 142030 522984 142030 0 qcpu_do\[3\]
rlabel metal2 524552 144438 524552 144438 0 qcpu_do\[4\]
rlabel metal2 526120 143766 526120 143766 0 qcpu_do\[5\]
rlabel metal3 275296 237048 275296 237048 0 qcpu_do\[6\]
rlabel metal2 275464 238490 275464 238490 0 qcpu_do\[7\]
rlabel metal3 277088 236936 277088 236936 0 qcpu_do\[8\]
rlabel metal3 278376 237048 278376 237048 0 qcpu_do\[9\]
rlabel metal3 331982 306824 331982 306824 0 qcpu_oeb\[0\]
rlabel metal1 332472 261352 332472 261352 0 qcpu_oeb\[10\]
rlabel metal3 327768 188104 327768 188104 0 qcpu_oeb\[11\]
rlabel metal3 330624 285656 330624 285656 0 qcpu_oeb\[12\]
rlabel metal3 332808 189784 332808 189784 0 qcpu_oeb\[13\]
rlabel metal3 335328 297192 335328 297192 0 qcpu_oeb\[14\]
rlabel metal4 472920 142921 472920 142921 0 qcpu_oeb\[15\]
rlabel metal5 329560 249570 329560 249570 0 qcpu_oeb\[16\]
rlabel metal3 331142 322056 331142 322056 0 qcpu_oeb\[17\]
rlabel metal3 332766 322952 332766 322952 0 qcpu_oeb\[18\]
rlabel metal3 330736 240296 330736 240296 0 qcpu_oeb\[19\]
rlabel metal2 335944 106344 335944 106344 0 qcpu_oeb\[1\]
rlabel metal5 456680 145350 456680 145350 0 qcpu_oeb\[20\]
rlabel metal3 334222 325640 334222 325640 0 qcpu_oeb\[21\]
rlabel metal5 330848 283770 330848 283770 0 qcpu_oeb\[22\]
rlabel metal4 468664 142775 468664 142775 0 qcpu_oeb\[23\]
rlabel metal3 332206 328328 332206 328328 0 qcpu_oeb\[24\]
rlabel metal5 329504 253710 329504 253710 0 qcpu_oeb\[25\]
rlabel metal4 327320 237690 327320 237690 0 qcpu_oeb\[26\]
rlabel metal5 329056 240390 329056 240390 0 qcpu_oeb\[27\]
rlabel metal4 333816 190841 333816 190841 0 qcpu_oeb\[28\]
rlabel metal3 332262 332808 332262 332808 0 qcpu_oeb\[29\]
rlabel metal3 331814 308616 331814 308616 0 qcpu_oeb\[2\]
rlabel metal4 329336 240390 329336 240390 0 qcpu_oeb\[30\]
rlabel metal3 333480 287448 333480 287448 0 qcpu_oeb\[31\]
rlabel metal3 335286 335496 335286 335496 0 qcpu_oeb\[32\]
rlabel metal3 334670 309512 334670 309512 0 qcpu_oeb\[3\]
rlabel metal3 335118 310408 335118 310408 0 qcpu_oeb\[4\]
rlabel metal4 335384 284480 335384 284480 0 qcpu_oeb\[5\]
rlabel metal3 335062 312200 335062 312200 0 qcpu_oeb\[6\]
rlabel metal3 328888 240296 328888 240296 0 qcpu_oeb\[7\]
rlabel metal4 329168 314010 329168 314010 0 qcpu_oeb\[8\]
rlabel metal4 327600 237330 327600 237330 0 qcpu_oeb\[9\]
rlabel metal3 576926 91112 576926 91112 0 qcpu_sram_addr\[0\]
rlabel metal3 575246 93128 575246 93128 0 qcpu_sram_addr\[1\]
rlabel metal3 575974 95144 575974 95144 0 qcpu_sram_addr\[2\]
rlabel metal4 290472 169680 290472 169680 0 qcpu_sram_addr\[3\]
rlabel metal1 301504 235816 301504 235816 0 qcpu_sram_addr\[4\]
rlabel metal3 303352 199416 303352 199416 0 qcpu_sram_addr\[5\]
rlabel metal3 314664 238168 314664 238168 0 qcpu_sram_gwe
rlabel metal4 305704 217392 305704 217392 0 qcpu_sram_in\[0\]
rlabel metal3 315112 238280 315112 238280 0 qcpu_sram_in\[1\]
rlabel metal3 574728 107366 574728 107366 0 qcpu_sram_in\[2\]
rlabel metal3 316568 238392 316568 238392 0 qcpu_sram_in\[3\]
rlabel metal4 308616 199136 308616 199136 0 qcpu_sram_in\[4\]
rlabel metal2 309512 221410 309512 221410 0 qcpu_sram_in\[5\]
rlabel metal3 310632 199416 310632 199416 0 qcpu_sram_in\[6\]
rlabel metal2 311598 240072 311598 240072 0 qcpu_sram_in\[7\]
rlabel metal3 335216 266280 335216 266280 0 qcpu_sram_out\[0\]
rlabel metal3 336224 265496 336224 265496 0 qcpu_sram_out\[1\]
rlabel metal3 335720 191576 335720 191576 0 qcpu_sram_out\[2\]
rlabel metal3 333424 156296 333424 156296 0 qcpu_sram_out\[3\]
rlabel metal2 332696 156968 332696 156968 0 qcpu_sram_out\[4\]
rlabel metal3 331478 340872 331478 340872 0 qcpu_sram_out\[5\]
rlabel metal3 331870 341768 331870 341768 0 qcpu_sram_out\[6\]
rlabel metal3 331982 342664 331982 342664 0 qcpu_sram_out\[7\]
rlabel metal3 331310 343560 331310 343560 0 rst_ay8913
rlabel metal3 228032 239512 228032 239512 0 rst_blinker
rlabel metal3 51912 364504 51912 364504 0 rst_diceroll
rlabel metal2 147784 302974 147784 302974 0 rst_hellorld
rlabel metal4 169624 265664 169624 265664 0 rst_mc14500
rlabel metal3 188202 421736 188202 421736 0 rst_pdp11
rlabel metal3 224336 216328 224336 216328 0 rst_qcpu
rlabel metal2 212296 48930 212296 48930 0 rst_sid
rlabel metal3 240688 220024 240688 220024 0 rst_sn76489
rlabel metal4 163800 332304 163800 332304 0 rst_tbb1143
rlabel metal4 196392 296968 196392 296968 0 rst_tholin_riscv
rlabel metal2 311976 383614 311976 383614 0 rst_ue1
rlabel metal3 271222 148792 271222 148792 0 sid_do\[0\]
rlabel metal3 179746 305928 179746 305928 0 sid_do\[10\]
rlabel metal4 180264 259056 180264 259056 0 sid_do\[11\]
rlabel metal4 171304 263200 171304 263200 0 sid_do\[12\]
rlabel metal3 177170 309288 177170 309288 0 sid_do\[13\]
rlabel metal3 177282 310408 177282 310408 0 sid_do\[14\]
rlabel metal4 169512 263872 169512 263872 0 sid_do\[15\]
rlabel metal3 178962 312648 178962 312648 0 sid_do\[16\]
rlabel metal3 178122 313768 178122 313768 0 sid_do\[17\]
rlabel metal3 222824 239736 222824 239736 0 sid_do\[18\]
rlabel metal4 180152 262528 180152 262528 0 sid_do\[19\]
rlabel metal3 178850 295848 178850 295848 0 sid_do\[1\]
rlabel metal3 179802 317128 179802 317128 0 sid_do\[20\]
rlabel metal3 178738 296968 178738 296968 0 sid_do\[2\]
rlabel metal4 270760 220050 270760 220050 0 sid_do\[3\]
rlabel metal3 226464 239624 226464 239624 0 sid_do\[4\]
rlabel metal3 271334 163352 271334 163352 0 sid_do\[5\]
rlabel metal4 172984 255416 172984 255416 0 sid_do\[6\]
rlabel metal4 166264 266224 166264 266224 0 sid_do\[7\]
rlabel metal3 178906 303688 178906 303688 0 sid_do\[8\]
rlabel metal4 167944 268184 167944 268184 0 sid_do\[9\]
rlabel metal2 154952 213374 154952 213374 0 sid_oeb
rlabel metal2 373618 99960 373618 99960 0 sn76489_do\[0\]
rlabel metal2 389018 99960 389018 99960 0 sn76489_do\[10\]
rlabel metal2 390586 99960 390586 99960 0 sn76489_do\[11\]
rlabel metal2 392154 99960 392154 99960 0 sn76489_do\[12\]
rlabel metal2 255752 226674 255752 226674 0 sn76489_do\[13\]
rlabel metal2 256648 227906 256648 227906 0 sn76489_do\[14\]
rlabel metal2 396858 99960 396858 99960 0 sn76489_do\[15\]
rlabel metal2 398706 99960 398706 99960 0 sn76489_do\[16\]
rlabel metal2 400274 99960 400274 99960 0 sn76489_do\[17\]
rlabel metal2 401842 99960 401842 99960 0 sn76489_do\[18\]
rlabel metal2 403354 99960 403354 99960 0 sn76489_do\[19\]
rlabel metal2 375186 99960 375186 99960 0 sn76489_do\[1\]
rlabel metal2 404978 99960 404978 99960 0 sn76489_do\[20\]
rlabel metal2 406686 99960 406686 99960 0 sn76489_do\[21\]
rlabel metal3 264880 237048 264880 237048 0 sn76489_do\[22\]
rlabel metal2 265384 238504 265384 238504 0 sn76489_do\[23\]
rlabel metal3 266560 236936 266560 236936 0 sn76489_do\[24\]
rlabel metal2 267064 238504 267064 238504 0 sn76489_do\[25\]
rlabel metal3 268408 237048 268408 237048 0 sn76489_do\[26\]
rlabel metal2 268632 238504 268632 238504 0 sn76489_do\[27\]
rlabel metal2 376698 99960 376698 99960 0 sn76489_do\[2\]
rlabel metal2 378210 99960 378210 99960 0 sn76489_do\[3\]
rlabel metal2 379890 99960 379890 99960 0 sn76489_do\[4\]
rlabel metal2 381458 99960 381458 99960 0 sn76489_do\[5\]
rlabel metal2 383166 99960 383166 99960 0 sn76489_do\[6\]
rlabel metal2 384594 99960 384594 99960 0 sn76489_do\[7\]
rlabel metal2 281848 183512 281848 183512 0 sn76489_do\[8\]
rlabel metal2 252168 238826 252168 238826 0 sn76489_do\[9\]
rlabel metal4 171416 354648 171416 354648 0 tbb1143_do\[0\]
rlabel metal3 161098 352968 161098 352968 0 tbb1143_do\[1\]
rlabel metal3 167902 356328 167902 356328 0 tbb1143_do\[2\]
rlabel metal3 161098 359688 161098 359688 0 tbb1143_do\[3\]
rlabel metal3 160888 363174 160888 363174 0 tbb1143_do\[4\]
rlabel metal2 344120 158970 344120 158970 0 tholin_riscv_do\[0\]
rlabel metal3 331702 354312 331702 354312 0 tholin_riscv_do\[10\]
rlabel metal2 425432 157234 425432 157234 0 tholin_riscv_do\[11\]
rlabel metal5 330400 242010 330400 242010 0 tholin_riscv_do\[12\]
rlabel metal3 335062 357000 335062 357000 0 tholin_riscv_do\[13\]
rlabel metal2 447608 158914 447608 158914 0 tholin_riscv_do\[14\]
rlabel metal2 420840 150976 420840 150976 0 tholin_riscv_do\[15\]
rlabel metal3 331632 307944 331632 307944 0 tholin_riscv_do\[16\]
rlabel metal3 332192 307384 332192 307384 0 tholin_riscv_do\[17\]
rlabel metal3 330862 361480 330862 361480 0 tholin_riscv_do\[18\]
rlabel metal5 333088 311670 333088 311670 0 tholin_riscv_do\[19\]
rlabel metal3 332024 308168 332024 308168 0 tholin_riscv_do\[1\]
rlabel metal3 329448 363090 329448 363090 0 tholin_riscv_do\[20\]
rlabel metal2 499352 158522 499352 158522 0 tholin_riscv_do\[21\]
rlabel metal3 330904 309176 330904 309176 0 tholin_riscv_do\[22\]
rlabel metal4 514136 157469 514136 157469 0 tholin_riscv_do\[23\]
rlabel metal3 330848 308392 330848 308392 0 tholin_riscv_do\[24\]
rlabel metal3 336168 277256 336168 277256 0 tholin_riscv_do\[25\]
rlabel metal3 335118 368648 335118 368648 0 tholin_riscv_do\[26\]
rlabel metal3 335608 275688 335608 275688 0 tholin_riscv_do\[27\]
rlabel metal3 335776 283864 335776 283864 0 tholin_riscv_do\[28\]
rlabel metal3 335230 371336 335230 371336 0 tholin_riscv_do\[29\]
rlabel metal3 334600 283864 334600 283864 0 tholin_riscv_do\[2\]
rlabel metal5 328720 260370 328720 260370 0 tholin_riscv_do\[30\]
rlabel metal3 330190 373128 330190 373128 0 tholin_riscv_do\[31\]
rlabel metal5 332248 283050 332248 283050 0 tholin_riscv_do\[32\]
rlabel metal3 331086 348040 331086 348040 0 tholin_riscv_do\[3\]
rlabel metal3 328776 237720 328776 237720 0 tholin_riscv_do\[4\]
rlabel metal3 330974 349832 330974 349832 0 tholin_riscv_do\[5\]
rlabel metal3 334278 350728 334278 350728 0 tholin_riscv_do\[6\]
rlabel metal3 332206 351624 332206 351624 0 tholin_riscv_do\[7\]
rlabel metal3 336112 277480 336112 277480 0 tholin_riscv_do\[8\]
rlabel metal3 329896 353234 329896 353234 0 tholin_riscv_do\[9\]
rlabel metal2 283080 388094 283080 388094 0 tholin_riscv_oeb\[0\]
rlabel metal2 289800 394198 289800 394198 0 tholin_riscv_oeb\[10\]
rlabel metal3 379008 406504 379008 406504 0 tholin_riscv_oeb\[11\]
rlabel metal4 342776 403872 342776 403872 0 tholin_riscv_oeb\[12\]
rlabel metal2 379736 409640 379736 409640 0 tholin_riscv_oeb\[13\]
rlabel metal3 354480 403144 354480 403144 0 tholin_riscv_oeb\[14\]
rlabel metal4 455000 403648 455000 403648 0 tholin_riscv_oeb\[15\]
rlabel metal3 316624 404152 316624 404152 0 tholin_riscv_oeb\[16\]
rlabel metal2 469784 406182 469784 406182 0 tholin_riscv_oeb\[17\]
rlabel metal2 383096 406952 383096 406952 0 tholin_riscv_oeb\[18\]
rlabel metal2 337064 397768 337064 397768 0 tholin_riscv_oeb\[19\]
rlabel metal2 283752 391286 283752 391286 0 tholin_riscv_oeb\[1\]
rlabel metal4 398440 404264 398440 404264 0 tholin_riscv_oeb\[20\]
rlabel metal2 499352 405790 499352 405790 0 tholin_riscv_oeb\[21\]
rlabel metal2 338072 403200 338072 403200 0 tholin_riscv_oeb\[22\]
rlabel metal2 514136 405790 514136 405790 0 tholin_riscv_oeb\[23\]
rlabel metal2 521528 406070 521528 406070 0 tholin_riscv_oeb\[24\]
rlabel metal4 339640 403461 339640 403461 0 tholin_riscv_oeb\[25\]
rlabel metal2 300552 380982 300552 380982 0 tholin_riscv_oeb\[26\]
rlabel metal2 543704 405790 543704 405790 0 tholin_riscv_oeb\[27\]
rlabel metal2 302078 379960 302078 379960 0 tholin_riscv_oeb\[28\]
rlabel metal2 302568 394310 302568 394310 0 tholin_riscv_oeb\[29\]
rlabel metal2 358904 406350 358904 406350 0 tholin_riscv_oeb\[2\]
rlabel metal2 303240 381038 303240 381038 0 tholin_riscv_oeb\[30\]
rlabel metal2 303912 380982 303912 380982 0 tholin_riscv_oeb\[31\]
rlabel metal2 304584 380814 304584 380814 0 tholin_riscv_oeb\[32\]
rlabel metal2 285096 392182 285096 392182 0 tholin_riscv_oeb\[3\]
rlabel metal4 373688 403592 373688 403592 0 tholin_riscv_oeb\[4\]
rlabel metal2 286440 394422 286440 394422 0 tholin_riscv_oeb\[5\]
rlabel metal2 287112 384510 287112 384510 0 tholin_riscv_oeb\[6\]
rlabel metal2 287784 388150 287784 388150 0 tholin_riscv_oeb\[7\]
rlabel metal2 288456 384566 288456 384566 0 tholin_riscv_oeb\[8\]
rlabel metal2 289128 389718 289128 389718 0 tholin_riscv_oeb\[9\]
rlabel metal2 313320 380982 313320 380982 0 ue1_do\[0\]
rlabel metal2 313992 387030 313992 387030 0 ue1_do\[1\]
rlabel metal2 66360 415478 66360 415478 0 ue1_do\[2\]
rlabel metal2 68600 415702 68600 415702 0 ue1_do\[3\]
rlabel metal2 70840 415590 70840 415590 0 ue1_do\[4\]
rlabel metal2 73080 415646 73080 415646 0 ue1_do\[5\]
rlabel metal2 75320 415534 75320 415534 0 ue1_do\[6\]
rlabel metal2 77560 415366 77560 415366 0 ue1_do\[7\]
rlabel metal3 83160 416696 83160 416696 0 ue1_do\[8\]
rlabel metal3 83552 413448 83552 413448 0 ue1_do\[9\]
rlabel metal2 312648 382942 312648 382942 0 ue1_oeb
rlabel metal2 580664 3990 580664 3990 0 user_irq[0]
rlabel metal4 217224 379319 217224 379319 0 user_irq[1]
rlabel metal2 584472 3150 584472 3150 0 user_irq[2]
rlabel metal2 46690 360360 46690 360360 0 wb_clk_i
rlabel metal2 185864 233898 185864 233898 0 wb_rst_i
rlabel metal3 329896 277550 329896 277550 0 wbs_ack_o
rlabel metal2 186760 236362 186760 236362 0 wbs_adr_i[0]
rlabel metal2 195720 237258 195720 237258 0 wbs_adr_i[10]
rlabel metal2 93240 25438 93240 25438 0 wbs_adr_i[11]
rlabel metal2 98952 25550 98952 25550 0 wbs_adr_i[12]
rlabel metal3 71456 49672 71456 49672 0 wbs_adr_i[13]
rlabel metal3 73640 49560 73640 49560 0 wbs_adr_i[14]
rlabel metal2 116088 21742 116088 21742 0 wbs_adr_i[15]
rlabel metal2 121800 16590 121800 16590 0 wbs_adr_i[16]
rlabel metal2 201992 236698 201992 236698 0 wbs_adr_i[17]
rlabel metal2 202888 236754 202888 236754 0 wbs_adr_i[18]
rlabel metal2 138936 16758 138936 16758 0 wbs_adr_i[19]
rlabel metal2 30408 111622 30408 111622 0 wbs_adr_i[1]
rlabel metal2 144648 21854 144648 21854 0 wbs_adr_i[20]
rlabel metal3 212408 46312 212408 46312 0 wbs_adr_i[21]
rlabel metal2 279160 136920 279160 136920 0 wbs_adr_i[22]
rlabel metal2 161784 23422 161784 23422 0 wbs_adr_i[23]
rlabel metal2 167496 25158 167496 25158 0 wbs_adr_i[24]
rlabel metal2 209160 235914 209160 235914 0 wbs_adr_i[25]
rlabel metal2 210056 233954 210056 233954 0 wbs_adr_i[26]
rlabel metal2 210952 234234 210952 234234 0 wbs_adr_i[27]
rlabel metal3 190400 50344 190400 50344 0 wbs_adr_i[28]
rlabel metal4 196056 50960 196056 50960 0 wbs_adr_i[29]
rlabel metal2 188552 234738 188552 234738 0 wbs_adr_i[2]
rlabel metal2 213640 237314 213640 237314 0 wbs_adr_i[30]
rlabel metal2 214536 235466 214536 235466 0 wbs_adr_i[31]
rlabel metal4 45640 50568 45640 50568 0 wbs_adr_i[3]
rlabel metal2 53256 25438 53256 25438 0 wbs_adr_i[4]
rlabel metal2 191240 236418 191240 236418 0 wbs_adr_i[5]
rlabel metal2 192136 226338 192136 226338 0 wbs_adr_i[6]
rlabel metal2 70392 2366 70392 2366 0 wbs_adr_i[7]
rlabel metal2 76104 25270 76104 25270 0 wbs_adr_i[8]
rlabel metal2 194824 235578 194824 235578 0 wbs_adr_i[9]
rlabel metal3 329896 275338 329896 275338 0 wbs_cyc_i
rlabel metal2 24696 106470 24696 106470 0 wbs_dat_i[0]
rlabel metal4 89432 50904 89432 50904 0 wbs_dat_i[10]
rlabel metal2 95144 21630 95144 21630 0 wbs_dat_i[11]
rlabel metal2 100856 23310 100856 23310 0 wbs_dat_i[12]
rlabel metal2 106568 21686 106568 21686 0 wbs_dat_i[13]
rlabel metal2 112280 21798 112280 21798 0 wbs_dat_i[14]
rlabel metal2 117992 19950 117992 19950 0 wbs_dat_i[15]
rlabel metal2 123704 20006 123704 20006 0 wbs_dat_i[16]
rlabel metal2 230664 237146 230664 237146 0 wbs_dat_i[17]
rlabel metal2 231784 238504 231784 238504 0 wbs_dat_i[18]
rlabel metal2 140840 18326 140840 18326 0 wbs_dat_i[19]
rlabel metal2 216328 231378 216328 231378 0 wbs_dat_i[1]
rlabel metal3 233408 236936 233408 236936 0 wbs_dat_i[20]
rlabel metal4 234248 237009 234248 237009 0 wbs_dat_i[21]
rlabel via4 235144 237155 235144 237155 0 wbs_dat_i[22]
rlabel metal2 236040 239050 236040 239050 0 wbs_dat_i[23]
rlabel metal2 169624 2310 169624 2310 0 wbs_dat_i[24]
rlabel metal2 237832 239106 237832 239106 0 wbs_dat_i[25]
rlabel metal2 238728 238882 238728 238882 0 wbs_dat_i[26]
rlabel metal2 239624 239218 239624 239218 0 wbs_dat_i[27]
rlabel metal2 240520 238938 240520 238938 0 wbs_dat_i[28]
rlabel metal4 241416 209496 241416 209496 0 wbs_dat_i[29]
rlabel metal2 217224 229754 217224 229754 0 wbs_dat_i[2]
rlabel metal2 242312 238994 242312 238994 0 wbs_dat_i[30]
rlabel metal4 209384 51072 209384 51072 0 wbs_dat_i[31]
rlabel metal2 218120 227178 218120 227178 0 wbs_dat_i[3]
rlabel metal2 55160 2646 55160 2646 0 wbs_dat_i[4]
rlabel metal2 219912 228858 219912 228858 0 wbs_dat_i[5]
rlabel metal2 66584 2422 66584 2422 0 wbs_dat_i[6]
rlabel metal2 72296 2310 72296 2310 0 wbs_dat_i[7]
rlabel metal2 78008 25214 78008 25214 0 wbs_dat_i[8]
rlabel metal3 62440 49784 62440 49784 0 wbs_dat_i[9]
rlabel metal2 26600 109830 26600 109830 0 wbs_dat_o[0]
rlabel metal2 91336 24206 91336 24206 0 wbs_dat_o[10]
rlabel metal4 328776 237771 328776 237771 0 wbs_dat_o[11]
rlabel metal3 329896 256354 329896 256354 0 wbs_dat_o[12]
rlabel metal3 199976 44520 199976 44520 0 wbs_dat_o[13]
rlabel metal5 329504 240750 329504 240750 0 wbs_dat_o[14]
rlabel metal2 119896 22526 119896 22526 0 wbs_dat_o[15]
rlabel metal3 329896 259938 329896 259938 0 wbs_dat_o[16]
rlabel metal4 326872 237857 326872 237857 0 wbs_dat_o[17]
rlabel metal5 329952 248310 329952 248310 0 wbs_dat_o[18]
rlabel metal3 329896 236544 329896 236544 0 wbs_dat_o[19]
rlabel metal2 34440 2310 34440 2310 0 wbs_dat_o[1]
rlabel metal2 327544 236376 327544 236376 0 wbs_dat_o[20]
rlabel metal3 331646 264712 331646 264712 0 wbs_dat_o[21]
rlabel metal4 329224 265590 329224 265590 0 wbs_dat_o[22]
rlabel metal3 331310 266504 331310 266504 0 wbs_dat_o[23]
rlabel metal3 330680 263816 330680 263816 0 wbs_dat_o[24]
rlabel metal3 334544 264040 334544 264040 0 wbs_dat_o[25]
rlabel metal2 281400 132832 281400 132832 0 wbs_dat_o[26]
rlabel metal2 327992 236992 327992 236992 0 wbs_dat_o[27]
rlabel metal2 194152 22862 194152 22862 0 wbs_dat_o[28]
rlabel metal2 329448 240912 329448 240912 0 wbs_dat_o[29]
rlabel metal2 331016 237496 331016 237496 0 wbs_dat_o[2]
rlabel metal3 333592 289128 333592 289128 0 wbs_dat_o[30]
rlabel metal3 334376 263816 334376 263816 0 wbs_dat_o[31]
rlabel metal4 289800 138936 289800 138936 0 wbs_dat_o[3]
rlabel metal4 288344 136151 288344 136151 0 wbs_dat_o[4]
rlabel metal4 286664 136528 286664 136528 0 wbs_dat_o[5]
rlabel metal2 68488 20958 68488 20958 0 wbs_dat_o[6]
rlabel metal2 74200 24262 74200 24262 0 wbs_dat_o[7]
rlabel metal2 285992 138320 285992 138320 0 wbs_dat_o[8]
rlabel metal4 286440 140605 286440 140605 0 wbs_dat_o[9]
rlabel metal3 333760 281400 333760 281400 0 wbs_stb_i
rlabel metal3 330736 287336 330736 287336 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
