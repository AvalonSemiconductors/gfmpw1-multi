magic
tech gf180mcuD
magscale 1 5
timestamp 1702241823
<< obsm1 >>
rect 672 1538 99288 108222
<< metal2 >>
rect 1568 109600 1624 110000
rect 4592 109600 4648 110000
rect 7616 109600 7672 110000
rect 10640 109600 10696 110000
rect 13664 109600 13720 110000
rect 16688 109600 16744 110000
rect 19712 109600 19768 110000
rect 22736 109600 22792 110000
rect 25760 109600 25816 110000
rect 28784 109600 28840 110000
rect 31808 109600 31864 110000
rect 34832 109600 34888 110000
rect 37856 109600 37912 110000
rect 40880 109600 40936 110000
rect 43904 109600 43960 110000
rect 46928 109600 46984 110000
rect 49952 109600 50008 110000
rect 52976 109600 53032 110000
rect 56000 109600 56056 110000
rect 59024 109600 59080 110000
rect 62048 109600 62104 110000
rect 65072 109600 65128 110000
rect 68096 109600 68152 110000
rect 71120 109600 71176 110000
rect 74144 109600 74200 110000
rect 77168 109600 77224 110000
rect 80192 109600 80248 110000
rect 83216 109600 83272 110000
rect 86240 109600 86296 110000
rect 89264 109600 89320 110000
rect 92288 109600 92344 110000
rect 95312 109600 95368 110000
rect 98336 109600 98392 110000
rect 1568 0 1624 400
rect 4592 0 4648 400
rect 7616 0 7672 400
rect 10640 0 10696 400
rect 13664 0 13720 400
rect 16688 0 16744 400
rect 19712 0 19768 400
rect 22736 0 22792 400
rect 25760 0 25816 400
rect 28784 0 28840 400
rect 31808 0 31864 400
rect 34832 0 34888 400
rect 37856 0 37912 400
rect 40880 0 40936 400
rect 43904 0 43960 400
rect 46928 0 46984 400
rect 49952 0 50008 400
rect 52976 0 53032 400
rect 56000 0 56056 400
rect 59024 0 59080 400
rect 62048 0 62104 400
rect 65072 0 65128 400
rect 68096 0 68152 400
rect 71120 0 71176 400
rect 74144 0 74200 400
rect 77168 0 77224 400
rect 80192 0 80248 400
rect 83216 0 83272 400
rect 86240 0 86296 400
rect 89264 0 89320 400
rect 92288 0 92344 400
rect 95312 0 95368 400
rect 98336 0 98392 400
<< obsm2 >>
rect 14 109570 1538 109600
rect 1654 109570 4562 109600
rect 4678 109570 7586 109600
rect 7702 109570 10610 109600
rect 10726 109570 13634 109600
rect 13750 109570 16658 109600
rect 16774 109570 19682 109600
rect 19798 109570 22706 109600
rect 22822 109570 25730 109600
rect 25846 109570 28754 109600
rect 28870 109570 31778 109600
rect 31894 109570 34802 109600
rect 34918 109570 37826 109600
rect 37942 109570 40850 109600
rect 40966 109570 43874 109600
rect 43990 109570 46898 109600
rect 47014 109570 49922 109600
rect 50038 109570 52946 109600
rect 53062 109570 55970 109600
rect 56086 109570 58994 109600
rect 59110 109570 62018 109600
rect 62134 109570 65042 109600
rect 65158 109570 68066 109600
rect 68182 109570 71090 109600
rect 71206 109570 74114 109600
rect 74230 109570 77138 109600
rect 77254 109570 80162 109600
rect 80278 109570 83186 109600
rect 83302 109570 86210 109600
rect 86326 109570 89234 109600
rect 89350 109570 92258 109600
rect 92374 109570 95282 109600
rect 95398 109570 98306 109600
rect 98422 109570 99386 109600
rect 14 430 99386 109570
rect 14 289 1538 430
rect 1654 289 4562 430
rect 4678 289 7586 430
rect 7702 289 10610 430
rect 10726 289 13634 430
rect 13750 289 16658 430
rect 16774 289 19682 430
rect 19798 289 22706 430
rect 22822 289 25730 430
rect 25846 289 28754 430
rect 28870 289 31778 430
rect 31894 289 34802 430
rect 34918 289 37826 430
rect 37942 289 40850 430
rect 40966 289 43874 430
rect 43990 289 46898 430
rect 47014 289 49922 430
rect 50038 289 52946 430
rect 53062 289 55970 430
rect 56086 289 58994 430
rect 59110 289 62018 430
rect 62134 289 65042 430
rect 65158 289 68066 430
rect 68182 289 71090 430
rect 71206 289 74114 430
rect 74230 289 77138 430
rect 77254 289 80162 430
rect 80278 289 83186 430
rect 83302 289 86210 430
rect 86326 289 89234 430
rect 89350 289 92258 430
rect 92374 289 95282 430
rect 95398 289 98306 430
rect 98422 289 99386 430
<< metal3 >>
rect 0 107296 400 107352
rect 0 104384 400 104440
rect 0 101472 400 101528
rect 0 98560 400 98616
rect 0 95648 400 95704
rect 0 92736 400 92792
rect 0 89824 400 89880
rect 0 86912 400 86968
rect 0 84000 400 84056
rect 0 81088 400 81144
rect 0 78176 400 78232
rect 0 75264 400 75320
rect 0 72352 400 72408
rect 0 69440 400 69496
rect 0 66528 400 66584
rect 0 63616 400 63672
rect 0 60704 400 60760
rect 0 57792 400 57848
rect 0 54880 400 54936
rect 0 51968 400 52024
rect 0 49056 400 49112
rect 0 46144 400 46200
rect 0 43232 400 43288
rect 0 40320 400 40376
rect 0 37408 400 37464
rect 0 34496 400 34552
rect 0 31584 400 31640
rect 0 28672 400 28728
rect 0 25760 400 25816
rect 0 22848 400 22904
rect 0 19936 400 19992
rect 0 17024 400 17080
rect 0 14112 400 14168
rect 0 11200 400 11256
rect 0 8288 400 8344
rect 0 5376 400 5432
rect 0 2464 400 2520
<< obsm3 >>
rect 9 107382 99391 108570
rect 430 107266 99391 107382
rect 9 104470 99391 107266
rect 430 104354 99391 104470
rect 9 101558 99391 104354
rect 430 101442 99391 101558
rect 9 98646 99391 101442
rect 430 98530 99391 98646
rect 9 95734 99391 98530
rect 430 95618 99391 95734
rect 9 92822 99391 95618
rect 430 92706 99391 92822
rect 9 89910 99391 92706
rect 430 89794 99391 89910
rect 9 86998 99391 89794
rect 430 86882 99391 86998
rect 9 84086 99391 86882
rect 430 83970 99391 84086
rect 9 81174 99391 83970
rect 430 81058 99391 81174
rect 9 78262 99391 81058
rect 430 78146 99391 78262
rect 9 75350 99391 78146
rect 430 75234 99391 75350
rect 9 72438 99391 75234
rect 430 72322 99391 72438
rect 9 69526 99391 72322
rect 430 69410 99391 69526
rect 9 66614 99391 69410
rect 430 66498 99391 66614
rect 9 63702 99391 66498
rect 430 63586 99391 63702
rect 9 60790 99391 63586
rect 430 60674 99391 60790
rect 9 57878 99391 60674
rect 430 57762 99391 57878
rect 9 54966 99391 57762
rect 430 54850 99391 54966
rect 9 52054 99391 54850
rect 430 51938 99391 52054
rect 9 49142 99391 51938
rect 430 49026 99391 49142
rect 9 46230 99391 49026
rect 430 46114 99391 46230
rect 9 43318 99391 46114
rect 430 43202 99391 43318
rect 9 40406 99391 43202
rect 430 40290 99391 40406
rect 9 37494 99391 40290
rect 430 37378 99391 37494
rect 9 34582 99391 37378
rect 430 34466 99391 34582
rect 9 31670 99391 34466
rect 430 31554 99391 31670
rect 9 28758 99391 31554
rect 430 28642 99391 28758
rect 9 25846 99391 28642
rect 430 25730 99391 25846
rect 9 22934 99391 25730
rect 430 22818 99391 22934
rect 9 20022 99391 22818
rect 430 19906 99391 20022
rect 9 17110 99391 19906
rect 430 16994 99391 17110
rect 9 14198 99391 16994
rect 430 14082 99391 14198
rect 9 11286 99391 14082
rect 430 11170 99391 11286
rect 9 8374 99391 11170
rect 430 8258 99391 8374
rect 9 5462 99391 8258
rect 430 5346 99391 5462
rect 9 2550 99391 5346
rect 430 2434 99391 2550
rect 9 294 99391 2434
<< metal4 >>
rect 2224 1538 2384 108222
rect 9904 1538 10064 108222
rect 17584 1538 17744 108222
rect 25264 1538 25424 108222
rect 32944 1538 33104 108222
rect 40624 1538 40784 108222
rect 48304 1538 48464 108222
rect 55984 1538 56144 108222
rect 63664 1538 63824 108222
rect 71344 1538 71504 108222
rect 79024 1538 79184 108222
rect 86704 1538 86864 108222
rect 94384 1538 94544 108222
<< obsm4 >>
rect 1134 108252 98938 108463
rect 1134 1508 2194 108252
rect 2414 1508 9874 108252
rect 10094 1508 17554 108252
rect 17774 1508 25234 108252
rect 25454 1508 32914 108252
rect 33134 1508 40594 108252
rect 40814 1508 48274 108252
rect 48494 1508 55954 108252
rect 56174 1508 63634 108252
rect 63854 1508 71314 108252
rect 71534 1508 78994 108252
rect 79214 1508 86674 108252
rect 86894 1508 94354 108252
rect 94574 1508 98938 108252
rect 1134 289 98938 1508
<< labels >>
rlabel metal3 s 0 8288 400 8344 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 11200 400 11256 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 0 14112 400 14168 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 0 43232 400 43288 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 0 46144 400 46200 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 49056 400 49112 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 0 51968 400 52024 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 0 54880 400 54936 6 io_in[14]
port 8 nsew signal input
rlabel metal3 s 0 57792 400 57848 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 60704 400 60760 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 0 63616 400 63672 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 66528 400 66584 6 io_in[18]
port 12 nsew signal input
rlabel metal3 s 0 69440 400 69496 6 io_in[19]
port 13 nsew signal input
rlabel metal3 s 0 17024 400 17080 6 io_in[1]
port 14 nsew signal input
rlabel metal3 s 0 72352 400 72408 6 io_in[20]
port 15 nsew signal input
rlabel metal3 s 0 75264 400 75320 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 78176 400 78232 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 81088 400 81144 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 0 84000 400 84056 6 io_in[24]
port 19 nsew signal input
rlabel metal3 s 0 86912 400 86968 6 io_in[25]
port 20 nsew signal input
rlabel metal3 s 0 89824 400 89880 6 io_in[26]
port 21 nsew signal input
rlabel metal3 s 0 92736 400 92792 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 95648 400 95704 6 io_in[28]
port 23 nsew signal input
rlabel metal3 s 0 98560 400 98616 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 19936 400 19992 6 io_in[2]
port 25 nsew signal input
rlabel metal3 s 0 101472 400 101528 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 104384 400 104440 6 io_in[31]
port 27 nsew signal input
rlabel metal3 s 0 107296 400 107352 6 io_in[32]
port 28 nsew signal input
rlabel metal3 s 0 22848 400 22904 6 io_in[3]
port 29 nsew signal input
rlabel metal3 s 0 25760 400 25816 6 io_in[4]
port 30 nsew signal input
rlabel metal3 s 0 28672 400 28728 6 io_in[5]
port 31 nsew signal input
rlabel metal3 s 0 31584 400 31640 6 io_in[6]
port 32 nsew signal input
rlabel metal3 s 0 34496 400 34552 6 io_in[7]
port 33 nsew signal input
rlabel metal3 s 0 37408 400 37464 6 io_in[8]
port 34 nsew signal input
rlabel metal3 s 0 40320 400 40376 6 io_in[9]
port 35 nsew signal input
rlabel metal2 s 1568 109600 1624 110000 6 io_oeb[0]
port 36 nsew signal output
rlabel metal2 s 31808 109600 31864 110000 6 io_oeb[10]
port 37 nsew signal output
rlabel metal2 s 34832 109600 34888 110000 6 io_oeb[11]
port 38 nsew signal output
rlabel metal2 s 37856 109600 37912 110000 6 io_oeb[12]
port 39 nsew signal output
rlabel metal2 s 40880 109600 40936 110000 6 io_oeb[13]
port 40 nsew signal output
rlabel metal2 s 43904 109600 43960 110000 6 io_oeb[14]
port 41 nsew signal output
rlabel metal2 s 46928 109600 46984 110000 6 io_oeb[15]
port 42 nsew signal output
rlabel metal2 s 49952 109600 50008 110000 6 io_oeb[16]
port 43 nsew signal output
rlabel metal2 s 52976 109600 53032 110000 6 io_oeb[17]
port 44 nsew signal output
rlabel metal2 s 56000 109600 56056 110000 6 io_oeb[18]
port 45 nsew signal output
rlabel metal2 s 59024 109600 59080 110000 6 io_oeb[19]
port 46 nsew signal output
rlabel metal2 s 4592 109600 4648 110000 6 io_oeb[1]
port 47 nsew signal output
rlabel metal2 s 62048 109600 62104 110000 6 io_oeb[20]
port 48 nsew signal output
rlabel metal2 s 65072 109600 65128 110000 6 io_oeb[21]
port 49 nsew signal output
rlabel metal2 s 68096 109600 68152 110000 6 io_oeb[22]
port 50 nsew signal output
rlabel metal2 s 71120 109600 71176 110000 6 io_oeb[23]
port 51 nsew signal output
rlabel metal2 s 74144 109600 74200 110000 6 io_oeb[24]
port 52 nsew signal output
rlabel metal2 s 77168 109600 77224 110000 6 io_oeb[25]
port 53 nsew signal output
rlabel metal2 s 80192 109600 80248 110000 6 io_oeb[26]
port 54 nsew signal output
rlabel metal2 s 83216 109600 83272 110000 6 io_oeb[27]
port 55 nsew signal output
rlabel metal2 s 86240 109600 86296 110000 6 io_oeb[28]
port 56 nsew signal output
rlabel metal2 s 89264 109600 89320 110000 6 io_oeb[29]
port 57 nsew signal output
rlabel metal2 s 7616 109600 7672 110000 6 io_oeb[2]
port 58 nsew signal output
rlabel metal2 s 92288 109600 92344 110000 6 io_oeb[30]
port 59 nsew signal output
rlabel metal2 s 95312 109600 95368 110000 6 io_oeb[31]
port 60 nsew signal output
rlabel metal2 s 98336 109600 98392 110000 6 io_oeb[32]
port 61 nsew signal output
rlabel metal2 s 10640 109600 10696 110000 6 io_oeb[3]
port 62 nsew signal output
rlabel metal2 s 13664 109600 13720 110000 6 io_oeb[4]
port 63 nsew signal output
rlabel metal2 s 16688 109600 16744 110000 6 io_oeb[5]
port 64 nsew signal output
rlabel metal2 s 19712 109600 19768 110000 6 io_oeb[6]
port 65 nsew signal output
rlabel metal2 s 22736 109600 22792 110000 6 io_oeb[7]
port 66 nsew signal output
rlabel metal2 s 25760 109600 25816 110000 6 io_oeb[8]
port 67 nsew signal output
rlabel metal2 s 28784 109600 28840 110000 6 io_oeb[9]
port 68 nsew signal output
rlabel metal2 s 1568 0 1624 400 6 io_out[0]
port 69 nsew signal output
rlabel metal2 s 31808 0 31864 400 6 io_out[10]
port 70 nsew signal output
rlabel metal2 s 34832 0 34888 400 6 io_out[11]
port 71 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 io_out[12]
port 72 nsew signal output
rlabel metal2 s 40880 0 40936 400 6 io_out[13]
port 73 nsew signal output
rlabel metal2 s 43904 0 43960 400 6 io_out[14]
port 74 nsew signal output
rlabel metal2 s 46928 0 46984 400 6 io_out[15]
port 75 nsew signal output
rlabel metal2 s 49952 0 50008 400 6 io_out[16]
port 76 nsew signal output
rlabel metal2 s 52976 0 53032 400 6 io_out[17]
port 77 nsew signal output
rlabel metal2 s 56000 0 56056 400 6 io_out[18]
port 78 nsew signal output
rlabel metal2 s 59024 0 59080 400 6 io_out[19]
port 79 nsew signal output
rlabel metal2 s 4592 0 4648 400 6 io_out[1]
port 80 nsew signal output
rlabel metal2 s 62048 0 62104 400 6 io_out[20]
port 81 nsew signal output
rlabel metal2 s 65072 0 65128 400 6 io_out[21]
port 82 nsew signal output
rlabel metal2 s 68096 0 68152 400 6 io_out[22]
port 83 nsew signal output
rlabel metal2 s 71120 0 71176 400 6 io_out[23]
port 84 nsew signal output
rlabel metal2 s 74144 0 74200 400 6 io_out[24]
port 85 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 io_out[25]
port 86 nsew signal output
rlabel metal2 s 80192 0 80248 400 6 io_out[26]
port 87 nsew signal output
rlabel metal2 s 83216 0 83272 400 6 io_out[27]
port 88 nsew signal output
rlabel metal2 s 86240 0 86296 400 6 io_out[28]
port 89 nsew signal output
rlabel metal2 s 89264 0 89320 400 6 io_out[29]
port 90 nsew signal output
rlabel metal2 s 7616 0 7672 400 6 io_out[2]
port 91 nsew signal output
rlabel metal2 s 92288 0 92344 400 6 io_out[30]
port 92 nsew signal output
rlabel metal2 s 95312 0 95368 400 6 io_out[31]
port 93 nsew signal output
rlabel metal2 s 98336 0 98392 400 6 io_out[32]
port 94 nsew signal output
rlabel metal2 s 10640 0 10696 400 6 io_out[3]
port 95 nsew signal output
rlabel metal2 s 13664 0 13720 400 6 io_out[4]
port 96 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 io_out[5]
port 97 nsew signal output
rlabel metal2 s 19712 0 19768 400 6 io_out[6]
port 98 nsew signal output
rlabel metal2 s 22736 0 22792 400 6 io_out[7]
port 99 nsew signal output
rlabel metal2 s 25760 0 25816 400 6 io_out[8]
port 100 nsew signal output
rlabel metal2 s 28784 0 28840 400 6 io_out[9]
port 101 nsew signal output
rlabel metal3 s 0 5376 400 5432 6 rst_n
port 102 nsew signal input
rlabel metal4 s 2224 1538 2384 108222 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 108222 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 108222 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 108222 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 108222 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 108222 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 108222 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 108222 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 108222 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 108222 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 108222 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 108222 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 108222 6 vss
port 104 nsew ground bidirectional
rlabel metal3 s 0 2464 400 2520 6 wb_clk_i
port 105 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 37709864
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_tholin_riscv/runs/23_12_10_21_06/results/signoff/wrapped_tholin_riscv.magic.gds
string GDS_START 552198
<< end >>

