magic
tech gf180mcuD
magscale 1 10
timestamp 1702046418
<< metal1 >>
rect 1344 22762 24640 22796
rect 1344 22710 4126 22762
rect 4178 22710 4230 22762
rect 4282 22710 4334 22762
rect 4386 22710 9950 22762
rect 10002 22710 10054 22762
rect 10106 22710 10158 22762
rect 10210 22710 15774 22762
rect 15826 22710 15878 22762
rect 15930 22710 15982 22762
rect 16034 22710 21598 22762
rect 21650 22710 21702 22762
rect 21754 22710 21806 22762
rect 21858 22710 24640 22762
rect 1344 22676 24640 22710
rect 22430 22594 22482 22606
rect 22430 22530 22482 22542
rect 12686 22482 12738 22494
rect 12686 22418 12738 22430
rect 19630 22370 19682 22382
rect 13346 22318 13358 22370
rect 13410 22318 13422 22370
rect 19954 22318 19966 22370
rect 20018 22318 20030 22370
rect 20850 22318 20862 22370
rect 20914 22318 20926 22370
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 19630 22306 19682 22318
rect 13134 22146 13186 22158
rect 13134 22082 13186 22094
rect 18734 22146 18786 22158
rect 18734 22082 18786 22094
rect 19182 22146 19234 22158
rect 19182 22082 19234 22094
rect 20190 22146 20242 22158
rect 20190 22082 20242 22094
rect 21086 22146 21138 22158
rect 21086 22082 21138 22094
rect 1344 21978 24800 22012
rect 1344 21926 7038 21978
rect 7090 21926 7142 21978
rect 7194 21926 7246 21978
rect 7298 21926 12862 21978
rect 12914 21926 12966 21978
rect 13018 21926 13070 21978
rect 13122 21926 18686 21978
rect 18738 21926 18790 21978
rect 18842 21926 18894 21978
rect 18946 21926 24510 21978
rect 24562 21926 24614 21978
rect 24666 21926 24718 21978
rect 24770 21926 24800 21978
rect 1344 21892 24800 21926
rect 8206 21810 8258 21822
rect 8206 21746 8258 21758
rect 17502 21698 17554 21710
rect 17502 21634 17554 21646
rect 16270 21586 16322 21598
rect 5058 21534 5070 21586
rect 5122 21534 5134 21586
rect 8418 21534 8430 21586
rect 8482 21534 8494 21586
rect 9650 21534 9662 21586
rect 9714 21534 9726 21586
rect 13010 21534 13022 21586
rect 13074 21534 13086 21586
rect 16270 21522 16322 21534
rect 17390 21586 17442 21598
rect 17938 21534 17950 21586
rect 18002 21534 18014 21586
rect 21186 21534 21198 21586
rect 21250 21534 21262 21586
rect 17390 21522 17442 21534
rect 5730 21422 5742 21474
rect 5794 21422 5806 21474
rect 7858 21422 7870 21474
rect 7922 21422 7934 21474
rect 10434 21422 10446 21474
rect 10498 21422 10510 21474
rect 12562 21422 12574 21474
rect 12626 21422 12638 21474
rect 13682 21422 13694 21474
rect 13746 21422 13758 21474
rect 15810 21422 15822 21474
rect 15874 21422 15886 21474
rect 18722 21422 18734 21474
rect 18786 21422 18798 21474
rect 20850 21422 20862 21474
rect 20914 21422 20926 21474
rect 21970 21422 21982 21474
rect 22034 21422 22046 21474
rect 24098 21422 24110 21474
rect 24162 21422 24174 21474
rect 17502 21362 17554 21374
rect 17502 21298 17554 21310
rect 1344 21194 24640 21228
rect 1344 21142 4126 21194
rect 4178 21142 4230 21194
rect 4282 21142 4334 21194
rect 4386 21142 9950 21194
rect 10002 21142 10054 21194
rect 10106 21142 10158 21194
rect 10210 21142 15774 21194
rect 15826 21142 15878 21194
rect 15930 21142 15982 21194
rect 16034 21142 21598 21194
rect 21650 21142 21702 21194
rect 21754 21142 21806 21194
rect 21858 21142 24640 21194
rect 1344 21108 24640 21142
rect 8866 20974 8878 21026
rect 8930 20974 8942 21026
rect 20414 20914 20466 20926
rect 5058 20862 5070 20914
rect 5122 20862 5134 20914
rect 18498 20862 18510 20914
rect 18562 20862 18574 20914
rect 19618 20862 19630 20914
rect 19682 20862 19694 20914
rect 20414 20850 20466 20862
rect 8094 20802 8146 20814
rect 23214 20802 23266 20814
rect 2258 20750 2270 20802
rect 2322 20750 2334 20802
rect 8642 20750 8654 20802
rect 8706 20750 8718 20802
rect 9314 20750 9326 20802
rect 9378 20750 9390 20802
rect 15586 20750 15598 20802
rect 15650 20750 15662 20802
rect 19506 20750 19518 20802
rect 19570 20750 19582 20802
rect 21970 20750 21982 20802
rect 22034 20750 22046 20802
rect 22418 20750 22430 20802
rect 22482 20750 22494 20802
rect 23538 20750 23550 20802
rect 23602 20750 23614 20802
rect 8094 20738 8146 20750
rect 23214 20738 23266 20750
rect 7646 20690 7698 20702
rect 9886 20690 9938 20702
rect 2930 20638 2942 20690
rect 2994 20638 3006 20690
rect 8306 20638 8318 20690
rect 8370 20638 8382 20690
rect 7646 20626 7698 20638
rect 9886 20626 9938 20638
rect 10446 20690 10498 20702
rect 19966 20690 20018 20702
rect 16370 20638 16382 20690
rect 16434 20638 16446 20690
rect 10446 20626 10498 20638
rect 19966 20626 20018 20638
rect 20302 20690 20354 20702
rect 20302 20626 20354 20638
rect 21758 20690 21810 20702
rect 21758 20626 21810 20638
rect 24110 20690 24162 20702
rect 24110 20626 24162 20638
rect 7758 20578 7810 20590
rect 7758 20514 7810 20526
rect 9998 20578 10050 20590
rect 9998 20514 10050 20526
rect 10222 20578 10274 20590
rect 10222 20514 10274 20526
rect 10558 20578 10610 20590
rect 10558 20514 10610 20526
rect 10782 20578 10834 20590
rect 10782 20514 10834 20526
rect 20526 20578 20578 20590
rect 20526 20514 20578 20526
rect 21534 20578 21586 20590
rect 21534 20514 21586 20526
rect 1344 20410 24800 20444
rect 1344 20358 7038 20410
rect 7090 20358 7142 20410
rect 7194 20358 7246 20410
rect 7298 20358 12862 20410
rect 12914 20358 12966 20410
rect 13018 20358 13070 20410
rect 13122 20358 18686 20410
rect 18738 20358 18790 20410
rect 18842 20358 18894 20410
rect 18946 20358 24510 20410
rect 24562 20358 24614 20410
rect 24666 20358 24718 20410
rect 24770 20358 24800 20410
rect 1344 20324 24800 20358
rect 6750 20242 6802 20254
rect 6750 20178 6802 20190
rect 8878 20242 8930 20254
rect 8878 20178 8930 20190
rect 13918 20242 13970 20254
rect 13918 20178 13970 20190
rect 9550 20130 9602 20142
rect 4946 20078 4958 20130
rect 5010 20078 5022 20130
rect 9550 20066 9602 20078
rect 9998 20130 10050 20142
rect 9998 20066 10050 20078
rect 11342 20130 11394 20142
rect 11342 20066 11394 20078
rect 12910 20130 12962 20142
rect 12910 20066 12962 20078
rect 14142 20130 14194 20142
rect 16494 20130 16546 20142
rect 14914 20078 14926 20130
rect 14978 20078 14990 20130
rect 14142 20066 14194 20078
rect 16494 20066 16546 20078
rect 16606 20130 16658 20142
rect 16606 20066 16658 20078
rect 18734 20130 18786 20142
rect 18734 20066 18786 20078
rect 19406 20130 19458 20142
rect 19406 20066 19458 20078
rect 19854 20130 19906 20142
rect 19854 20066 19906 20078
rect 20414 20130 20466 20142
rect 20414 20066 20466 20078
rect 20638 20130 20690 20142
rect 20638 20066 20690 20078
rect 21310 20130 21362 20142
rect 21310 20066 21362 20078
rect 21870 20130 21922 20142
rect 21870 20066 21922 20078
rect 22094 20130 22146 20142
rect 22094 20066 22146 20078
rect 22430 20130 22482 20142
rect 22430 20066 22482 20078
rect 7982 20018 8034 20030
rect 4386 19966 4398 20018
rect 4450 19966 4462 20018
rect 7746 19966 7758 20018
rect 7810 19966 7822 20018
rect 7982 19954 8034 19966
rect 8990 20018 9042 20030
rect 11230 20018 11282 20030
rect 9762 19966 9774 20018
rect 9826 19966 9838 20018
rect 8990 19954 9042 19966
rect 11230 19954 11282 19966
rect 11566 20018 11618 20030
rect 11566 19954 11618 19966
rect 13134 20018 13186 20030
rect 13134 19954 13186 19966
rect 13582 20018 13634 20030
rect 13582 19954 13634 19966
rect 13806 20018 13858 20030
rect 13806 19954 13858 19966
rect 14254 20018 14306 20030
rect 14254 19954 14306 19966
rect 15262 20018 15314 20030
rect 16830 20018 16882 20030
rect 19630 20018 19682 20030
rect 16034 19966 16046 20018
rect 16098 19966 16110 20018
rect 18162 19966 18174 20018
rect 18226 19966 18238 20018
rect 15262 19954 15314 19966
rect 16830 19954 16882 19966
rect 19630 19954 19682 19966
rect 19966 20018 20018 20030
rect 22766 20018 22818 20030
rect 21074 19966 21086 20018
rect 21138 19966 21150 20018
rect 21634 19966 21646 20018
rect 21698 19966 21710 20018
rect 19966 19954 20018 19966
rect 22766 19954 22818 19966
rect 23214 20018 23266 20030
rect 23650 19966 23662 20018
rect 23714 19966 23726 20018
rect 23214 19954 23266 19966
rect 6638 19906 6690 19918
rect 4498 19854 4510 19906
rect 4562 19854 4574 19906
rect 6638 19842 6690 19854
rect 7086 19906 7138 19918
rect 7086 19842 7138 19854
rect 9886 19906 9938 19918
rect 9886 19842 9938 19854
rect 13358 19906 13410 19918
rect 17950 19906 18002 19918
rect 24110 19906 24162 19918
rect 16482 19854 16494 19906
rect 16546 19854 16558 19906
rect 20290 19854 20302 19906
rect 20354 19854 20366 19906
rect 21970 19854 21982 19906
rect 22034 19854 22046 19906
rect 13358 19842 13410 19854
rect 17950 19842 18002 19854
rect 24110 19842 24162 19854
rect 8878 19794 8930 19806
rect 8878 19730 8930 19742
rect 17838 19794 17890 19806
rect 17838 19730 17890 19742
rect 1344 19626 24640 19660
rect 1344 19574 4126 19626
rect 4178 19574 4230 19626
rect 4282 19574 4334 19626
rect 4386 19574 9950 19626
rect 10002 19574 10054 19626
rect 10106 19574 10158 19626
rect 10210 19574 15774 19626
rect 15826 19574 15878 19626
rect 15930 19574 15982 19626
rect 16034 19574 21598 19626
rect 21650 19574 21702 19626
rect 21754 19574 21806 19626
rect 21858 19574 24640 19626
rect 1344 19540 24640 19574
rect 7534 19458 7586 19470
rect 7534 19394 7586 19406
rect 11790 19458 11842 19470
rect 11790 19394 11842 19406
rect 11902 19458 11954 19470
rect 11902 19394 11954 19406
rect 12574 19458 12626 19470
rect 12574 19394 12626 19406
rect 16718 19458 16770 19470
rect 21646 19458 21698 19470
rect 20402 19406 20414 19458
rect 20466 19455 20478 19458
rect 20850 19455 20862 19458
rect 20466 19409 20862 19455
rect 20466 19406 20478 19409
rect 20850 19406 20862 19409
rect 20914 19406 20926 19458
rect 16718 19394 16770 19406
rect 21646 19394 21698 19406
rect 13806 19346 13858 19358
rect 13806 19282 13858 19294
rect 15486 19346 15538 19358
rect 20526 19346 20578 19358
rect 17938 19294 17950 19346
rect 18002 19294 18014 19346
rect 20066 19294 20078 19346
rect 20130 19294 20142 19346
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 22866 19294 22878 19346
rect 22930 19294 22942 19346
rect 15486 19282 15538 19294
rect 20526 19282 20578 19294
rect 7422 19234 7474 19246
rect 8094 19234 8146 19246
rect 4386 19182 4398 19234
rect 4450 19182 4462 19234
rect 7858 19182 7870 19234
rect 7922 19182 7934 19234
rect 7422 19170 7474 19182
rect 8094 19170 8146 19182
rect 8206 19234 8258 19246
rect 8206 19170 8258 19182
rect 9102 19234 9154 19246
rect 9102 19170 9154 19182
rect 10670 19234 10722 19246
rect 10670 19170 10722 19182
rect 10894 19234 10946 19246
rect 10894 19170 10946 19182
rect 11902 19234 11954 19246
rect 11902 19170 11954 19182
rect 12350 19234 12402 19246
rect 12350 19170 12402 19182
rect 13918 19234 13970 19246
rect 13918 19170 13970 19182
rect 14366 19234 14418 19246
rect 14366 19170 14418 19182
rect 14590 19234 14642 19246
rect 14590 19170 14642 19182
rect 14814 19234 14866 19246
rect 14814 19170 14866 19182
rect 14926 19234 14978 19246
rect 14926 19170 14978 19182
rect 15374 19234 15426 19246
rect 15374 19170 15426 19182
rect 16942 19234 16994 19246
rect 17266 19182 17278 19234
rect 17330 19182 17342 19234
rect 22978 19182 22990 19234
rect 23042 19182 23054 19234
rect 16942 19170 16994 19182
rect 3278 19122 3330 19134
rect 9438 19122 9490 19134
rect 3938 19070 3950 19122
rect 4002 19070 4014 19122
rect 4274 19070 4286 19122
rect 4338 19070 4350 19122
rect 8642 19070 8654 19122
rect 8706 19070 8718 19122
rect 3278 19058 3330 19070
rect 9438 19058 9490 19070
rect 9774 19122 9826 19134
rect 9774 19058 9826 19070
rect 10110 19122 10162 19134
rect 10110 19058 10162 19070
rect 10334 19122 10386 19134
rect 10334 19058 10386 19070
rect 21422 19122 21474 19134
rect 21422 19058 21474 19070
rect 21982 19122 22034 19134
rect 21982 19058 22034 19070
rect 23662 19122 23714 19134
rect 23662 19058 23714 19070
rect 9326 19010 9378 19022
rect 9326 18946 9378 18958
rect 9998 19010 10050 19022
rect 14478 19010 14530 19022
rect 11218 18958 11230 19010
rect 11282 18958 11294 19010
rect 9998 18946 10050 18958
rect 14478 18946 14530 18958
rect 16382 19010 16434 19022
rect 16382 18946 16434 18958
rect 16606 19010 16658 19022
rect 16606 18946 16658 18958
rect 22094 19010 22146 19022
rect 22094 18946 22146 18958
rect 22206 19010 22258 19022
rect 22206 18946 22258 18958
rect 24110 19010 24162 19022
rect 24110 18946 24162 18958
rect 1344 18842 24800 18876
rect 1344 18790 7038 18842
rect 7090 18790 7142 18842
rect 7194 18790 7246 18842
rect 7298 18790 12862 18842
rect 12914 18790 12966 18842
rect 13018 18790 13070 18842
rect 13122 18790 18686 18842
rect 18738 18790 18790 18842
rect 18842 18790 18894 18842
rect 18946 18790 24510 18842
rect 24562 18790 24614 18842
rect 24666 18790 24718 18842
rect 24770 18790 24800 18842
rect 1344 18756 24800 18790
rect 11118 18674 11170 18686
rect 11118 18610 11170 18622
rect 11342 18674 11394 18686
rect 11342 18610 11394 18622
rect 14254 18674 14306 18686
rect 14254 18610 14306 18622
rect 14366 18674 14418 18686
rect 14366 18610 14418 18622
rect 11566 18562 11618 18574
rect 14142 18562 14194 18574
rect 5170 18510 5182 18562
rect 5234 18510 5246 18562
rect 7746 18510 7758 18562
rect 7810 18510 7822 18562
rect 12226 18510 12238 18562
rect 12290 18510 12302 18562
rect 12562 18510 12574 18562
rect 12626 18510 12638 18562
rect 11566 18498 11618 18510
rect 14142 18498 14194 18510
rect 15262 18562 15314 18574
rect 17378 18510 17390 18562
rect 17442 18510 17454 18562
rect 15262 18498 15314 18510
rect 4958 18450 5010 18462
rect 6862 18450 6914 18462
rect 1810 18398 1822 18450
rect 1874 18398 1886 18450
rect 5506 18398 5518 18450
rect 5570 18398 5582 18450
rect 6402 18398 6414 18450
rect 6466 18398 6478 18450
rect 4958 18386 5010 18398
rect 6862 18386 6914 18398
rect 7198 18450 7250 18462
rect 8430 18450 8482 18462
rect 7970 18398 7982 18450
rect 8034 18398 8046 18450
rect 7198 18386 7250 18398
rect 8430 18386 8482 18398
rect 8990 18450 9042 18462
rect 12910 18450 12962 18462
rect 10770 18398 10782 18450
rect 10834 18398 10846 18450
rect 12002 18398 12014 18450
rect 12066 18398 12078 18450
rect 8990 18386 9042 18398
rect 12910 18386 12962 18398
rect 14814 18450 14866 18462
rect 14814 18386 14866 18398
rect 15150 18450 15202 18462
rect 19966 18450 20018 18462
rect 17602 18398 17614 18450
rect 17666 18398 17678 18450
rect 19170 18398 19182 18450
rect 19234 18398 19246 18450
rect 15150 18386 15202 18398
rect 19966 18386 20018 18398
rect 20078 18450 20130 18462
rect 24110 18450 24162 18462
rect 23538 18398 23550 18450
rect 23602 18398 23614 18450
rect 20078 18386 20130 18398
rect 24110 18386 24162 18398
rect 9774 18338 9826 18350
rect 2482 18286 2494 18338
rect 2546 18286 2558 18338
rect 4610 18286 4622 18338
rect 4674 18286 4686 18338
rect 9774 18274 9826 18286
rect 19406 18338 19458 18350
rect 19406 18274 19458 18286
rect 20414 18338 20466 18350
rect 20738 18286 20750 18338
rect 20802 18286 20814 18338
rect 22866 18286 22878 18338
rect 22930 18286 22942 18338
rect 20414 18274 20466 18286
rect 4846 18226 4898 18238
rect 4846 18162 4898 18174
rect 11006 18226 11058 18238
rect 11006 18162 11058 18174
rect 15038 18226 15090 18238
rect 15038 18162 15090 18174
rect 19518 18226 19570 18238
rect 19518 18162 19570 18174
rect 20302 18226 20354 18238
rect 20302 18162 20354 18174
rect 1344 18058 24640 18092
rect 1344 18006 4126 18058
rect 4178 18006 4230 18058
rect 4282 18006 4334 18058
rect 4386 18006 9950 18058
rect 10002 18006 10054 18058
rect 10106 18006 10158 18058
rect 10210 18006 15774 18058
rect 15826 18006 15878 18058
rect 15930 18006 15982 18058
rect 16034 18006 21598 18058
rect 21650 18006 21702 18058
rect 21754 18006 21806 18058
rect 21858 18006 24640 18058
rect 1344 17972 24640 18006
rect 3614 17890 3666 17902
rect 3614 17826 3666 17838
rect 9550 17890 9602 17902
rect 9550 17826 9602 17838
rect 14366 17890 14418 17902
rect 14366 17826 14418 17838
rect 16494 17890 16546 17902
rect 20526 17890 20578 17902
rect 20178 17838 20190 17890
rect 20242 17838 20254 17890
rect 16494 17826 16546 17838
rect 20526 17826 20578 17838
rect 3838 17778 3890 17790
rect 9326 17778 9378 17790
rect 12014 17778 12066 17790
rect 5618 17726 5630 17778
rect 5682 17726 5694 17778
rect 10882 17726 10894 17778
rect 10946 17726 10958 17778
rect 3838 17714 3890 17726
rect 9326 17714 9378 17726
rect 12014 17714 12066 17726
rect 15934 17778 15986 17790
rect 15934 17714 15986 17726
rect 20750 17778 20802 17790
rect 21970 17726 21982 17778
rect 22034 17726 22046 17778
rect 20750 17714 20802 17726
rect 4398 17666 4450 17678
rect 11342 17666 11394 17678
rect 2930 17614 2942 17666
rect 2994 17614 3006 17666
rect 6738 17614 6750 17666
rect 6802 17614 6814 17666
rect 7186 17614 7198 17666
rect 7250 17614 7262 17666
rect 8754 17614 8766 17666
rect 8818 17614 8830 17666
rect 4398 17602 4450 17614
rect 11342 17602 11394 17614
rect 16158 17666 16210 17678
rect 16158 17602 16210 17614
rect 16830 17666 16882 17678
rect 16830 17602 16882 17614
rect 17166 17666 17218 17678
rect 19182 17666 19234 17678
rect 18050 17614 18062 17666
rect 18114 17614 18126 17666
rect 22306 17614 22318 17666
rect 22370 17614 22382 17666
rect 24098 17614 24110 17666
rect 24162 17614 24174 17666
rect 17166 17602 17218 17614
rect 19182 17602 19234 17614
rect 14478 17554 14530 17566
rect 8530 17502 8542 17554
rect 8594 17502 8606 17554
rect 14478 17490 14530 17502
rect 16942 17554 16994 17566
rect 16942 17490 16994 17502
rect 22766 17554 22818 17566
rect 22766 17490 22818 17502
rect 2382 17442 2434 17454
rect 4286 17442 4338 17454
rect 11902 17442 11954 17454
rect 3266 17390 3278 17442
rect 3330 17390 3342 17442
rect 9874 17390 9886 17442
rect 9938 17390 9950 17442
rect 2382 17378 2434 17390
rect 4286 17378 4338 17390
rect 11902 17378 11954 17390
rect 14366 17442 14418 17454
rect 23886 17442 23938 17454
rect 18274 17390 18286 17442
rect 18338 17390 18350 17442
rect 19506 17390 19518 17442
rect 19570 17390 19582 17442
rect 14366 17378 14418 17390
rect 23886 17378 23938 17390
rect 1344 17274 24800 17308
rect 1344 17222 7038 17274
rect 7090 17222 7142 17274
rect 7194 17222 7246 17274
rect 7298 17222 12862 17274
rect 12914 17222 12966 17274
rect 13018 17222 13070 17274
rect 13122 17222 18686 17274
rect 18738 17222 18790 17274
rect 18842 17222 18894 17274
rect 18946 17222 24510 17274
rect 24562 17222 24614 17274
rect 24666 17222 24718 17274
rect 24770 17222 24800 17274
rect 1344 17188 24800 17222
rect 2046 17106 2098 17118
rect 2046 17042 2098 17054
rect 4398 17106 4450 17118
rect 16146 17054 16158 17106
rect 16210 17054 16222 17106
rect 23090 17054 23102 17106
rect 23154 17054 23166 17106
rect 4398 17042 4450 17054
rect 1934 16994 1986 17006
rect 1934 16930 1986 16942
rect 3054 16994 3106 17006
rect 3054 16930 3106 16942
rect 3166 16994 3218 17006
rect 3166 16930 3218 16942
rect 7870 16994 7922 17006
rect 14254 16994 14306 17006
rect 9650 16942 9662 16994
rect 9714 16942 9726 16994
rect 7870 16930 7922 16942
rect 14254 16930 14306 16942
rect 14366 16994 14418 17006
rect 14802 16942 14814 16994
rect 14866 16942 14878 16994
rect 16258 16942 16270 16994
rect 16322 16942 16334 16994
rect 20626 16942 20638 16994
rect 20690 16942 20702 16994
rect 14366 16930 14418 16942
rect 6302 16882 6354 16894
rect 23662 16882 23714 16894
rect 4722 16830 4734 16882
rect 4786 16830 4798 16882
rect 10994 16830 11006 16882
rect 11058 16830 11070 16882
rect 14690 16830 14702 16882
rect 14754 16830 14766 16882
rect 15698 16830 15710 16882
rect 15762 16830 15774 16882
rect 17378 16830 17390 16882
rect 17442 16830 17454 16882
rect 23426 16830 23438 16882
rect 23490 16830 23502 16882
rect 6302 16818 6354 16830
rect 23662 16818 23714 16830
rect 23886 16882 23938 16894
rect 23886 16818 23938 16830
rect 24222 16882 24274 16894
rect 24222 16818 24274 16830
rect 7310 16770 7362 16782
rect 3938 16718 3950 16770
rect 4002 16718 4014 16770
rect 6738 16718 6750 16770
rect 6802 16718 6814 16770
rect 7310 16706 7362 16718
rect 10110 16770 10162 16782
rect 10110 16706 10162 16718
rect 10334 16770 10386 16782
rect 11778 16718 11790 16770
rect 11842 16718 11854 16770
rect 13906 16718 13918 16770
rect 13970 16718 13982 16770
rect 10334 16706 10386 16718
rect 3054 16658 3106 16670
rect 3054 16594 3106 16606
rect 5742 16658 5794 16670
rect 5742 16594 5794 16606
rect 10446 16658 10498 16670
rect 10446 16594 10498 16606
rect 1344 16490 24640 16524
rect 1344 16438 4126 16490
rect 4178 16438 4230 16490
rect 4282 16438 4334 16490
rect 4386 16438 9950 16490
rect 10002 16438 10054 16490
rect 10106 16438 10158 16490
rect 10210 16438 15774 16490
rect 15826 16438 15878 16490
rect 15930 16438 15982 16490
rect 16034 16438 21598 16490
rect 21650 16438 21702 16490
rect 21754 16438 21806 16490
rect 21858 16438 24640 16490
rect 1344 16404 24640 16438
rect 6078 16322 6130 16334
rect 2482 16270 2494 16322
rect 2546 16270 2558 16322
rect 6078 16258 6130 16270
rect 6302 16322 6354 16334
rect 6302 16258 6354 16270
rect 13582 16322 13634 16334
rect 21858 16270 21870 16322
rect 21922 16270 21934 16322
rect 13582 16258 13634 16270
rect 4958 16210 5010 16222
rect 4162 16158 4174 16210
rect 4226 16158 4238 16210
rect 4958 16146 5010 16158
rect 5070 16210 5122 16222
rect 20638 16210 20690 16222
rect 9538 16158 9550 16210
rect 9602 16158 9614 16210
rect 20178 16158 20190 16210
rect 20242 16158 20254 16210
rect 5070 16146 5122 16158
rect 20638 16146 20690 16158
rect 21310 16210 21362 16222
rect 21310 16146 21362 16158
rect 2718 16098 2770 16110
rect 2482 16046 2494 16098
rect 2546 16046 2558 16098
rect 2718 16034 2770 16046
rect 3390 16098 3442 16110
rect 6526 16098 6578 16110
rect 15038 16098 15090 16110
rect 16494 16098 16546 16110
rect 21534 16098 21586 16110
rect 4050 16046 4062 16098
rect 4114 16046 4126 16098
rect 5842 16046 5854 16098
rect 5906 16046 5918 16098
rect 8754 16046 8766 16098
rect 8818 16046 8830 16098
rect 14578 16046 14590 16098
rect 14642 16046 14654 16098
rect 15810 16046 15822 16098
rect 15874 16046 15886 16098
rect 17266 16046 17278 16098
rect 17330 16046 17342 16098
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 23538 16046 23550 16098
rect 23602 16046 23614 16098
rect 3390 16034 3442 16046
rect 6526 16034 6578 16046
rect 15038 16034 15090 16046
rect 16494 16034 16546 16046
rect 21534 16034 21586 16046
rect 3054 15986 3106 15998
rect 3054 15922 3106 15934
rect 3726 15986 3778 15998
rect 3726 15922 3778 15934
rect 13582 15986 13634 15998
rect 13582 15922 13634 15934
rect 13694 15986 13746 15998
rect 13694 15922 13746 15934
rect 14142 15986 14194 15998
rect 14142 15922 14194 15934
rect 15486 15986 15538 15998
rect 15486 15922 15538 15934
rect 15598 15986 15650 15998
rect 18050 15934 18062 15986
rect 18114 15934 18126 15986
rect 22530 15934 22542 15986
rect 22594 15934 22606 15986
rect 24098 15934 24110 15986
rect 24162 15934 24174 15986
rect 15598 15922 15650 15934
rect 3614 15874 3666 15886
rect 2594 15822 2606 15874
rect 2658 15822 2670 15874
rect 3614 15810 3666 15822
rect 6414 15874 6466 15886
rect 16146 15822 16158 15874
rect 16210 15822 16222 15874
rect 23202 15822 23214 15874
rect 23266 15822 23278 15874
rect 6414 15810 6466 15822
rect 1344 15706 24800 15740
rect 1344 15654 7038 15706
rect 7090 15654 7142 15706
rect 7194 15654 7246 15706
rect 7298 15654 12862 15706
rect 12914 15654 12966 15706
rect 13018 15654 13070 15706
rect 13122 15654 18686 15706
rect 18738 15654 18790 15706
rect 18842 15654 18894 15706
rect 18946 15654 24510 15706
rect 24562 15654 24614 15706
rect 24666 15654 24718 15706
rect 24770 15654 24800 15706
rect 1344 15620 24800 15654
rect 6862 15538 6914 15550
rect 6862 15474 6914 15486
rect 14254 15538 14306 15550
rect 14254 15474 14306 15486
rect 15598 15538 15650 15550
rect 15598 15474 15650 15486
rect 16270 15538 16322 15550
rect 16270 15474 16322 15486
rect 21982 15538 22034 15550
rect 23986 15486 23998 15538
rect 24050 15486 24062 15538
rect 21982 15474 22034 15486
rect 8430 15426 8482 15438
rect 3266 15374 3278 15426
rect 3330 15374 3342 15426
rect 3826 15374 3838 15426
rect 3890 15374 3902 15426
rect 5394 15374 5406 15426
rect 5458 15374 5470 15426
rect 8082 15374 8094 15426
rect 8146 15374 8158 15426
rect 8430 15362 8482 15374
rect 15038 15426 15090 15438
rect 15038 15362 15090 15374
rect 15486 15426 15538 15438
rect 15486 15362 15538 15374
rect 17390 15426 17442 15438
rect 17390 15362 17442 15374
rect 20078 15426 20130 15438
rect 20078 15362 20130 15374
rect 21758 15426 21810 15438
rect 22642 15374 22654 15426
rect 22706 15374 22718 15426
rect 24098 15374 24110 15426
rect 24162 15374 24174 15426
rect 21758 15362 21810 15374
rect 2494 15314 2546 15326
rect 6302 15314 6354 15326
rect 14590 15314 14642 15326
rect 3154 15262 3166 15314
rect 3218 15262 3230 15314
rect 4386 15262 4398 15314
rect 4450 15262 4462 15314
rect 4722 15262 4734 15314
rect 4786 15262 4798 15314
rect 6626 15262 6638 15314
rect 6690 15262 6702 15314
rect 7634 15262 7646 15314
rect 7698 15262 7710 15314
rect 9538 15262 9550 15314
rect 9602 15262 9614 15314
rect 14354 15262 14366 15314
rect 14418 15262 14430 15314
rect 2494 15250 2546 15262
rect 6302 15250 6354 15262
rect 14590 15250 14642 15262
rect 14702 15314 14754 15326
rect 14702 15250 14754 15262
rect 15710 15314 15762 15326
rect 20190 15314 20242 15326
rect 16482 15262 16494 15314
rect 16546 15262 16558 15314
rect 17602 15262 17614 15314
rect 17666 15262 17678 15314
rect 15710 15250 15762 15262
rect 20190 15250 20242 15262
rect 20414 15314 20466 15326
rect 20414 15250 20466 15262
rect 20526 15314 20578 15326
rect 20526 15250 20578 15262
rect 22318 15314 22370 15326
rect 22530 15262 22542 15314
rect 22594 15262 22606 15314
rect 23538 15262 23550 15314
rect 23602 15262 23614 15314
rect 22318 15250 22370 15262
rect 7198 15202 7250 15214
rect 4834 15150 4846 15202
rect 4898 15150 4910 15202
rect 6738 15150 6750 15202
rect 6802 15150 6814 15202
rect 10322 15150 10334 15202
rect 10386 15150 10398 15202
rect 12450 15150 12462 15202
rect 12514 15150 12526 15202
rect 7198 15138 7250 15150
rect 2158 15090 2210 15102
rect 2158 15026 2210 15038
rect 21646 15090 21698 15102
rect 21646 15026 21698 15038
rect 1344 14922 24640 14956
rect 1344 14870 4126 14922
rect 4178 14870 4230 14922
rect 4282 14870 4334 14922
rect 4386 14870 9950 14922
rect 10002 14870 10054 14922
rect 10106 14870 10158 14922
rect 10210 14870 15774 14922
rect 15826 14870 15878 14922
rect 15930 14870 15982 14922
rect 16034 14870 21598 14922
rect 21650 14870 21702 14922
rect 21754 14870 21806 14922
rect 21858 14870 24640 14922
rect 1344 14836 24640 14870
rect 2046 14754 2098 14766
rect 2046 14690 2098 14702
rect 14590 14754 14642 14766
rect 14590 14690 14642 14702
rect 15598 14754 15650 14766
rect 15598 14690 15650 14702
rect 12910 14642 12962 14654
rect 10546 14590 10558 14642
rect 10610 14590 10622 14642
rect 12910 14578 12962 14590
rect 15374 14642 15426 14654
rect 22766 14642 22818 14654
rect 20402 14590 20414 14642
rect 20466 14590 20478 14642
rect 21970 14590 21982 14642
rect 22034 14590 22046 14642
rect 15374 14578 15426 14590
rect 22766 14578 22818 14590
rect 23662 14642 23714 14654
rect 23662 14578 23714 14590
rect 1934 14530 1986 14542
rect 3166 14530 3218 14542
rect 2818 14478 2830 14530
rect 2882 14478 2894 14530
rect 1934 14466 1986 14478
rect 3166 14466 3218 14478
rect 4174 14530 4226 14542
rect 4174 14466 4226 14478
rect 4622 14530 4674 14542
rect 4622 14466 4674 14478
rect 4846 14530 4898 14542
rect 7086 14530 7138 14542
rect 16606 14530 16658 14542
rect 24222 14530 24274 14542
rect 6738 14478 6750 14530
rect 6802 14478 6814 14530
rect 7746 14478 7758 14530
rect 7810 14478 7822 14530
rect 8418 14478 8430 14530
rect 8482 14478 8494 14530
rect 16370 14478 16382 14530
rect 16434 14478 16446 14530
rect 17490 14478 17502 14530
rect 17554 14478 17566 14530
rect 22306 14478 22318 14530
rect 22370 14478 22382 14530
rect 4846 14466 4898 14478
rect 7086 14466 7138 14478
rect 16606 14466 16658 14478
rect 24222 14466 24274 14478
rect 1822 14418 1874 14430
rect 1822 14354 1874 14366
rect 7198 14418 7250 14430
rect 7198 14354 7250 14366
rect 14478 14418 14530 14430
rect 14478 14354 14530 14366
rect 16718 14418 16770 14430
rect 23886 14418 23938 14430
rect 18274 14366 18286 14418
rect 18338 14366 18350 14418
rect 16718 14354 16770 14366
rect 23886 14354 23938 14366
rect 2494 14306 2546 14318
rect 2494 14242 2546 14254
rect 2606 14306 2658 14318
rect 2606 14242 2658 14254
rect 2718 14306 2770 14318
rect 2718 14242 2770 14254
rect 4398 14306 4450 14318
rect 4398 14242 4450 14254
rect 12350 14306 12402 14318
rect 21422 14306 21474 14318
rect 15922 14254 15934 14306
rect 15986 14254 15998 14306
rect 17154 14254 17166 14306
rect 17218 14254 17230 14306
rect 12350 14242 12402 14254
rect 21422 14242 21474 14254
rect 1344 14138 24800 14172
rect 1344 14086 7038 14138
rect 7090 14086 7142 14138
rect 7194 14086 7246 14138
rect 7298 14086 12862 14138
rect 12914 14086 12966 14138
rect 13018 14086 13070 14138
rect 13122 14086 18686 14138
rect 18738 14086 18790 14138
rect 18842 14086 18894 14138
rect 18946 14086 24510 14138
rect 24562 14086 24614 14138
rect 24666 14086 24718 14138
rect 24770 14086 24800 14138
rect 1344 14052 24800 14086
rect 6078 13970 6130 13982
rect 6078 13906 6130 13918
rect 9886 13970 9938 13982
rect 9886 13906 9938 13918
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 18286 13970 18338 13982
rect 18286 13906 18338 13918
rect 23886 13970 23938 13982
rect 23886 13906 23938 13918
rect 6862 13858 6914 13870
rect 6862 13794 6914 13806
rect 6974 13858 7026 13870
rect 6974 13794 7026 13806
rect 7758 13858 7810 13870
rect 17950 13858 18002 13870
rect 14914 13806 14926 13858
rect 14978 13806 14990 13858
rect 19618 13806 19630 13858
rect 19682 13806 19694 13858
rect 7758 13794 7810 13806
rect 17950 13794 18002 13806
rect 5070 13746 5122 13758
rect 6190 13746 6242 13758
rect 5954 13694 5966 13746
rect 6018 13694 6030 13746
rect 5070 13682 5122 13694
rect 6190 13682 6242 13694
rect 6414 13746 6466 13758
rect 6414 13682 6466 13694
rect 9550 13746 9602 13758
rect 9550 13682 9602 13694
rect 11230 13746 11282 13758
rect 19966 13746 20018 13758
rect 11554 13694 11566 13746
rect 11618 13694 11630 13746
rect 20402 13694 20414 13746
rect 20466 13694 20478 13746
rect 24098 13694 24110 13746
rect 24162 13694 24174 13746
rect 11230 13682 11282 13694
rect 19966 13682 20018 13694
rect 7982 13634 8034 13646
rect 7982 13570 8034 13582
rect 8318 13634 8370 13646
rect 8318 13570 8370 13582
rect 17502 13634 17554 13646
rect 21074 13582 21086 13634
rect 21138 13582 21150 13634
rect 23202 13582 23214 13634
rect 23266 13582 23278 13634
rect 17502 13570 17554 13582
rect 5294 13522 5346 13534
rect 5294 13458 5346 13470
rect 5630 13522 5682 13534
rect 5630 13458 5682 13470
rect 6974 13522 7026 13534
rect 6974 13458 7026 13470
rect 1344 13354 24640 13388
rect 1344 13302 4126 13354
rect 4178 13302 4230 13354
rect 4282 13302 4334 13354
rect 4386 13302 9950 13354
rect 10002 13302 10054 13354
rect 10106 13302 10158 13354
rect 10210 13302 15774 13354
rect 15826 13302 15878 13354
rect 15930 13302 15982 13354
rect 16034 13302 21598 13354
rect 21650 13302 21702 13354
rect 21754 13302 21806 13354
rect 21858 13302 24640 13354
rect 1344 13268 24640 13302
rect 21310 13186 21362 13198
rect 21310 13122 21362 13134
rect 18286 13074 18338 13086
rect 2482 13022 2494 13074
rect 2546 13022 2558 13074
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 8642 13022 8654 13074
rect 8706 13022 8718 13074
rect 10770 13022 10782 13074
rect 10834 13022 10846 13074
rect 14242 13022 14254 13074
rect 14306 13022 14318 13074
rect 18286 13010 18338 13022
rect 20190 13074 20242 13086
rect 20190 13010 20242 13022
rect 23886 13074 23938 13086
rect 23886 13010 23938 13022
rect 6190 12962 6242 12974
rect 19182 12962 19234 12974
rect 22990 12962 23042 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 7074 12910 7086 12962
rect 7138 12910 7150 12962
rect 7858 12910 7870 12962
rect 7922 12910 7934 12962
rect 17154 12910 17166 12962
rect 17218 12910 17230 12962
rect 18946 12910 18958 12962
rect 19010 12910 19022 12962
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 21298 12910 21310 12962
rect 21362 12910 21374 12962
rect 23202 12910 23214 12962
rect 23266 12910 23278 12962
rect 6190 12898 6242 12910
rect 19182 12898 19234 12910
rect 22990 12898 23042 12910
rect 20750 12850 20802 12862
rect 16370 12798 16382 12850
rect 16434 12798 16446 12850
rect 20750 12786 20802 12798
rect 21646 12850 21698 12862
rect 21646 12786 21698 12798
rect 22206 12850 22258 12862
rect 22206 12786 22258 12798
rect 6526 12738 6578 12750
rect 6526 12674 6578 12686
rect 6862 12738 6914 12750
rect 6862 12674 6914 12686
rect 22542 12738 22594 12750
rect 22542 12674 22594 12686
rect 1344 12570 24800 12604
rect 1344 12518 7038 12570
rect 7090 12518 7142 12570
rect 7194 12518 7246 12570
rect 7298 12518 12862 12570
rect 12914 12518 12966 12570
rect 13018 12518 13070 12570
rect 13122 12518 18686 12570
rect 18738 12518 18790 12570
rect 18842 12518 18894 12570
rect 18946 12518 24510 12570
rect 24562 12518 24614 12570
rect 24666 12518 24718 12570
rect 24770 12518 24800 12570
rect 1344 12484 24800 12518
rect 15486 12402 15538 12414
rect 15486 12338 15538 12350
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 19294 12402 19346 12414
rect 19294 12338 19346 12350
rect 22766 12402 22818 12414
rect 22766 12338 22818 12350
rect 20862 12290 20914 12302
rect 6626 12238 6638 12290
rect 6690 12238 6702 12290
rect 10322 12238 10334 12290
rect 10386 12238 10398 12290
rect 10658 12238 10670 12290
rect 10722 12238 10734 12290
rect 12450 12238 12462 12290
rect 12514 12238 12526 12290
rect 16370 12238 16382 12290
rect 16434 12238 16446 12290
rect 19730 12238 19742 12290
rect 19794 12238 19806 12290
rect 20862 12226 20914 12238
rect 22206 12290 22258 12302
rect 22206 12226 22258 12238
rect 23102 12290 23154 12302
rect 23102 12226 23154 12238
rect 10894 12178 10946 12190
rect 15262 12178 15314 12190
rect 2034 12126 2046 12178
rect 2098 12126 2110 12178
rect 5954 12126 5966 12178
rect 6018 12126 6030 12178
rect 11666 12126 11678 12178
rect 11730 12126 11742 12178
rect 15026 12126 15038 12178
rect 15090 12126 15102 12178
rect 10894 12114 10946 12126
rect 15262 12114 15314 12126
rect 15598 12178 15650 12190
rect 19182 12178 19234 12190
rect 16146 12126 16158 12178
rect 16210 12126 16222 12178
rect 15598 12114 15650 12126
rect 19182 12114 19234 12126
rect 20078 12178 20130 12190
rect 20078 12114 20130 12126
rect 20302 12178 20354 12190
rect 23998 12178 24050 12190
rect 20626 12126 20638 12178
rect 20690 12126 20702 12178
rect 21746 12126 21758 12178
rect 21810 12126 21822 12178
rect 23538 12126 23550 12178
rect 23602 12126 23614 12178
rect 20302 12114 20354 12126
rect 23998 12114 24050 12126
rect 15374 12066 15426 12078
rect 2706 12014 2718 12066
rect 2770 12014 2782 12066
rect 4834 12014 4846 12066
rect 4898 12014 4910 12066
rect 8754 12014 8766 12066
rect 8818 12014 8830 12066
rect 14578 12014 14590 12066
rect 14642 12014 14654 12066
rect 15374 12002 15426 12014
rect 16830 12066 16882 12078
rect 16830 12002 16882 12014
rect 20974 12066 21026 12078
rect 21298 12014 21310 12066
rect 21362 12014 21374 12066
rect 20974 12002 21026 12014
rect 11230 11954 11282 11966
rect 11230 11890 11282 11902
rect 19294 11954 19346 11966
rect 19294 11890 19346 11902
rect 1344 11786 24640 11820
rect 1344 11734 4126 11786
rect 4178 11734 4230 11786
rect 4282 11734 4334 11786
rect 4386 11734 9950 11786
rect 10002 11734 10054 11786
rect 10106 11734 10158 11786
rect 10210 11734 15774 11786
rect 15826 11734 15878 11786
rect 15930 11734 15982 11786
rect 16034 11734 21598 11786
rect 21650 11734 21702 11786
rect 21754 11734 21806 11786
rect 21858 11734 24640 11786
rect 1344 11700 24640 11734
rect 13918 11618 13970 11630
rect 13918 11554 13970 11566
rect 21198 11618 21250 11630
rect 21198 11554 21250 11566
rect 3166 11506 3218 11518
rect 23762 11454 23774 11506
rect 23826 11454 23838 11506
rect 3166 11442 3218 11454
rect 21422 11394 21474 11406
rect 3378 11342 3390 11394
rect 3442 11342 3454 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 14690 11342 14702 11394
rect 14754 11342 14766 11394
rect 15474 11342 15486 11394
rect 15538 11342 15550 11394
rect 21422 11330 21474 11342
rect 21870 11394 21922 11406
rect 21870 11330 21922 11342
rect 22094 11394 22146 11406
rect 23090 11342 23102 11394
rect 23154 11342 23166 11394
rect 23538 11342 23550 11394
rect 23602 11342 23614 11394
rect 22094 11330 22146 11342
rect 3054 11282 3106 11294
rect 12686 11282 12738 11294
rect 9314 11230 9326 11282
rect 9378 11230 9390 11282
rect 3054 11218 3106 11230
rect 12686 11218 12738 11230
rect 13582 11282 13634 11294
rect 21982 11282 22034 11294
rect 14466 11230 14478 11282
rect 14530 11230 14542 11282
rect 17490 11230 17502 11282
rect 17554 11230 17566 11282
rect 22530 11230 22542 11282
rect 22594 11230 22606 11282
rect 24098 11230 24110 11282
rect 24162 11230 24174 11282
rect 13582 11218 13634 11230
rect 21982 11218 22034 11230
rect 12350 11170 12402 11182
rect 12350 11106 12402 11118
rect 1344 11002 24800 11036
rect 1344 10950 7038 11002
rect 7090 10950 7142 11002
rect 7194 10950 7246 11002
rect 7298 10950 12862 11002
rect 12914 10950 12966 11002
rect 13018 10950 13070 11002
rect 13122 10950 18686 11002
rect 18738 10950 18790 11002
rect 18842 10950 18894 11002
rect 18946 10950 24510 11002
rect 24562 10950 24614 11002
rect 24666 10950 24718 11002
rect 24770 10950 24800 11002
rect 1344 10916 24800 10950
rect 3166 10834 3218 10846
rect 3166 10770 3218 10782
rect 14926 10834 14978 10846
rect 14926 10770 14978 10782
rect 15934 10834 15986 10846
rect 15934 10770 15986 10782
rect 16494 10834 16546 10846
rect 16494 10770 16546 10782
rect 24222 10834 24274 10846
rect 24222 10770 24274 10782
rect 2494 10722 2546 10734
rect 22654 10722 22706 10734
rect 4274 10670 4286 10722
rect 4338 10670 4350 10722
rect 5506 10670 5518 10722
rect 5570 10670 5582 10722
rect 9762 10670 9774 10722
rect 9826 10670 9838 10722
rect 10210 10670 10222 10722
rect 10274 10670 10286 10722
rect 12114 10670 12126 10722
rect 12178 10670 12190 10722
rect 2494 10658 2546 10670
rect 22654 10658 22706 10670
rect 3502 10610 3554 10622
rect 10446 10610 10498 10622
rect 16382 10610 16434 10622
rect 21422 10610 21474 10622
rect 2258 10558 2270 10610
rect 2322 10558 2334 10610
rect 3938 10558 3950 10610
rect 4002 10558 4014 10610
rect 4834 10558 4846 10610
rect 4898 10558 4910 10610
rect 11330 10558 11342 10610
rect 11394 10558 11406 10610
rect 17378 10558 17390 10610
rect 17442 10558 17454 10610
rect 3502 10546 3554 10558
rect 10446 10546 10498 10558
rect 16382 10546 16434 10558
rect 21422 10546 21474 10558
rect 21646 10610 21698 10622
rect 21646 10546 21698 10558
rect 21982 10610 22034 10622
rect 23202 10558 23214 10610
rect 23266 10558 23278 10610
rect 21982 10546 22034 10558
rect 21534 10498 21586 10510
rect 7634 10446 7646 10498
rect 7698 10446 7710 10498
rect 14242 10446 14254 10498
rect 14306 10446 14318 10498
rect 15474 10446 15486 10498
rect 15538 10446 15550 10498
rect 18162 10446 18174 10498
rect 18226 10446 18238 10498
rect 20290 10446 20302 10498
rect 20354 10446 20366 10498
rect 23426 10446 23438 10498
rect 23490 10446 23502 10498
rect 21534 10434 21586 10446
rect 10782 10386 10834 10398
rect 10782 10322 10834 10334
rect 16270 10386 16322 10398
rect 16270 10322 16322 10334
rect 1344 10218 24640 10252
rect 1344 10166 4126 10218
rect 4178 10166 4230 10218
rect 4282 10166 4334 10218
rect 4386 10166 9950 10218
rect 10002 10166 10054 10218
rect 10106 10166 10158 10218
rect 10210 10166 15774 10218
rect 15826 10166 15878 10218
rect 15930 10166 15982 10218
rect 16034 10166 21598 10218
rect 21650 10166 21702 10218
rect 21754 10166 21806 10218
rect 21858 10166 24640 10218
rect 1344 10132 24640 10166
rect 18174 10050 18226 10062
rect 18174 9986 18226 9998
rect 20302 9938 20354 9950
rect 2482 9886 2494 9938
rect 2546 9886 2558 9938
rect 4610 9886 4622 9938
rect 4674 9886 4686 9938
rect 12002 9886 12014 9938
rect 12066 9886 12078 9938
rect 19170 9886 19182 9938
rect 19234 9886 19246 9938
rect 24210 9886 24222 9938
rect 24274 9886 24286 9938
rect 20302 9874 20354 9886
rect 15038 9826 15090 9838
rect 1810 9774 1822 9826
rect 1874 9774 1886 9826
rect 8530 9774 8542 9826
rect 8594 9774 8606 9826
rect 9202 9774 9214 9826
rect 9266 9774 9278 9826
rect 15038 9762 15090 9774
rect 15262 9826 15314 9838
rect 20526 9826 20578 9838
rect 19506 9774 19518 9826
rect 19570 9774 19582 9826
rect 20738 9774 20750 9826
rect 20802 9774 20814 9826
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 15262 9762 15314 9774
rect 20526 9762 20578 9774
rect 14814 9714 14866 9726
rect 9874 9662 9886 9714
rect 9938 9662 9950 9714
rect 14814 9650 14866 9662
rect 18286 9714 18338 9726
rect 18286 9650 18338 9662
rect 18510 9714 18562 9726
rect 18510 9650 18562 9662
rect 18846 9714 18898 9726
rect 18846 9650 18898 9662
rect 20190 9714 20242 9726
rect 22082 9662 22094 9714
rect 22146 9662 22158 9714
rect 20190 9650 20242 9662
rect 8766 9602 8818 9614
rect 8766 9538 8818 9550
rect 14926 9602 14978 9614
rect 14926 9538 14978 9550
rect 1344 9434 24800 9468
rect 1344 9382 7038 9434
rect 7090 9382 7142 9434
rect 7194 9382 7246 9434
rect 7298 9382 12862 9434
rect 12914 9382 12966 9434
rect 13018 9382 13070 9434
rect 13122 9382 18686 9434
rect 18738 9382 18790 9434
rect 18842 9382 18894 9434
rect 18946 9382 24510 9434
rect 24562 9382 24614 9434
rect 24666 9382 24718 9434
rect 24770 9382 24800 9434
rect 1344 9348 24800 9382
rect 4510 9266 4562 9278
rect 4510 9202 4562 9214
rect 7310 9266 7362 9278
rect 7310 9202 7362 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 16046 9266 16098 9278
rect 16046 9202 16098 9214
rect 16382 9266 16434 9278
rect 16382 9202 16434 9214
rect 20974 9266 21026 9278
rect 20974 9202 21026 9214
rect 21198 9266 21250 9278
rect 21198 9202 21250 9214
rect 22766 9266 22818 9278
rect 22766 9202 22818 9214
rect 21870 9154 21922 9166
rect 3826 9102 3838 9154
rect 3890 9102 3902 9154
rect 5394 9102 5406 9154
rect 5458 9102 5470 9154
rect 10322 9102 10334 9154
rect 10386 9102 10398 9154
rect 10770 9102 10782 9154
rect 10834 9102 10846 9154
rect 14690 9102 14702 9154
rect 14754 9102 14766 9154
rect 18162 9102 18174 9154
rect 18226 9102 18238 9154
rect 21870 9090 21922 9102
rect 24110 9154 24162 9166
rect 24110 9090 24162 9102
rect 4846 9042 4898 9054
rect 9998 9042 10050 9054
rect 3938 8990 3950 9042
rect 4002 8990 4014 9042
rect 5618 8990 5630 9042
rect 5682 8990 5694 9042
rect 7074 8990 7086 9042
rect 7138 8990 7150 9042
rect 4846 8978 4898 8990
rect 9998 8978 10050 8990
rect 11902 9042 11954 9054
rect 16270 9042 16322 9054
rect 21982 9042 22034 9054
rect 15474 8990 15486 9042
rect 15538 8990 15550 9042
rect 15810 8990 15822 9042
rect 15874 8990 15886 9042
rect 17378 8990 17390 9042
rect 17442 8990 17454 9042
rect 20738 8990 20750 9042
rect 20802 8990 20814 9042
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 23426 8990 23438 9042
rect 23490 8990 23502 9042
rect 23874 8990 23886 9042
rect 23938 8990 23950 9042
rect 11902 8978 11954 8990
rect 16270 8978 16322 8990
rect 21982 8978 22034 8990
rect 11342 8930 11394 8942
rect 16158 8930 16210 8942
rect 22206 8930 22258 8942
rect 12562 8878 12574 8930
rect 12626 8878 12638 8930
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 11342 8866 11394 8878
rect 16158 8866 16210 8878
rect 22206 8866 22258 8878
rect 2830 8818 2882 8830
rect 2830 8754 2882 8766
rect 3166 8818 3218 8830
rect 3166 8754 3218 8766
rect 1344 8650 24640 8684
rect 1344 8598 4126 8650
rect 4178 8598 4230 8650
rect 4282 8598 4334 8650
rect 4386 8598 9950 8650
rect 10002 8598 10054 8650
rect 10106 8598 10158 8650
rect 10210 8598 15774 8650
rect 15826 8598 15878 8650
rect 15930 8598 15982 8650
rect 16034 8598 21598 8650
rect 21650 8598 21702 8650
rect 21754 8598 21806 8650
rect 21858 8598 24640 8650
rect 1344 8564 24640 8598
rect 21646 8482 21698 8494
rect 20290 8430 20302 8482
rect 20354 8430 20366 8482
rect 21646 8418 21698 8430
rect 22094 8482 22146 8494
rect 22094 8418 22146 8430
rect 11790 8370 11842 8382
rect 4610 8318 4622 8370
rect 4674 8318 4686 8370
rect 7522 8318 7534 8370
rect 7586 8318 7598 8370
rect 9650 8318 9662 8370
rect 9714 8318 9726 8370
rect 10098 8318 10110 8370
rect 10162 8318 10174 8370
rect 11790 8306 11842 8318
rect 15262 8370 15314 8382
rect 15262 8306 15314 8318
rect 15374 8370 15426 8382
rect 15374 8306 15426 8318
rect 15710 8370 15762 8382
rect 15710 8306 15762 8318
rect 23102 8370 23154 8382
rect 23538 8318 23550 8370
rect 23602 8318 23614 8370
rect 23102 8306 23154 8318
rect 19630 8258 19682 8270
rect 1810 8206 1822 8258
rect 1874 8206 1886 8258
rect 6850 8206 6862 8258
rect 6914 8206 6926 8258
rect 10434 8206 10446 8258
rect 10498 8206 10510 8258
rect 19630 8194 19682 8206
rect 19854 8258 19906 8270
rect 19854 8194 19906 8206
rect 21758 8258 21810 8270
rect 21758 8194 21810 8206
rect 21982 8258 22034 8270
rect 22530 8206 22542 8258
rect 22594 8206 22606 8258
rect 23762 8206 23774 8258
rect 23826 8206 23838 8258
rect 21982 8194 22034 8206
rect 19742 8146 19794 8158
rect 2482 8094 2494 8146
rect 2546 8094 2558 8146
rect 10994 8094 11006 8146
rect 11058 8094 11070 8146
rect 11554 8094 11566 8146
rect 11618 8094 11630 8146
rect 19742 8082 19794 8094
rect 22766 8146 22818 8158
rect 22766 8082 22818 8094
rect 12126 8034 12178 8046
rect 12126 7970 12178 7982
rect 15822 8034 15874 8046
rect 15822 7970 15874 7982
rect 1344 7866 24800 7900
rect 1344 7814 7038 7866
rect 7090 7814 7142 7866
rect 7194 7814 7246 7866
rect 7298 7814 12862 7866
rect 12914 7814 12966 7866
rect 13018 7814 13070 7866
rect 13122 7814 18686 7866
rect 18738 7814 18790 7866
rect 18842 7814 18894 7866
rect 18946 7814 24510 7866
rect 24562 7814 24614 7866
rect 24666 7814 24718 7866
rect 24770 7814 24800 7866
rect 1344 7780 24800 7814
rect 2494 7698 2546 7710
rect 2494 7634 2546 7646
rect 3838 7698 3890 7710
rect 21534 7698 21586 7710
rect 19730 7646 19742 7698
rect 19794 7646 19806 7698
rect 3838 7634 3890 7646
rect 21534 7634 21586 7646
rect 22654 7698 22706 7710
rect 22654 7634 22706 7646
rect 7198 7586 7250 7598
rect 21310 7586 21362 7598
rect 4946 7534 4958 7586
rect 5010 7534 5022 7586
rect 6626 7534 6638 7586
rect 6690 7534 6702 7586
rect 7746 7534 7758 7586
rect 7810 7534 7822 7586
rect 8306 7534 8318 7586
rect 8370 7534 8382 7586
rect 10546 7534 10558 7586
rect 10610 7534 10622 7586
rect 11106 7534 11118 7586
rect 11170 7534 11182 7586
rect 12562 7534 12574 7586
rect 12626 7534 12638 7586
rect 16034 7534 16046 7586
rect 16098 7534 16110 7586
rect 7198 7522 7250 7534
rect 21310 7522 21362 7534
rect 22878 7586 22930 7598
rect 22878 7522 22930 7534
rect 4174 7474 4226 7486
rect 7534 7474 7586 7486
rect 2258 7422 2270 7474
rect 2322 7422 2334 7474
rect 4834 7422 4846 7474
rect 4898 7422 4910 7474
rect 6402 7422 6414 7474
rect 6466 7422 6478 7474
rect 4174 7410 4226 7422
rect 7534 7410 7586 7422
rect 10334 7474 10386 7486
rect 10334 7410 10386 7422
rect 12014 7474 12066 7486
rect 20078 7474 20130 7486
rect 12786 7422 12798 7474
rect 12850 7422 12862 7474
rect 16818 7422 16830 7474
rect 16882 7422 16894 7474
rect 23314 7422 23326 7474
rect 23378 7422 23390 7474
rect 12014 7410 12066 7422
rect 20078 7410 20130 7422
rect 13906 7310 13918 7362
rect 13970 7310 13982 7362
rect 21634 7310 21646 7362
rect 21698 7310 21710 7362
rect 23650 7310 23662 7362
rect 23714 7310 23726 7362
rect 5518 7250 5570 7262
rect 5518 7186 5570 7198
rect 5854 7250 5906 7262
rect 5854 7186 5906 7198
rect 9998 7250 10050 7262
rect 9998 7186 10050 7198
rect 11678 7250 11730 7262
rect 11678 7186 11730 7198
rect 1344 7082 24640 7116
rect 1344 7030 4126 7082
rect 4178 7030 4230 7082
rect 4282 7030 4334 7082
rect 4386 7030 9950 7082
rect 10002 7030 10054 7082
rect 10106 7030 10158 7082
rect 10210 7030 15774 7082
rect 15826 7030 15878 7082
rect 15930 7030 15982 7082
rect 16034 7030 21598 7082
rect 21650 7030 21702 7082
rect 21754 7030 21806 7082
rect 21858 7030 24640 7082
rect 1344 6996 24640 7030
rect 9214 6914 9266 6926
rect 9214 6850 9266 6862
rect 19954 6750 19966 6802
rect 20018 6750 20030 6802
rect 20738 6750 20750 6802
rect 20802 6750 20814 6802
rect 24210 6750 24222 6802
rect 24274 6750 24286 6802
rect 4734 6690 4786 6702
rect 4734 6626 4786 6638
rect 8318 6690 8370 6702
rect 8318 6626 8370 6638
rect 8878 6690 8930 6702
rect 11790 6690 11842 6702
rect 9986 6638 9998 6690
rect 10050 6638 10062 6690
rect 17042 6638 17054 6690
rect 17106 6638 17118 6690
rect 21410 6638 21422 6690
rect 21474 6638 21486 6690
rect 8878 6626 8930 6638
rect 11790 6626 11842 6638
rect 20414 6578 20466 6590
rect 9762 6526 9774 6578
rect 9826 6526 9838 6578
rect 17826 6526 17838 6578
rect 17890 6526 17902 6578
rect 20414 6514 20466 6526
rect 20638 6578 20690 6590
rect 22082 6526 22094 6578
rect 22146 6526 22158 6578
rect 20638 6514 20690 6526
rect 4398 6466 4450 6478
rect 4398 6402 4450 6414
rect 7982 6466 8034 6478
rect 7982 6402 8034 6414
rect 12126 6466 12178 6478
rect 12126 6402 12178 6414
rect 1344 6298 24800 6332
rect 1344 6246 7038 6298
rect 7090 6246 7142 6298
rect 7194 6246 7246 6298
rect 7298 6246 12862 6298
rect 12914 6246 12966 6298
rect 13018 6246 13070 6298
rect 13122 6246 18686 6298
rect 18738 6246 18790 6298
rect 18842 6246 18894 6298
rect 18946 6246 24510 6298
rect 24562 6246 24614 6298
rect 24666 6246 24718 6298
rect 24770 6246 24800 6298
rect 1344 6212 24800 6246
rect 18510 6130 18562 6142
rect 18510 6066 18562 6078
rect 22766 6130 22818 6142
rect 22766 6066 22818 6078
rect 18398 6018 18450 6030
rect 24110 6018 24162 6030
rect 4050 5966 4062 6018
rect 4114 5966 4126 6018
rect 13458 5966 13470 6018
rect 13522 5966 13534 6018
rect 22418 5966 22430 6018
rect 22482 5966 22494 6018
rect 18398 5954 18450 5966
rect 24110 5954 24162 5966
rect 20414 5906 20466 5918
rect 3378 5854 3390 5906
rect 3442 5854 3454 5906
rect 14242 5854 14254 5906
rect 14306 5854 14318 5906
rect 18722 5854 18734 5906
rect 18786 5854 18798 5906
rect 19730 5854 19742 5906
rect 19794 5854 19806 5906
rect 20414 5842 20466 5854
rect 23214 5906 23266 5918
rect 23650 5854 23662 5906
rect 23714 5854 23726 5906
rect 23214 5842 23266 5854
rect 20526 5794 20578 5806
rect 6178 5742 6190 5794
rect 6242 5742 6254 5794
rect 11330 5742 11342 5794
rect 11394 5742 11406 5794
rect 20526 5730 20578 5742
rect 1344 5514 24640 5548
rect 1344 5462 4126 5514
rect 4178 5462 4230 5514
rect 4282 5462 4334 5514
rect 4386 5462 9950 5514
rect 10002 5462 10054 5514
rect 10106 5462 10158 5514
rect 10210 5462 15774 5514
rect 15826 5462 15878 5514
rect 15930 5462 15982 5514
rect 16034 5462 21598 5514
rect 21650 5462 21702 5514
rect 21754 5462 21806 5514
rect 21858 5462 24640 5514
rect 1344 5428 24640 5462
rect 23662 5234 23714 5246
rect 7746 5182 7758 5234
rect 7810 5182 7822 5234
rect 9874 5182 9886 5234
rect 9938 5182 9950 5234
rect 23662 5170 23714 5182
rect 24222 5122 24274 5134
rect 6962 5070 6974 5122
rect 7026 5070 7038 5122
rect 24222 5058 24274 5070
rect 23886 5010 23938 5022
rect 23886 4946 23938 4958
rect 1344 4730 24800 4764
rect 1344 4678 7038 4730
rect 7090 4678 7142 4730
rect 7194 4678 7246 4730
rect 7298 4678 12862 4730
rect 12914 4678 12966 4730
rect 13018 4678 13070 4730
rect 13122 4678 18686 4730
rect 18738 4678 18790 4730
rect 18842 4678 18894 4730
rect 18946 4678 24510 4730
rect 24562 4678 24614 4730
rect 24666 4678 24718 4730
rect 24770 4678 24800 4730
rect 1344 4644 24800 4678
rect 23886 4562 23938 4574
rect 23886 4498 23938 4510
rect 24222 4338 24274 4350
rect 24222 4274 24274 4286
rect 23662 4226 23714 4238
rect 23662 4162 23714 4174
rect 1344 3946 24640 3980
rect 1344 3894 4126 3946
rect 4178 3894 4230 3946
rect 4282 3894 4334 3946
rect 4386 3894 9950 3946
rect 10002 3894 10054 3946
rect 10106 3894 10158 3946
rect 10210 3894 15774 3946
rect 15826 3894 15878 3946
rect 15930 3894 15982 3946
rect 16034 3894 21598 3946
rect 21650 3894 21702 3946
rect 21754 3894 21806 3946
rect 21858 3894 24640 3946
rect 1344 3860 24640 3894
rect 23438 3442 23490 3454
rect 23438 3378 23490 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 1344 3162 24800 3196
rect 1344 3110 7038 3162
rect 7090 3110 7142 3162
rect 7194 3110 7246 3162
rect 7298 3110 12862 3162
rect 12914 3110 12966 3162
rect 13018 3110 13070 3162
rect 13122 3110 18686 3162
rect 18738 3110 18790 3162
rect 18842 3110 18894 3162
rect 18946 3110 24510 3162
rect 24562 3110 24614 3162
rect 24666 3110 24718 3162
rect 24770 3110 24800 3162
rect 1344 3076 24800 3110
<< via1 >>
rect 4126 22710 4178 22762
rect 4230 22710 4282 22762
rect 4334 22710 4386 22762
rect 9950 22710 10002 22762
rect 10054 22710 10106 22762
rect 10158 22710 10210 22762
rect 15774 22710 15826 22762
rect 15878 22710 15930 22762
rect 15982 22710 16034 22762
rect 21598 22710 21650 22762
rect 21702 22710 21754 22762
rect 21806 22710 21858 22762
rect 22430 22542 22482 22594
rect 12686 22430 12738 22482
rect 13358 22318 13410 22370
rect 19630 22318 19682 22370
rect 19966 22318 20018 22370
rect 20862 22318 20914 22370
rect 21422 22318 21474 22370
rect 13134 22094 13186 22146
rect 18734 22094 18786 22146
rect 19182 22094 19234 22146
rect 20190 22094 20242 22146
rect 21086 22094 21138 22146
rect 7038 21926 7090 21978
rect 7142 21926 7194 21978
rect 7246 21926 7298 21978
rect 12862 21926 12914 21978
rect 12966 21926 13018 21978
rect 13070 21926 13122 21978
rect 18686 21926 18738 21978
rect 18790 21926 18842 21978
rect 18894 21926 18946 21978
rect 24510 21926 24562 21978
rect 24614 21926 24666 21978
rect 24718 21926 24770 21978
rect 8206 21758 8258 21810
rect 17502 21646 17554 21698
rect 5070 21534 5122 21586
rect 8430 21534 8482 21586
rect 9662 21534 9714 21586
rect 13022 21534 13074 21586
rect 16270 21534 16322 21586
rect 17390 21534 17442 21586
rect 17950 21534 18002 21586
rect 21198 21534 21250 21586
rect 5742 21422 5794 21474
rect 7870 21422 7922 21474
rect 10446 21422 10498 21474
rect 12574 21422 12626 21474
rect 13694 21422 13746 21474
rect 15822 21422 15874 21474
rect 18734 21422 18786 21474
rect 20862 21422 20914 21474
rect 21982 21422 22034 21474
rect 24110 21422 24162 21474
rect 17502 21310 17554 21362
rect 4126 21142 4178 21194
rect 4230 21142 4282 21194
rect 4334 21142 4386 21194
rect 9950 21142 10002 21194
rect 10054 21142 10106 21194
rect 10158 21142 10210 21194
rect 15774 21142 15826 21194
rect 15878 21142 15930 21194
rect 15982 21142 16034 21194
rect 21598 21142 21650 21194
rect 21702 21142 21754 21194
rect 21806 21142 21858 21194
rect 8878 20974 8930 21026
rect 5070 20862 5122 20914
rect 18510 20862 18562 20914
rect 19630 20862 19682 20914
rect 20414 20862 20466 20914
rect 2270 20750 2322 20802
rect 8094 20750 8146 20802
rect 8654 20750 8706 20802
rect 9326 20750 9378 20802
rect 15598 20750 15650 20802
rect 19518 20750 19570 20802
rect 21982 20750 22034 20802
rect 22430 20750 22482 20802
rect 23214 20750 23266 20802
rect 23550 20750 23602 20802
rect 2942 20638 2994 20690
rect 7646 20638 7698 20690
rect 8318 20638 8370 20690
rect 9886 20638 9938 20690
rect 10446 20638 10498 20690
rect 16382 20638 16434 20690
rect 19966 20638 20018 20690
rect 20302 20638 20354 20690
rect 21758 20638 21810 20690
rect 24110 20638 24162 20690
rect 7758 20526 7810 20578
rect 9998 20526 10050 20578
rect 10222 20526 10274 20578
rect 10558 20526 10610 20578
rect 10782 20526 10834 20578
rect 20526 20526 20578 20578
rect 21534 20526 21586 20578
rect 7038 20358 7090 20410
rect 7142 20358 7194 20410
rect 7246 20358 7298 20410
rect 12862 20358 12914 20410
rect 12966 20358 13018 20410
rect 13070 20358 13122 20410
rect 18686 20358 18738 20410
rect 18790 20358 18842 20410
rect 18894 20358 18946 20410
rect 24510 20358 24562 20410
rect 24614 20358 24666 20410
rect 24718 20358 24770 20410
rect 6750 20190 6802 20242
rect 8878 20190 8930 20242
rect 13918 20190 13970 20242
rect 4958 20078 5010 20130
rect 9550 20078 9602 20130
rect 9998 20078 10050 20130
rect 11342 20078 11394 20130
rect 12910 20078 12962 20130
rect 14142 20078 14194 20130
rect 14926 20078 14978 20130
rect 16494 20078 16546 20130
rect 16606 20078 16658 20130
rect 18734 20078 18786 20130
rect 19406 20078 19458 20130
rect 19854 20078 19906 20130
rect 20414 20078 20466 20130
rect 20638 20078 20690 20130
rect 21310 20078 21362 20130
rect 21870 20078 21922 20130
rect 22094 20078 22146 20130
rect 22430 20078 22482 20130
rect 4398 19966 4450 20018
rect 7758 19966 7810 20018
rect 7982 19966 8034 20018
rect 8990 19966 9042 20018
rect 9774 19966 9826 20018
rect 11230 19966 11282 20018
rect 11566 19966 11618 20018
rect 13134 19966 13186 20018
rect 13582 19966 13634 20018
rect 13806 19966 13858 20018
rect 14254 19966 14306 20018
rect 15262 19966 15314 20018
rect 16046 19966 16098 20018
rect 16830 19966 16882 20018
rect 18174 19966 18226 20018
rect 19630 19966 19682 20018
rect 19966 19966 20018 20018
rect 21086 19966 21138 20018
rect 21646 19966 21698 20018
rect 22766 19966 22818 20018
rect 23214 19966 23266 20018
rect 23662 19966 23714 20018
rect 4510 19854 4562 19906
rect 6638 19854 6690 19906
rect 7086 19854 7138 19906
rect 9886 19854 9938 19906
rect 13358 19854 13410 19906
rect 16494 19854 16546 19906
rect 17950 19854 18002 19906
rect 20302 19854 20354 19906
rect 21982 19854 22034 19906
rect 24110 19854 24162 19906
rect 8878 19742 8930 19794
rect 17838 19742 17890 19794
rect 4126 19574 4178 19626
rect 4230 19574 4282 19626
rect 4334 19574 4386 19626
rect 9950 19574 10002 19626
rect 10054 19574 10106 19626
rect 10158 19574 10210 19626
rect 15774 19574 15826 19626
rect 15878 19574 15930 19626
rect 15982 19574 16034 19626
rect 21598 19574 21650 19626
rect 21702 19574 21754 19626
rect 21806 19574 21858 19626
rect 7534 19406 7586 19458
rect 11790 19406 11842 19458
rect 11902 19406 11954 19458
rect 12574 19406 12626 19458
rect 16718 19406 16770 19458
rect 20414 19406 20466 19458
rect 20862 19406 20914 19458
rect 21646 19406 21698 19458
rect 13806 19294 13858 19346
rect 15486 19294 15538 19346
rect 17950 19294 18002 19346
rect 20078 19294 20130 19346
rect 20526 19294 20578 19346
rect 21422 19294 21474 19346
rect 22878 19294 22930 19346
rect 4398 19182 4450 19234
rect 7422 19182 7474 19234
rect 7870 19182 7922 19234
rect 8094 19182 8146 19234
rect 8206 19182 8258 19234
rect 9102 19182 9154 19234
rect 10670 19182 10722 19234
rect 10894 19182 10946 19234
rect 11902 19182 11954 19234
rect 12350 19182 12402 19234
rect 13918 19182 13970 19234
rect 14366 19182 14418 19234
rect 14590 19182 14642 19234
rect 14814 19182 14866 19234
rect 14926 19182 14978 19234
rect 15374 19182 15426 19234
rect 16942 19182 16994 19234
rect 17278 19182 17330 19234
rect 22990 19182 23042 19234
rect 3278 19070 3330 19122
rect 3950 19070 4002 19122
rect 4286 19070 4338 19122
rect 8654 19070 8706 19122
rect 9438 19070 9490 19122
rect 9774 19070 9826 19122
rect 10110 19070 10162 19122
rect 10334 19070 10386 19122
rect 21422 19070 21474 19122
rect 21982 19070 22034 19122
rect 23662 19070 23714 19122
rect 9326 18958 9378 19010
rect 9998 18958 10050 19010
rect 11230 18958 11282 19010
rect 14478 18958 14530 19010
rect 16382 18958 16434 19010
rect 16606 18958 16658 19010
rect 22094 18958 22146 19010
rect 22206 18958 22258 19010
rect 24110 18958 24162 19010
rect 7038 18790 7090 18842
rect 7142 18790 7194 18842
rect 7246 18790 7298 18842
rect 12862 18790 12914 18842
rect 12966 18790 13018 18842
rect 13070 18790 13122 18842
rect 18686 18790 18738 18842
rect 18790 18790 18842 18842
rect 18894 18790 18946 18842
rect 24510 18790 24562 18842
rect 24614 18790 24666 18842
rect 24718 18790 24770 18842
rect 11118 18622 11170 18674
rect 11342 18622 11394 18674
rect 14254 18622 14306 18674
rect 14366 18622 14418 18674
rect 5182 18510 5234 18562
rect 7758 18510 7810 18562
rect 11566 18510 11618 18562
rect 12238 18510 12290 18562
rect 12574 18510 12626 18562
rect 14142 18510 14194 18562
rect 15262 18510 15314 18562
rect 17390 18510 17442 18562
rect 1822 18398 1874 18450
rect 4958 18398 5010 18450
rect 5518 18398 5570 18450
rect 6414 18398 6466 18450
rect 6862 18398 6914 18450
rect 7198 18398 7250 18450
rect 7982 18398 8034 18450
rect 8430 18398 8482 18450
rect 8990 18398 9042 18450
rect 10782 18398 10834 18450
rect 12014 18398 12066 18450
rect 12910 18398 12962 18450
rect 14814 18398 14866 18450
rect 15150 18398 15202 18450
rect 17614 18398 17666 18450
rect 19182 18398 19234 18450
rect 19966 18398 20018 18450
rect 20078 18398 20130 18450
rect 23550 18398 23602 18450
rect 24110 18398 24162 18450
rect 2494 18286 2546 18338
rect 4622 18286 4674 18338
rect 9774 18286 9826 18338
rect 19406 18286 19458 18338
rect 20414 18286 20466 18338
rect 20750 18286 20802 18338
rect 22878 18286 22930 18338
rect 4846 18174 4898 18226
rect 11006 18174 11058 18226
rect 15038 18174 15090 18226
rect 19518 18174 19570 18226
rect 20302 18174 20354 18226
rect 4126 18006 4178 18058
rect 4230 18006 4282 18058
rect 4334 18006 4386 18058
rect 9950 18006 10002 18058
rect 10054 18006 10106 18058
rect 10158 18006 10210 18058
rect 15774 18006 15826 18058
rect 15878 18006 15930 18058
rect 15982 18006 16034 18058
rect 21598 18006 21650 18058
rect 21702 18006 21754 18058
rect 21806 18006 21858 18058
rect 3614 17838 3666 17890
rect 9550 17838 9602 17890
rect 14366 17838 14418 17890
rect 16494 17838 16546 17890
rect 20190 17838 20242 17890
rect 20526 17838 20578 17890
rect 3838 17726 3890 17778
rect 5630 17726 5682 17778
rect 9326 17726 9378 17778
rect 10894 17726 10946 17778
rect 12014 17726 12066 17778
rect 15934 17726 15986 17778
rect 20750 17726 20802 17778
rect 21982 17726 22034 17778
rect 2942 17614 2994 17666
rect 4398 17614 4450 17666
rect 6750 17614 6802 17666
rect 7198 17614 7250 17666
rect 8766 17614 8818 17666
rect 11342 17614 11394 17666
rect 16158 17614 16210 17666
rect 16830 17614 16882 17666
rect 17166 17614 17218 17666
rect 18062 17614 18114 17666
rect 19182 17614 19234 17666
rect 22318 17614 22370 17666
rect 24110 17614 24162 17666
rect 8542 17502 8594 17554
rect 14478 17502 14530 17554
rect 16942 17502 16994 17554
rect 22766 17502 22818 17554
rect 2382 17390 2434 17442
rect 3278 17390 3330 17442
rect 4286 17390 4338 17442
rect 9886 17390 9938 17442
rect 11902 17390 11954 17442
rect 14366 17390 14418 17442
rect 18286 17390 18338 17442
rect 19518 17390 19570 17442
rect 23886 17390 23938 17442
rect 7038 17222 7090 17274
rect 7142 17222 7194 17274
rect 7246 17222 7298 17274
rect 12862 17222 12914 17274
rect 12966 17222 13018 17274
rect 13070 17222 13122 17274
rect 18686 17222 18738 17274
rect 18790 17222 18842 17274
rect 18894 17222 18946 17274
rect 24510 17222 24562 17274
rect 24614 17222 24666 17274
rect 24718 17222 24770 17274
rect 2046 17054 2098 17106
rect 4398 17054 4450 17106
rect 16158 17054 16210 17106
rect 23102 17054 23154 17106
rect 1934 16942 1986 16994
rect 3054 16942 3106 16994
rect 3166 16942 3218 16994
rect 7870 16942 7922 16994
rect 9662 16942 9714 16994
rect 14254 16942 14306 16994
rect 14366 16942 14418 16994
rect 14814 16942 14866 16994
rect 16270 16942 16322 16994
rect 20638 16942 20690 16994
rect 4734 16830 4786 16882
rect 6302 16830 6354 16882
rect 11006 16830 11058 16882
rect 14702 16830 14754 16882
rect 15710 16830 15762 16882
rect 17390 16830 17442 16882
rect 23438 16830 23490 16882
rect 23662 16830 23714 16882
rect 23886 16830 23938 16882
rect 24222 16830 24274 16882
rect 3950 16718 4002 16770
rect 6750 16718 6802 16770
rect 7310 16718 7362 16770
rect 10110 16718 10162 16770
rect 10334 16718 10386 16770
rect 11790 16718 11842 16770
rect 13918 16718 13970 16770
rect 3054 16606 3106 16658
rect 5742 16606 5794 16658
rect 10446 16606 10498 16658
rect 4126 16438 4178 16490
rect 4230 16438 4282 16490
rect 4334 16438 4386 16490
rect 9950 16438 10002 16490
rect 10054 16438 10106 16490
rect 10158 16438 10210 16490
rect 15774 16438 15826 16490
rect 15878 16438 15930 16490
rect 15982 16438 16034 16490
rect 21598 16438 21650 16490
rect 21702 16438 21754 16490
rect 21806 16438 21858 16490
rect 2494 16270 2546 16322
rect 6078 16270 6130 16322
rect 6302 16270 6354 16322
rect 13582 16270 13634 16322
rect 21870 16270 21922 16322
rect 4174 16158 4226 16210
rect 4958 16158 5010 16210
rect 5070 16158 5122 16210
rect 9550 16158 9602 16210
rect 20190 16158 20242 16210
rect 20638 16158 20690 16210
rect 21310 16158 21362 16210
rect 2494 16046 2546 16098
rect 2718 16046 2770 16098
rect 3390 16046 3442 16098
rect 4062 16046 4114 16098
rect 5854 16046 5906 16098
rect 6526 16046 6578 16098
rect 8766 16046 8818 16098
rect 14590 16046 14642 16098
rect 15038 16046 15090 16098
rect 15822 16046 15874 16098
rect 16494 16046 16546 16098
rect 17278 16046 17330 16098
rect 21534 16046 21586 16098
rect 23102 16046 23154 16098
rect 23550 16046 23602 16098
rect 3054 15934 3106 15986
rect 3726 15934 3778 15986
rect 13582 15934 13634 15986
rect 13694 15934 13746 15986
rect 14142 15934 14194 15986
rect 15486 15934 15538 15986
rect 15598 15934 15650 15986
rect 18062 15934 18114 15986
rect 22542 15934 22594 15986
rect 24110 15934 24162 15986
rect 2606 15822 2658 15874
rect 3614 15822 3666 15874
rect 6414 15822 6466 15874
rect 16158 15822 16210 15874
rect 23214 15822 23266 15874
rect 7038 15654 7090 15706
rect 7142 15654 7194 15706
rect 7246 15654 7298 15706
rect 12862 15654 12914 15706
rect 12966 15654 13018 15706
rect 13070 15654 13122 15706
rect 18686 15654 18738 15706
rect 18790 15654 18842 15706
rect 18894 15654 18946 15706
rect 24510 15654 24562 15706
rect 24614 15654 24666 15706
rect 24718 15654 24770 15706
rect 6862 15486 6914 15538
rect 14254 15486 14306 15538
rect 15598 15486 15650 15538
rect 16270 15486 16322 15538
rect 21982 15486 22034 15538
rect 23998 15486 24050 15538
rect 3278 15374 3330 15426
rect 3838 15374 3890 15426
rect 5406 15374 5458 15426
rect 8094 15374 8146 15426
rect 8430 15374 8482 15426
rect 15038 15374 15090 15426
rect 15486 15374 15538 15426
rect 17390 15374 17442 15426
rect 20078 15374 20130 15426
rect 21758 15374 21810 15426
rect 22654 15374 22706 15426
rect 24110 15374 24162 15426
rect 2494 15262 2546 15314
rect 3166 15262 3218 15314
rect 4398 15262 4450 15314
rect 4734 15262 4786 15314
rect 6302 15262 6354 15314
rect 6638 15262 6690 15314
rect 7646 15262 7698 15314
rect 9550 15262 9602 15314
rect 14366 15262 14418 15314
rect 14590 15262 14642 15314
rect 14702 15262 14754 15314
rect 15710 15262 15762 15314
rect 16494 15262 16546 15314
rect 17614 15262 17666 15314
rect 20190 15262 20242 15314
rect 20414 15262 20466 15314
rect 20526 15262 20578 15314
rect 22318 15262 22370 15314
rect 22542 15262 22594 15314
rect 23550 15262 23602 15314
rect 4846 15150 4898 15202
rect 6750 15150 6802 15202
rect 7198 15150 7250 15202
rect 10334 15150 10386 15202
rect 12462 15150 12514 15202
rect 2158 15038 2210 15090
rect 21646 15038 21698 15090
rect 4126 14870 4178 14922
rect 4230 14870 4282 14922
rect 4334 14870 4386 14922
rect 9950 14870 10002 14922
rect 10054 14870 10106 14922
rect 10158 14870 10210 14922
rect 15774 14870 15826 14922
rect 15878 14870 15930 14922
rect 15982 14870 16034 14922
rect 21598 14870 21650 14922
rect 21702 14870 21754 14922
rect 21806 14870 21858 14922
rect 2046 14702 2098 14754
rect 14590 14702 14642 14754
rect 15598 14702 15650 14754
rect 10558 14590 10610 14642
rect 12910 14590 12962 14642
rect 15374 14590 15426 14642
rect 20414 14590 20466 14642
rect 21982 14590 22034 14642
rect 22766 14590 22818 14642
rect 23662 14590 23714 14642
rect 1934 14478 1986 14530
rect 2830 14478 2882 14530
rect 3166 14478 3218 14530
rect 4174 14478 4226 14530
rect 4622 14478 4674 14530
rect 4846 14478 4898 14530
rect 6750 14478 6802 14530
rect 7086 14478 7138 14530
rect 7758 14478 7810 14530
rect 8430 14478 8482 14530
rect 16382 14478 16434 14530
rect 16606 14478 16658 14530
rect 17502 14478 17554 14530
rect 22318 14478 22370 14530
rect 24222 14478 24274 14530
rect 1822 14366 1874 14418
rect 7198 14366 7250 14418
rect 14478 14366 14530 14418
rect 16718 14366 16770 14418
rect 18286 14366 18338 14418
rect 23886 14366 23938 14418
rect 2494 14254 2546 14306
rect 2606 14254 2658 14306
rect 2718 14254 2770 14306
rect 4398 14254 4450 14306
rect 12350 14254 12402 14306
rect 15934 14254 15986 14306
rect 17166 14254 17218 14306
rect 21422 14254 21474 14306
rect 7038 14086 7090 14138
rect 7142 14086 7194 14138
rect 7246 14086 7298 14138
rect 12862 14086 12914 14138
rect 12966 14086 13018 14138
rect 13070 14086 13122 14138
rect 18686 14086 18738 14138
rect 18790 14086 18842 14138
rect 18894 14086 18946 14138
rect 24510 14086 24562 14138
rect 24614 14086 24666 14138
rect 24718 14086 24770 14138
rect 6078 13918 6130 13970
rect 9886 13918 9938 13970
rect 17390 13918 17442 13970
rect 18286 13918 18338 13970
rect 23886 13918 23938 13970
rect 6862 13806 6914 13858
rect 6974 13806 7026 13858
rect 7758 13806 7810 13858
rect 14926 13806 14978 13858
rect 17950 13806 18002 13858
rect 19630 13806 19682 13858
rect 5070 13694 5122 13746
rect 5966 13694 6018 13746
rect 6190 13694 6242 13746
rect 6414 13694 6466 13746
rect 9550 13694 9602 13746
rect 11230 13694 11282 13746
rect 11566 13694 11618 13746
rect 19966 13694 20018 13746
rect 20414 13694 20466 13746
rect 24110 13694 24162 13746
rect 7982 13582 8034 13634
rect 8318 13582 8370 13634
rect 17502 13582 17554 13634
rect 21086 13582 21138 13634
rect 23214 13582 23266 13634
rect 5294 13470 5346 13522
rect 5630 13470 5682 13522
rect 6974 13470 7026 13522
rect 4126 13302 4178 13354
rect 4230 13302 4282 13354
rect 4334 13302 4386 13354
rect 9950 13302 10002 13354
rect 10054 13302 10106 13354
rect 10158 13302 10210 13354
rect 15774 13302 15826 13354
rect 15878 13302 15930 13354
rect 15982 13302 16034 13354
rect 21598 13302 21650 13354
rect 21702 13302 21754 13354
rect 21806 13302 21858 13354
rect 21310 13134 21362 13186
rect 2494 13022 2546 13074
rect 4622 13022 4674 13074
rect 8654 13022 8706 13074
rect 10782 13022 10834 13074
rect 14254 13022 14306 13074
rect 18286 13022 18338 13074
rect 20190 13022 20242 13074
rect 23886 13022 23938 13074
rect 1822 12910 1874 12962
rect 6190 12910 6242 12962
rect 7086 12910 7138 12962
rect 7870 12910 7922 12962
rect 17166 12910 17218 12962
rect 18958 12910 19010 12962
rect 19182 12910 19234 12962
rect 20526 12910 20578 12962
rect 21310 12910 21362 12962
rect 22990 12910 23042 12962
rect 23214 12910 23266 12962
rect 16382 12798 16434 12850
rect 20750 12798 20802 12850
rect 21646 12798 21698 12850
rect 22206 12798 22258 12850
rect 6526 12686 6578 12738
rect 6862 12686 6914 12738
rect 22542 12686 22594 12738
rect 7038 12518 7090 12570
rect 7142 12518 7194 12570
rect 7246 12518 7298 12570
rect 12862 12518 12914 12570
rect 12966 12518 13018 12570
rect 13070 12518 13122 12570
rect 18686 12518 18738 12570
rect 18790 12518 18842 12570
rect 18894 12518 18946 12570
rect 24510 12518 24562 12570
rect 24614 12518 24666 12570
rect 24718 12518 24770 12570
rect 15486 12350 15538 12402
rect 16718 12350 16770 12402
rect 19294 12350 19346 12402
rect 22766 12350 22818 12402
rect 6638 12238 6690 12290
rect 10334 12238 10386 12290
rect 10670 12238 10722 12290
rect 12462 12238 12514 12290
rect 16382 12238 16434 12290
rect 19742 12238 19794 12290
rect 20862 12238 20914 12290
rect 22206 12238 22258 12290
rect 23102 12238 23154 12290
rect 2046 12126 2098 12178
rect 5966 12126 6018 12178
rect 10894 12126 10946 12178
rect 11678 12126 11730 12178
rect 15038 12126 15090 12178
rect 15262 12126 15314 12178
rect 15598 12126 15650 12178
rect 16158 12126 16210 12178
rect 19182 12126 19234 12178
rect 20078 12126 20130 12178
rect 20302 12126 20354 12178
rect 20638 12126 20690 12178
rect 21758 12126 21810 12178
rect 23550 12126 23602 12178
rect 23998 12126 24050 12178
rect 2718 12014 2770 12066
rect 4846 12014 4898 12066
rect 8766 12014 8818 12066
rect 14590 12014 14642 12066
rect 15374 12014 15426 12066
rect 16830 12014 16882 12066
rect 20974 12014 21026 12066
rect 21310 12014 21362 12066
rect 11230 11902 11282 11954
rect 19294 11902 19346 11954
rect 4126 11734 4178 11786
rect 4230 11734 4282 11786
rect 4334 11734 4386 11786
rect 9950 11734 10002 11786
rect 10054 11734 10106 11786
rect 10158 11734 10210 11786
rect 15774 11734 15826 11786
rect 15878 11734 15930 11786
rect 15982 11734 16034 11786
rect 21598 11734 21650 11786
rect 21702 11734 21754 11786
rect 21806 11734 21858 11786
rect 13918 11566 13970 11618
rect 21198 11566 21250 11618
rect 3166 11454 3218 11506
rect 23774 11454 23826 11506
rect 3390 11342 3442 11394
rect 11454 11342 11506 11394
rect 14702 11342 14754 11394
rect 15486 11342 15538 11394
rect 21422 11342 21474 11394
rect 21870 11342 21922 11394
rect 22094 11342 22146 11394
rect 23102 11342 23154 11394
rect 23550 11342 23602 11394
rect 3054 11230 3106 11282
rect 9326 11230 9378 11282
rect 12686 11230 12738 11282
rect 13582 11230 13634 11282
rect 14478 11230 14530 11282
rect 17502 11230 17554 11282
rect 21982 11230 22034 11282
rect 22542 11230 22594 11282
rect 24110 11230 24162 11282
rect 12350 11118 12402 11170
rect 7038 10950 7090 11002
rect 7142 10950 7194 11002
rect 7246 10950 7298 11002
rect 12862 10950 12914 11002
rect 12966 10950 13018 11002
rect 13070 10950 13122 11002
rect 18686 10950 18738 11002
rect 18790 10950 18842 11002
rect 18894 10950 18946 11002
rect 24510 10950 24562 11002
rect 24614 10950 24666 11002
rect 24718 10950 24770 11002
rect 3166 10782 3218 10834
rect 14926 10782 14978 10834
rect 15934 10782 15986 10834
rect 16494 10782 16546 10834
rect 24222 10782 24274 10834
rect 2494 10670 2546 10722
rect 4286 10670 4338 10722
rect 5518 10670 5570 10722
rect 9774 10670 9826 10722
rect 10222 10670 10274 10722
rect 12126 10670 12178 10722
rect 22654 10670 22706 10722
rect 2270 10558 2322 10610
rect 3502 10558 3554 10610
rect 3950 10558 4002 10610
rect 4846 10558 4898 10610
rect 10446 10558 10498 10610
rect 11342 10558 11394 10610
rect 16382 10558 16434 10610
rect 17390 10558 17442 10610
rect 21422 10558 21474 10610
rect 21646 10558 21698 10610
rect 21982 10558 22034 10610
rect 23214 10558 23266 10610
rect 7646 10446 7698 10498
rect 14254 10446 14306 10498
rect 15486 10446 15538 10498
rect 18174 10446 18226 10498
rect 20302 10446 20354 10498
rect 21534 10446 21586 10498
rect 23438 10446 23490 10498
rect 10782 10334 10834 10386
rect 16270 10334 16322 10386
rect 4126 10166 4178 10218
rect 4230 10166 4282 10218
rect 4334 10166 4386 10218
rect 9950 10166 10002 10218
rect 10054 10166 10106 10218
rect 10158 10166 10210 10218
rect 15774 10166 15826 10218
rect 15878 10166 15930 10218
rect 15982 10166 16034 10218
rect 21598 10166 21650 10218
rect 21702 10166 21754 10218
rect 21806 10166 21858 10218
rect 18174 9998 18226 10050
rect 2494 9886 2546 9938
rect 4622 9886 4674 9938
rect 12014 9886 12066 9938
rect 19182 9886 19234 9938
rect 20302 9886 20354 9938
rect 24222 9886 24274 9938
rect 1822 9774 1874 9826
rect 8542 9774 8594 9826
rect 9214 9774 9266 9826
rect 15038 9774 15090 9826
rect 15262 9774 15314 9826
rect 19518 9774 19570 9826
rect 20526 9774 20578 9826
rect 20750 9774 20802 9826
rect 21310 9774 21362 9826
rect 9886 9662 9938 9714
rect 14814 9662 14866 9714
rect 18286 9662 18338 9714
rect 18510 9662 18562 9714
rect 18846 9662 18898 9714
rect 20190 9662 20242 9714
rect 22094 9662 22146 9714
rect 8766 9550 8818 9602
rect 14926 9550 14978 9602
rect 7038 9382 7090 9434
rect 7142 9382 7194 9434
rect 7246 9382 7298 9434
rect 12862 9382 12914 9434
rect 12966 9382 13018 9434
rect 13070 9382 13122 9434
rect 18686 9382 18738 9434
rect 18790 9382 18842 9434
rect 18894 9382 18946 9434
rect 24510 9382 24562 9434
rect 24614 9382 24666 9434
rect 24718 9382 24770 9434
rect 4510 9214 4562 9266
rect 7310 9214 7362 9266
rect 9662 9214 9714 9266
rect 16046 9214 16098 9266
rect 16382 9214 16434 9266
rect 20974 9214 21026 9266
rect 21198 9214 21250 9266
rect 22766 9214 22818 9266
rect 3838 9102 3890 9154
rect 5406 9102 5458 9154
rect 10334 9102 10386 9154
rect 10782 9102 10834 9154
rect 14702 9102 14754 9154
rect 18174 9102 18226 9154
rect 21870 9102 21922 9154
rect 24110 9102 24162 9154
rect 3950 8990 4002 9042
rect 4846 8990 4898 9042
rect 5630 8990 5682 9042
rect 7086 8990 7138 9042
rect 9998 8990 10050 9042
rect 11902 8990 11954 9042
rect 15486 8990 15538 9042
rect 15822 8990 15874 9042
rect 16270 8990 16322 9042
rect 17390 8990 17442 9042
rect 20750 8990 20802 9042
rect 21646 8990 21698 9042
rect 21982 8990 22034 9042
rect 23438 8990 23490 9042
rect 23886 8990 23938 9042
rect 11342 8878 11394 8930
rect 12574 8878 12626 8930
rect 16158 8878 16210 8930
rect 20302 8878 20354 8930
rect 22206 8878 22258 8930
rect 2830 8766 2882 8818
rect 3166 8766 3218 8818
rect 4126 8598 4178 8650
rect 4230 8598 4282 8650
rect 4334 8598 4386 8650
rect 9950 8598 10002 8650
rect 10054 8598 10106 8650
rect 10158 8598 10210 8650
rect 15774 8598 15826 8650
rect 15878 8598 15930 8650
rect 15982 8598 16034 8650
rect 21598 8598 21650 8650
rect 21702 8598 21754 8650
rect 21806 8598 21858 8650
rect 20302 8430 20354 8482
rect 21646 8430 21698 8482
rect 22094 8430 22146 8482
rect 4622 8318 4674 8370
rect 7534 8318 7586 8370
rect 9662 8318 9714 8370
rect 10110 8318 10162 8370
rect 11790 8318 11842 8370
rect 15262 8318 15314 8370
rect 15374 8318 15426 8370
rect 15710 8318 15762 8370
rect 23102 8318 23154 8370
rect 23550 8318 23602 8370
rect 1822 8206 1874 8258
rect 6862 8206 6914 8258
rect 10446 8206 10498 8258
rect 19630 8206 19682 8258
rect 19854 8206 19906 8258
rect 21758 8206 21810 8258
rect 21982 8206 22034 8258
rect 22542 8206 22594 8258
rect 23774 8206 23826 8258
rect 2494 8094 2546 8146
rect 11006 8094 11058 8146
rect 11566 8094 11618 8146
rect 19742 8094 19794 8146
rect 22766 8094 22818 8146
rect 12126 7982 12178 8034
rect 15822 7982 15874 8034
rect 7038 7814 7090 7866
rect 7142 7814 7194 7866
rect 7246 7814 7298 7866
rect 12862 7814 12914 7866
rect 12966 7814 13018 7866
rect 13070 7814 13122 7866
rect 18686 7814 18738 7866
rect 18790 7814 18842 7866
rect 18894 7814 18946 7866
rect 24510 7814 24562 7866
rect 24614 7814 24666 7866
rect 24718 7814 24770 7866
rect 2494 7646 2546 7698
rect 3838 7646 3890 7698
rect 19742 7646 19794 7698
rect 21534 7646 21586 7698
rect 22654 7646 22706 7698
rect 4958 7534 5010 7586
rect 6638 7534 6690 7586
rect 7198 7534 7250 7586
rect 7758 7534 7810 7586
rect 8318 7534 8370 7586
rect 10558 7534 10610 7586
rect 11118 7534 11170 7586
rect 12574 7534 12626 7586
rect 16046 7534 16098 7586
rect 21310 7534 21362 7586
rect 22878 7534 22930 7586
rect 2270 7422 2322 7474
rect 4174 7422 4226 7474
rect 4846 7422 4898 7474
rect 6414 7422 6466 7474
rect 7534 7422 7586 7474
rect 10334 7422 10386 7474
rect 12014 7422 12066 7474
rect 12798 7422 12850 7474
rect 16830 7422 16882 7474
rect 20078 7422 20130 7474
rect 23326 7422 23378 7474
rect 13918 7310 13970 7362
rect 21646 7310 21698 7362
rect 23662 7310 23714 7362
rect 5518 7198 5570 7250
rect 5854 7198 5906 7250
rect 9998 7198 10050 7250
rect 11678 7198 11730 7250
rect 4126 7030 4178 7082
rect 4230 7030 4282 7082
rect 4334 7030 4386 7082
rect 9950 7030 10002 7082
rect 10054 7030 10106 7082
rect 10158 7030 10210 7082
rect 15774 7030 15826 7082
rect 15878 7030 15930 7082
rect 15982 7030 16034 7082
rect 21598 7030 21650 7082
rect 21702 7030 21754 7082
rect 21806 7030 21858 7082
rect 9214 6862 9266 6914
rect 19966 6750 20018 6802
rect 20750 6750 20802 6802
rect 24222 6750 24274 6802
rect 4734 6638 4786 6690
rect 8318 6638 8370 6690
rect 8878 6638 8930 6690
rect 9998 6638 10050 6690
rect 11790 6638 11842 6690
rect 17054 6638 17106 6690
rect 21422 6638 21474 6690
rect 9774 6526 9826 6578
rect 17838 6526 17890 6578
rect 20414 6526 20466 6578
rect 20638 6526 20690 6578
rect 22094 6526 22146 6578
rect 4398 6414 4450 6466
rect 7982 6414 8034 6466
rect 12126 6414 12178 6466
rect 7038 6246 7090 6298
rect 7142 6246 7194 6298
rect 7246 6246 7298 6298
rect 12862 6246 12914 6298
rect 12966 6246 13018 6298
rect 13070 6246 13122 6298
rect 18686 6246 18738 6298
rect 18790 6246 18842 6298
rect 18894 6246 18946 6298
rect 24510 6246 24562 6298
rect 24614 6246 24666 6298
rect 24718 6246 24770 6298
rect 18510 6078 18562 6130
rect 22766 6078 22818 6130
rect 4062 5966 4114 6018
rect 13470 5966 13522 6018
rect 18398 5966 18450 6018
rect 22430 5966 22482 6018
rect 24110 5966 24162 6018
rect 3390 5854 3442 5906
rect 14254 5854 14306 5906
rect 18734 5854 18786 5906
rect 19742 5854 19794 5906
rect 20414 5854 20466 5906
rect 23214 5854 23266 5906
rect 23662 5854 23714 5906
rect 6190 5742 6242 5794
rect 11342 5742 11394 5794
rect 20526 5742 20578 5794
rect 4126 5462 4178 5514
rect 4230 5462 4282 5514
rect 4334 5462 4386 5514
rect 9950 5462 10002 5514
rect 10054 5462 10106 5514
rect 10158 5462 10210 5514
rect 15774 5462 15826 5514
rect 15878 5462 15930 5514
rect 15982 5462 16034 5514
rect 21598 5462 21650 5514
rect 21702 5462 21754 5514
rect 21806 5462 21858 5514
rect 7758 5182 7810 5234
rect 9886 5182 9938 5234
rect 23662 5182 23714 5234
rect 6974 5070 7026 5122
rect 24222 5070 24274 5122
rect 23886 4958 23938 5010
rect 7038 4678 7090 4730
rect 7142 4678 7194 4730
rect 7246 4678 7298 4730
rect 12862 4678 12914 4730
rect 12966 4678 13018 4730
rect 13070 4678 13122 4730
rect 18686 4678 18738 4730
rect 18790 4678 18842 4730
rect 18894 4678 18946 4730
rect 24510 4678 24562 4730
rect 24614 4678 24666 4730
rect 24718 4678 24770 4730
rect 23886 4510 23938 4562
rect 24222 4286 24274 4338
rect 23662 4174 23714 4226
rect 4126 3894 4178 3946
rect 4230 3894 4282 3946
rect 4334 3894 4386 3946
rect 9950 3894 10002 3946
rect 10054 3894 10106 3946
rect 10158 3894 10210 3946
rect 15774 3894 15826 3946
rect 15878 3894 15930 3946
rect 15982 3894 16034 3946
rect 21598 3894 21650 3946
rect 21702 3894 21754 3946
rect 21806 3894 21858 3946
rect 23438 3390 23490 3442
rect 23662 3390 23714 3442
rect 23998 3390 24050 3442
rect 7038 3110 7090 3162
rect 7142 3110 7194 3162
rect 7246 3110 7298 3162
rect 12862 3110 12914 3162
rect 12966 3110 13018 3162
rect 13070 3110 13122 3162
rect 18686 3110 18738 3162
rect 18790 3110 18842 3162
rect 18894 3110 18946 3162
rect 24510 3110 24562 3162
rect 24614 3110 24666 3162
rect 24718 3110 24770 3162
<< metal2 >>
rect 4256 25200 4368 26000
rect 12768 25200 12880 26000
rect 21280 25200 21392 26000
rect 4284 22932 4340 25200
rect 4284 22876 4788 22932
rect 4124 22764 4388 22774
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4124 22698 4388 22708
rect 2268 21364 2324 21374
rect 2268 20804 2324 21308
rect 4124 21196 4388 21206
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4124 21130 4388 21140
rect 1820 20802 2324 20804
rect 1820 20750 2270 20802
rect 2322 20750 2324 20802
rect 1820 20748 2324 20750
rect 1820 18450 1876 20748
rect 2268 20738 2324 20748
rect 2940 20690 2996 20702
rect 2940 20638 2942 20690
rect 2994 20638 2996 20690
rect 2940 20188 2996 20638
rect 2044 20132 2996 20188
rect 1820 18398 1822 18450
rect 1874 18398 1876 18450
rect 1820 18386 1876 18398
rect 1932 18564 1988 18574
rect 1932 16994 1988 18508
rect 1932 16942 1934 16994
rect 1986 16942 1988 16994
rect 1932 16930 1988 16942
rect 2044 17106 2100 20132
rect 4396 20018 4452 20030
rect 4396 19966 4398 20018
rect 4450 19966 4452 20018
rect 4396 19796 4452 19966
rect 3948 19740 4452 19796
rect 4508 19906 4564 19918
rect 4508 19854 4510 19906
rect 4562 19854 4564 19906
rect 3276 19124 3332 19134
rect 2940 19122 3332 19124
rect 2940 19070 3278 19122
rect 3330 19070 3332 19122
rect 2940 19068 3332 19070
rect 2940 18564 2996 19068
rect 3276 19058 3332 19068
rect 3948 19122 4004 19740
rect 4124 19628 4388 19638
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4124 19562 4388 19572
rect 4396 19234 4452 19246
rect 4396 19182 4398 19234
rect 4450 19182 4452 19234
rect 3948 19070 3950 19122
rect 4002 19070 4004 19122
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2492 17892 2548 18286
rect 2492 17826 2548 17836
rect 2940 17666 2996 18508
rect 3612 18452 3668 18462
rect 2940 17614 2942 17666
rect 2994 17614 2996 17666
rect 2940 17602 2996 17614
rect 3164 18228 3220 18238
rect 2044 17054 2046 17106
rect 2098 17054 2100 17106
rect 2044 16324 2100 17054
rect 2044 16258 2100 16268
rect 2380 17442 2436 17454
rect 2380 17390 2382 17442
rect 2434 17390 2436 17442
rect 2380 16100 2436 17390
rect 3052 16996 3108 17006
rect 2940 16994 3108 16996
rect 2940 16942 3054 16994
rect 3106 16942 3108 16994
rect 2940 16940 3108 16942
rect 2940 16772 2996 16940
rect 3052 16930 3108 16940
rect 3164 16996 3220 18172
rect 3612 17890 3668 18396
rect 3612 17838 3614 17890
rect 3666 17838 3668 17890
rect 3612 17826 3668 17838
rect 3836 18340 3892 18350
rect 3836 17778 3892 18284
rect 3836 17726 3838 17778
rect 3890 17726 3892 17778
rect 3836 17714 3892 17726
rect 3948 17556 4004 19070
rect 4284 19122 4340 19134
rect 4284 19070 4286 19122
rect 4338 19070 4340 19122
rect 4284 18340 4340 19070
rect 4396 18452 4452 19182
rect 4396 18386 4452 18396
rect 4284 18274 4340 18284
rect 4124 18060 4388 18070
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4124 17994 4388 18004
rect 3948 17490 4004 17500
rect 4284 17892 4340 17902
rect 3164 16902 3220 16940
rect 3276 17442 3332 17454
rect 3276 17390 3278 17442
rect 3330 17390 3332 17442
rect 2716 16716 2996 16772
rect 2492 16324 2548 16362
rect 2492 16258 2548 16268
rect 2044 15316 2100 15326
rect 1820 15092 1876 15102
rect 1820 14418 1876 15036
rect 2044 14754 2100 15260
rect 2380 15316 2436 16044
rect 2492 16098 2548 16110
rect 2492 16046 2494 16098
rect 2546 16046 2548 16098
rect 2492 15876 2548 16046
rect 2716 16098 2772 16716
rect 3052 16660 3108 16670
rect 2716 16046 2718 16098
rect 2770 16046 2772 16098
rect 2492 15810 2548 15820
rect 2604 15874 2660 15886
rect 2604 15822 2606 15874
rect 2658 15822 2660 15874
rect 2492 15316 2548 15326
rect 2436 15314 2548 15316
rect 2436 15262 2494 15314
rect 2546 15262 2548 15314
rect 2436 15260 2548 15262
rect 2380 15222 2436 15260
rect 2492 15250 2548 15260
rect 2044 14702 2046 14754
rect 2098 14702 2100 14754
rect 2044 14690 2100 14702
rect 2156 15090 2212 15102
rect 2156 15038 2158 15090
rect 2210 15038 2212 15090
rect 1932 14532 1988 14542
rect 1932 14438 1988 14476
rect 1820 14366 1822 14418
rect 1874 14366 1876 14418
rect 1820 14354 1876 14366
rect 2156 14308 2212 15038
rect 2604 14980 2660 15822
rect 2716 15428 2772 16046
rect 2940 16658 3108 16660
rect 2940 16606 3054 16658
rect 3106 16606 3108 16658
rect 2940 16604 3108 16606
rect 2940 15540 2996 16604
rect 3052 16594 3108 16604
rect 2716 15362 2772 15372
rect 2828 15484 2996 15540
rect 3052 15986 3108 15998
rect 3052 15934 3054 15986
rect 3106 15934 3108 15986
rect 2604 14914 2660 14924
rect 2828 14530 2884 15484
rect 3052 15092 3108 15934
rect 3276 15540 3332 17390
rect 4284 17442 4340 17836
rect 4396 17668 4452 17678
rect 4508 17668 4564 19854
rect 4620 18564 4676 18574
rect 4620 18338 4676 18508
rect 4620 18286 4622 18338
rect 4674 18286 4676 18338
rect 4620 18274 4676 18286
rect 4396 17666 4676 17668
rect 4396 17614 4398 17666
rect 4450 17614 4676 17666
rect 4396 17612 4676 17614
rect 4396 17602 4452 17612
rect 4284 17390 4286 17442
rect 4338 17390 4340 17442
rect 3724 16996 3780 17006
rect 3388 16324 3444 16334
rect 3388 16098 3444 16268
rect 3388 16046 3390 16098
rect 3442 16046 3444 16098
rect 3388 16034 3444 16046
rect 3724 15986 3780 16940
rect 3948 16770 4004 16782
rect 3948 16718 3950 16770
rect 4002 16718 4004 16770
rect 3948 16100 4004 16718
rect 4284 16660 4340 17390
rect 4396 17108 4452 17118
rect 4396 17014 4452 17052
rect 4620 16884 4676 17612
rect 4732 17444 4788 22876
rect 9948 22764 10212 22774
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 9948 22698 10212 22708
rect 12684 22484 12740 22494
rect 12796 22484 12852 25200
rect 20300 24052 20356 24062
rect 15772 22764 16036 22774
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 15772 22698 16036 22708
rect 12684 22482 13412 22484
rect 12684 22430 12686 22482
rect 12738 22430 13412 22482
rect 12684 22428 13412 22430
rect 12684 22418 12740 22428
rect 13356 22370 13412 22428
rect 13356 22318 13358 22370
rect 13410 22318 13412 22370
rect 13356 22306 13412 22318
rect 19628 22372 19684 22382
rect 19964 22372 20020 22382
rect 20300 22372 20356 23996
rect 21308 22596 21364 25200
rect 21596 22764 21860 22774
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21596 22698 21860 22708
rect 21308 22530 21364 22540
rect 22428 22596 22484 22606
rect 22428 22502 22484 22540
rect 19628 22370 20356 22372
rect 19628 22318 19630 22370
rect 19682 22318 19966 22370
rect 20018 22318 20356 22370
rect 19628 22316 20356 22318
rect 20860 22370 20916 22382
rect 20860 22318 20862 22370
rect 20914 22318 20916 22370
rect 19628 22306 19684 22316
rect 19964 22306 20020 22316
rect 13132 22148 13188 22158
rect 18732 22148 18788 22158
rect 12012 22146 13188 22148
rect 12012 22094 13134 22146
rect 13186 22094 13188 22146
rect 12012 22092 13188 22094
rect 7036 21980 7300 21990
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7036 21914 7300 21924
rect 7644 21812 7700 21822
rect 5068 21586 5124 21598
rect 5068 21534 5070 21586
rect 5122 21534 5124 21586
rect 5068 21364 5124 21534
rect 5068 21298 5124 21308
rect 5740 21474 5796 21486
rect 5740 21422 5742 21474
rect 5794 21422 5796 21474
rect 5068 20916 5124 20926
rect 5068 20914 5348 20916
rect 5068 20862 5070 20914
rect 5122 20862 5348 20914
rect 5068 20860 5348 20862
rect 5068 20850 5124 20860
rect 4956 20132 5012 20142
rect 4956 20130 5236 20132
rect 4956 20078 4958 20130
rect 5010 20078 5236 20130
rect 4956 20076 5236 20078
rect 4956 20066 5012 20076
rect 5180 18676 5236 20076
rect 5292 19908 5348 20860
rect 5404 19908 5460 19918
rect 5292 19852 5404 19908
rect 5404 19842 5460 19852
rect 5180 18562 5236 18620
rect 5180 18510 5182 18562
rect 5234 18510 5236 18562
rect 5180 18498 5236 18510
rect 4956 18452 5012 18462
rect 4956 18358 5012 18396
rect 5516 18450 5572 18462
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 4844 18228 4900 18238
rect 4844 18134 4900 18172
rect 5516 18228 5572 18398
rect 5516 18162 5572 18172
rect 5628 18452 5684 18462
rect 5628 17778 5684 18396
rect 5628 17726 5630 17778
rect 5682 17726 5684 17778
rect 5628 17714 5684 17726
rect 4732 17388 4900 17444
rect 4732 16884 4788 16894
rect 4620 16882 4788 16884
rect 4620 16830 4734 16882
rect 4786 16830 4788 16882
rect 4620 16828 4788 16830
rect 4732 16818 4788 16828
rect 4284 16604 4564 16660
rect 4124 16492 4388 16502
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4124 16426 4388 16436
rect 4172 16210 4228 16222
rect 4172 16158 4174 16210
rect 4226 16158 4228 16210
rect 4060 16100 4116 16110
rect 3948 16098 4116 16100
rect 3948 16046 4062 16098
rect 4114 16046 4116 16098
rect 3948 16044 4116 16046
rect 3724 15934 3726 15986
rect 3778 15934 3780 15986
rect 3724 15922 3780 15934
rect 3612 15876 3668 15886
rect 3612 15782 3668 15820
rect 3276 15484 3892 15540
rect 3276 15426 3332 15484
rect 3276 15374 3278 15426
rect 3330 15374 3332 15426
rect 3276 15362 3332 15374
rect 3836 15426 3892 15484
rect 3836 15374 3838 15426
rect 3890 15374 3892 15426
rect 3836 15362 3892 15374
rect 3164 15316 3220 15326
rect 3164 15222 3220 15260
rect 4060 15316 4116 16044
rect 4060 15250 4116 15260
rect 4172 15148 4228 16158
rect 4508 15876 4564 16604
rect 4844 15988 4900 17388
rect 4956 17108 5012 17118
rect 4956 16210 5012 17052
rect 5740 16884 5796 21422
rect 7644 20690 7700 21756
rect 8204 21812 8260 21822
rect 8204 21718 8260 21756
rect 8428 21586 8484 21598
rect 8428 21534 8430 21586
rect 8482 21534 8484 21586
rect 7868 21476 7924 21486
rect 8428 21476 8484 21534
rect 7868 21474 8484 21476
rect 7868 21422 7870 21474
rect 7922 21422 8484 21474
rect 7868 21420 8484 21422
rect 7868 21410 7924 21420
rect 7644 20638 7646 20690
rect 7698 20638 7700 20690
rect 7036 20412 7300 20422
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7036 20346 7300 20356
rect 7644 20356 7700 20638
rect 7868 20804 7924 20814
rect 7756 20580 7812 20590
rect 7756 20486 7812 20524
rect 7644 20290 7700 20300
rect 6748 20244 6804 20254
rect 6748 20150 6804 20188
rect 7756 20020 7812 20030
rect 7868 20020 7924 20748
rect 8092 20802 8148 20814
rect 8092 20750 8094 20802
rect 8146 20750 8148 20802
rect 8092 20244 8148 20750
rect 8316 20692 8372 20702
rect 8428 20692 8484 21420
rect 9660 21586 9716 21598
rect 9660 21534 9662 21586
rect 9714 21534 9716 21586
rect 9660 21364 9716 21534
rect 10444 21476 10500 21486
rect 10444 21474 10724 21476
rect 10444 21422 10446 21474
rect 10498 21422 10724 21474
rect 10444 21420 10724 21422
rect 10444 21410 10500 21420
rect 8876 21026 8932 21038
rect 8876 20974 8878 21026
rect 8930 20974 8932 21026
rect 8652 20804 8708 20814
rect 8652 20710 8708 20748
rect 8316 20690 8484 20692
rect 8316 20638 8318 20690
rect 8370 20638 8484 20690
rect 8316 20636 8484 20638
rect 8316 20626 8372 20636
rect 8428 20468 8484 20478
rect 8316 20356 8372 20366
rect 8092 20178 8148 20188
rect 8204 20300 8316 20356
rect 7532 20018 7924 20020
rect 7532 19966 7758 20018
rect 7810 19966 7924 20018
rect 7532 19964 7924 19966
rect 7980 20020 8036 20030
rect 8204 20020 8260 20300
rect 8316 20290 8372 20300
rect 8428 20132 8484 20412
rect 8876 20244 8932 20974
rect 9324 20804 9380 20814
rect 6636 19908 6692 19918
rect 6412 18450 6468 18462
rect 6412 18398 6414 18450
rect 6466 18398 6468 18450
rect 6412 18340 6468 18398
rect 6636 18340 6692 19852
rect 7084 19906 7140 19918
rect 7084 19854 7086 19906
rect 7138 19854 7140 19906
rect 7084 19012 7140 19854
rect 7532 19458 7588 19964
rect 7756 19954 7812 19964
rect 7980 19926 8036 19964
rect 8092 19964 8260 20020
rect 8316 20076 8484 20132
rect 8764 20242 8932 20244
rect 8764 20190 8878 20242
rect 8930 20190 8932 20242
rect 8764 20188 8932 20190
rect 7532 19406 7534 19458
rect 7586 19406 7588 19458
rect 7532 19394 7588 19406
rect 7420 19236 7476 19246
rect 7868 19236 7924 19246
rect 7420 19234 7924 19236
rect 7420 19182 7422 19234
rect 7474 19182 7870 19234
rect 7922 19182 7924 19234
rect 7420 19180 7924 19182
rect 7420 19170 7476 19180
rect 6860 18956 7140 19012
rect 6748 18676 6804 18686
rect 6860 18676 6916 18956
rect 7036 18844 7300 18854
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7036 18778 7300 18788
rect 6860 18620 7588 18676
rect 6748 18452 6804 18620
rect 6860 18452 6916 18462
rect 6748 18450 6916 18452
rect 6748 18398 6862 18450
rect 6914 18398 6916 18450
rect 6748 18396 6916 18398
rect 6860 18386 6916 18396
rect 7196 18450 7252 18620
rect 7196 18398 7198 18450
rect 7250 18398 7252 18450
rect 7196 18386 7252 18398
rect 7308 18452 7364 18462
rect 6636 18284 6804 18340
rect 6412 18274 6468 18284
rect 6748 17666 6804 18284
rect 6748 17614 6750 17666
rect 6802 17614 6804 17666
rect 6748 17602 6804 17614
rect 7196 17668 7252 17678
rect 7308 17668 7364 18396
rect 7196 17666 7364 17668
rect 7196 17614 7198 17666
rect 7250 17614 7364 17666
rect 7196 17612 7364 17614
rect 7196 17602 7252 17612
rect 7036 17276 7300 17286
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7036 17210 7300 17220
rect 6300 16884 6356 16894
rect 5628 16828 5740 16884
rect 5180 16324 5236 16334
rect 4956 16158 4958 16210
rect 5010 16158 5012 16210
rect 4956 16146 5012 16158
rect 5068 16268 5180 16324
rect 5068 16210 5124 16268
rect 5180 16258 5236 16268
rect 5068 16158 5070 16210
rect 5122 16158 5124 16210
rect 5068 16146 5124 16158
rect 4844 15932 5012 15988
rect 4732 15876 4788 15886
rect 4508 15820 4732 15876
rect 4620 15428 4676 15438
rect 4396 15316 4452 15326
rect 4396 15222 4452 15260
rect 3052 15026 3108 15036
rect 3948 15092 4228 15148
rect 3164 14980 3220 14990
rect 3220 14924 3332 14980
rect 3164 14914 3220 14924
rect 2828 14478 2830 14530
rect 2882 14478 2884 14530
rect 2828 14466 2884 14478
rect 2940 14532 2996 14542
rect 3164 14532 3220 14542
rect 2996 14530 3220 14532
rect 2996 14478 3166 14530
rect 3218 14478 3220 14530
rect 2996 14476 3220 14478
rect 2940 14466 2996 14476
rect 3164 14466 3220 14476
rect 2492 14308 2548 14318
rect 2156 14306 2548 14308
rect 2156 14254 2494 14306
rect 2546 14254 2548 14306
rect 2156 14252 2548 14254
rect 2492 14242 2548 14252
rect 2604 14306 2660 14318
rect 2604 14254 2606 14306
rect 2658 14254 2660 14306
rect 2492 13076 2548 13086
rect 2604 13076 2660 14254
rect 2716 14306 2772 14318
rect 2716 14254 2718 14306
rect 2770 14254 2772 14306
rect 2716 13636 2772 14254
rect 2716 13570 2772 13580
rect 2492 13074 2660 13076
rect 2492 13022 2494 13074
rect 2546 13022 2660 13074
rect 2492 13020 2660 13022
rect 2492 13010 2548 13020
rect 1820 12962 1876 12974
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1820 12180 1876 12910
rect 2044 12180 2100 12190
rect 1820 12178 2100 12180
rect 1820 12126 2046 12178
rect 2098 12126 2100 12178
rect 1820 12124 2100 12126
rect 2044 10612 2100 12124
rect 2716 12068 2772 12078
rect 2716 12066 3220 12068
rect 2716 12014 2718 12066
rect 2770 12014 3220 12066
rect 2716 12012 3220 12014
rect 2716 12002 2772 12012
rect 3164 11506 3220 12012
rect 3164 11454 3166 11506
rect 3218 11454 3220 11506
rect 3164 11442 3220 11454
rect 3052 11284 3108 11294
rect 3276 11284 3332 14924
rect 3948 14532 4004 15092
rect 4124 14924 4388 14934
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4124 14858 4388 14868
rect 4172 14532 4228 14542
rect 3948 14530 4228 14532
rect 3948 14478 4174 14530
rect 4226 14478 4228 14530
rect 3948 14476 4228 14478
rect 4172 14466 4228 14476
rect 4620 14530 4676 15372
rect 4732 15314 4788 15820
rect 4732 15262 4734 15314
rect 4786 15262 4788 15314
rect 4732 15250 4788 15262
rect 4620 14478 4622 14530
rect 4674 14478 4676 14530
rect 4620 14466 4676 14478
rect 4844 15202 4900 15214
rect 4844 15150 4846 15202
rect 4898 15150 4900 15202
rect 4844 14530 4900 15150
rect 4844 14478 4846 14530
rect 4898 14478 4900 14530
rect 4396 14308 4452 14318
rect 4396 14214 4452 14252
rect 4844 13748 4900 14478
rect 4956 13972 5012 15932
rect 5516 15876 5572 15886
rect 5404 15428 5460 15438
rect 5516 15428 5572 15820
rect 5460 15372 5572 15428
rect 5404 15334 5460 15372
rect 5628 15092 5684 16828
rect 5740 16818 5796 16828
rect 6076 16882 6356 16884
rect 6076 16830 6302 16882
rect 6354 16830 6356 16882
rect 6076 16828 6356 16830
rect 5740 16660 5796 16670
rect 5740 16566 5796 16604
rect 6076 16324 6132 16828
rect 6300 16818 6356 16828
rect 6748 16884 6804 16894
rect 6748 16770 6804 16828
rect 6748 16718 6750 16770
rect 6802 16718 6804 16770
rect 6748 16706 6804 16718
rect 7308 16770 7364 16782
rect 7308 16718 7310 16770
rect 7362 16718 7364 16770
rect 6076 16230 6132 16268
rect 6300 16660 6356 16670
rect 6300 16324 6356 16604
rect 6300 16322 6916 16324
rect 6300 16270 6302 16322
rect 6354 16270 6916 16322
rect 6300 16268 6916 16270
rect 6300 16258 6356 16268
rect 5852 16100 5908 16110
rect 6524 16100 6580 16110
rect 5908 16044 6356 16100
rect 5852 16006 5908 16044
rect 6300 15314 6356 16044
rect 6524 16006 6580 16044
rect 6412 15876 6468 15886
rect 6412 15874 6580 15876
rect 6412 15822 6414 15874
rect 6466 15822 6580 15874
rect 6412 15820 6580 15822
rect 6412 15810 6468 15820
rect 6300 15262 6302 15314
rect 6354 15262 6356 15314
rect 6300 15250 6356 15262
rect 5628 14084 5684 15036
rect 6412 14532 6468 14542
rect 5628 14028 6020 14084
rect 4956 13906 5012 13916
rect 5068 13748 5124 13758
rect 4844 13746 5124 13748
rect 4844 13694 5070 13746
rect 5122 13694 5124 13746
rect 4844 13692 5124 13694
rect 5068 13682 5124 13692
rect 5964 13746 6020 14028
rect 5964 13694 5966 13746
rect 6018 13694 6020 13746
rect 5964 13682 6020 13694
rect 6076 13970 6132 13982
rect 6076 13918 6078 13970
rect 6130 13918 6132 13970
rect 5292 13524 5348 13534
rect 5292 13430 5348 13468
rect 5628 13524 5684 13534
rect 6076 13524 6132 13918
rect 6188 13860 6244 13870
rect 6188 13746 6244 13804
rect 6188 13694 6190 13746
rect 6242 13694 6244 13746
rect 6188 13682 6244 13694
rect 6412 13748 6468 14476
rect 6524 14308 6580 15820
rect 6860 15538 6916 16268
rect 7308 15876 7364 16718
rect 7308 15810 7364 15820
rect 7036 15708 7300 15718
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7036 15642 7300 15652
rect 6860 15486 6862 15538
rect 6914 15486 6916 15538
rect 6636 15316 6692 15326
rect 6636 15222 6692 15260
rect 6748 15202 6804 15214
rect 6748 15150 6750 15202
rect 6802 15150 6804 15202
rect 6748 14530 6804 15150
rect 6748 14478 6750 14530
rect 6802 14478 6804 14530
rect 6748 14466 6804 14478
rect 6524 14252 6804 14308
rect 6412 13654 6468 13692
rect 5628 13522 6020 13524
rect 5628 13470 5630 13522
rect 5682 13470 6020 13522
rect 5628 13468 6020 13470
rect 5628 13458 5684 13468
rect 4124 13356 4388 13366
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4124 13290 4388 13300
rect 5964 13188 6020 13468
rect 6076 13458 6132 13468
rect 5964 13132 6244 13188
rect 4620 13076 4676 13086
rect 4620 13074 4788 13076
rect 4620 13022 4622 13074
rect 4674 13022 4788 13074
rect 4620 13020 4788 13022
rect 4620 13010 4676 13020
rect 4124 11788 4388 11798
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4124 11722 4388 11732
rect 3388 11508 3444 11518
rect 3388 11394 3444 11452
rect 3388 11342 3390 11394
rect 3442 11342 3444 11394
rect 3388 11330 3444 11342
rect 3052 11282 3332 11284
rect 3052 11230 3054 11282
rect 3106 11230 3332 11282
rect 3052 11228 3332 11230
rect 3052 11218 3108 11228
rect 1820 9828 1876 9838
rect 2044 9828 2100 10556
rect 2268 10892 3220 10948
rect 2268 10610 2324 10892
rect 3164 10834 3220 10892
rect 3164 10782 3166 10834
rect 3218 10782 3220 10834
rect 3164 10770 3220 10782
rect 2268 10558 2270 10610
rect 2322 10558 2324 10610
rect 2268 10546 2324 10558
rect 2492 10722 2548 10734
rect 2492 10670 2494 10722
rect 2546 10670 2548 10722
rect 2492 9938 2548 10670
rect 3500 10724 3556 10734
rect 2492 9886 2494 9938
rect 2546 9886 2548 9938
rect 2492 9874 2548 9886
rect 3276 10612 3332 10622
rect 1820 9826 2100 9828
rect 1820 9774 1822 9826
rect 1874 9774 2100 9826
rect 1820 9772 2100 9774
rect 1820 9762 1876 9772
rect 2044 8428 2100 9772
rect 2828 8818 2884 8830
rect 2828 8766 2830 8818
rect 2882 8766 2884 8818
rect 2828 8428 2884 8766
rect 3164 8820 3220 8830
rect 3164 8726 3220 8764
rect 1820 8372 2100 8428
rect 2268 8372 2884 8428
rect 1820 8258 1876 8372
rect 1820 8206 1822 8258
rect 1874 8206 1876 8258
rect 1820 8194 1876 8206
rect 2268 7474 2324 8372
rect 2492 8146 2548 8158
rect 2492 8094 2494 8146
rect 2546 8094 2548 8146
rect 2492 7698 2548 8094
rect 2492 7646 2494 7698
rect 2546 7646 2548 7698
rect 2492 7634 2548 7646
rect 2268 7422 2270 7474
rect 2322 7422 2324 7474
rect 2268 7410 2324 7422
rect 3276 6804 3332 10556
rect 3500 10610 3556 10668
rect 4284 10724 4340 10734
rect 4620 10724 4676 10734
rect 4284 10722 4564 10724
rect 4284 10670 4286 10722
rect 4338 10670 4564 10722
rect 4284 10668 4564 10670
rect 4284 10658 4340 10668
rect 3500 10558 3502 10610
rect 3554 10558 3556 10610
rect 3500 10546 3556 10558
rect 3948 10610 4004 10622
rect 3948 10558 3950 10610
rect 4002 10558 4004 10610
rect 3948 9380 4004 10558
rect 4124 10220 4388 10230
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4124 10154 4388 10164
rect 3724 9324 4004 9380
rect 3724 8372 3780 9324
rect 3724 8306 3780 8316
rect 3836 9154 3892 9166
rect 3836 9102 3838 9154
rect 3890 9102 3892 9154
rect 3836 7698 3892 9102
rect 3948 9042 4004 9324
rect 4508 9266 4564 10668
rect 4620 9938 4676 10668
rect 4620 9886 4622 9938
rect 4674 9886 4676 9938
rect 4620 9874 4676 9886
rect 4508 9214 4510 9266
rect 4562 9214 4564 9266
rect 4508 9202 4564 9214
rect 3948 8990 3950 9042
rect 4002 8990 4004 9042
rect 3948 8978 4004 8990
rect 4124 8652 4388 8662
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4732 8596 4788 13020
rect 5964 12964 6020 12974
rect 5964 12178 6020 12908
rect 6188 12962 6244 13132
rect 6188 12910 6190 12962
rect 6242 12910 6244 12962
rect 6188 12898 6244 12910
rect 6748 12964 6804 14252
rect 6860 13860 6916 15486
rect 7196 15202 7252 15214
rect 7196 15150 7198 15202
rect 7250 15150 7252 15202
rect 7196 15148 7252 15150
rect 7084 15092 7252 15148
rect 7084 14532 7140 15092
rect 7084 14438 7140 14476
rect 7196 14420 7252 14430
rect 7196 14418 7476 14420
rect 7196 14366 7198 14418
rect 7250 14366 7476 14418
rect 7196 14364 7476 14366
rect 7196 14354 7252 14364
rect 7036 14140 7300 14150
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7036 14074 7300 14084
rect 6860 13766 6916 13804
rect 6972 13860 7028 13870
rect 6972 13858 7140 13860
rect 6972 13806 6974 13858
rect 7026 13806 7140 13858
rect 6972 13804 7140 13806
rect 6972 13794 7028 13804
rect 7084 13748 7140 13804
rect 7084 13682 7140 13692
rect 6972 13636 7028 13646
rect 6972 13522 7028 13580
rect 6972 13470 6974 13522
rect 7026 13470 7028 13522
rect 6972 13458 7028 13470
rect 7084 12964 7140 12974
rect 6748 12962 7140 12964
rect 6748 12910 7086 12962
rect 7138 12910 7140 12962
rect 6748 12908 7140 12910
rect 7084 12898 7140 12908
rect 6524 12740 6580 12750
rect 6524 12738 6692 12740
rect 6524 12686 6526 12738
rect 6578 12686 6692 12738
rect 6524 12684 6692 12686
rect 6524 12674 6580 12684
rect 6636 12290 6692 12684
rect 6636 12238 6638 12290
rect 6690 12238 6692 12290
rect 6636 12226 6692 12238
rect 6860 12738 6916 12750
rect 6860 12686 6862 12738
rect 6914 12686 6916 12738
rect 5964 12126 5966 12178
rect 6018 12126 6020 12178
rect 4844 12068 4900 12078
rect 4844 12066 5012 12068
rect 4844 12014 4846 12066
rect 4898 12014 5012 12066
rect 4844 12012 5012 12014
rect 4844 12002 4900 12012
rect 4844 11732 4900 11742
rect 4844 10612 4900 11676
rect 4844 10518 4900 10556
rect 4844 9044 4900 9054
rect 4956 9044 5012 12012
rect 5964 11732 6020 12126
rect 5964 11666 6020 11676
rect 5516 11508 5572 11518
rect 5516 10722 5572 11452
rect 6860 11508 6916 12686
rect 7036 12572 7300 12582
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7036 12506 7300 12516
rect 6860 11442 6916 11452
rect 5516 10670 5518 10722
rect 5570 10670 5572 10722
rect 5516 10658 5572 10670
rect 6860 11284 6916 11294
rect 4844 9042 5012 9044
rect 4844 8990 4846 9042
rect 4898 8990 5012 9042
rect 4844 8988 5012 8990
rect 5404 9154 5460 9166
rect 5404 9102 5406 9154
rect 5458 9102 5460 9154
rect 4844 8978 4900 8988
rect 4124 8586 4388 8596
rect 4508 8540 4788 8596
rect 4844 8820 4900 8830
rect 4508 8428 4564 8540
rect 4844 8428 4900 8764
rect 5404 8428 5460 9102
rect 3836 7646 3838 7698
rect 3890 7646 3892 7698
rect 3836 7634 3892 7646
rect 4172 8372 4564 8428
rect 4620 8372 5460 8428
rect 5628 9042 5684 9054
rect 5628 8990 5630 9042
rect 5682 8990 5684 9042
rect 4172 7474 4228 8372
rect 4620 8370 4676 8372
rect 4620 8318 4622 8370
rect 4674 8318 4676 8370
rect 4620 8306 4676 8318
rect 4956 7588 5012 7598
rect 4956 7494 5012 7532
rect 4172 7422 4174 7474
rect 4226 7422 4228 7474
rect 4172 7410 4228 7422
rect 4844 7476 4900 7486
rect 4844 7382 4900 7420
rect 5628 7476 5684 8990
rect 6412 8372 6468 8382
rect 5628 7410 5684 7420
rect 5852 7588 5908 7598
rect 4732 7252 4788 7262
rect 4124 7084 4388 7094
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4124 7018 4388 7028
rect 3276 6748 3444 6804
rect 3388 5906 3444 6748
rect 4732 6690 4788 7196
rect 5516 7252 5572 7262
rect 5516 7158 5572 7196
rect 5852 7250 5908 7532
rect 6412 7474 6468 8316
rect 6860 8258 6916 11228
rect 7036 11004 7300 11014
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7036 10938 7300 10948
rect 7036 9436 7300 9446
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7036 9370 7300 9380
rect 7420 9380 7476 14364
rect 7532 13860 7588 18620
rect 7756 18564 7812 18574
rect 7868 18564 7924 19180
rect 8092 19234 8148 19964
rect 8316 19908 8372 20076
rect 8092 19182 8094 19234
rect 8146 19182 8148 19234
rect 8092 19170 8148 19182
rect 8204 19236 8260 19246
rect 8316 19236 8372 19852
rect 8204 19234 8372 19236
rect 8204 19182 8206 19234
rect 8258 19182 8372 19234
rect 8204 19180 8372 19182
rect 8204 19170 8260 19180
rect 8652 19124 8708 19134
rect 8652 19030 8708 19068
rect 7812 18508 7924 18564
rect 7756 18470 7812 18508
rect 7980 18452 8036 18462
rect 8428 18452 8484 18462
rect 7980 18450 8484 18452
rect 7980 18398 7982 18450
rect 8034 18398 8430 18450
rect 8482 18398 8484 18450
rect 7980 18396 8484 18398
rect 7980 18386 8036 18396
rect 8428 18386 8484 18396
rect 8540 18228 8596 18238
rect 8540 17554 8596 18172
rect 8764 17666 8820 20188
rect 8876 20178 8932 20188
rect 9212 20802 9380 20804
rect 9212 20750 9326 20802
rect 9378 20750 9380 20802
rect 9212 20748 9380 20750
rect 8988 20020 9044 20030
rect 8988 20018 9156 20020
rect 8988 19966 8990 20018
rect 9042 19966 9156 20018
rect 8988 19964 9156 19966
rect 8988 19954 9044 19964
rect 8876 19796 8932 19806
rect 8876 19794 9044 19796
rect 8876 19742 8878 19794
rect 8930 19742 9044 19794
rect 8876 19740 9044 19742
rect 8876 19730 8932 19740
rect 8988 18676 9044 19740
rect 9100 19234 9156 19964
rect 9100 19182 9102 19234
rect 9154 19182 9156 19234
rect 9100 19170 9156 19182
rect 9212 19012 9268 20748
rect 9324 20738 9380 20748
rect 9548 20130 9604 20142
rect 9548 20078 9550 20130
rect 9602 20078 9604 20130
rect 9548 20020 9604 20078
rect 9548 19954 9604 19964
rect 9660 19348 9716 21308
rect 9948 21196 10212 21206
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 9948 21130 10212 21140
rect 9884 20690 9940 20702
rect 9884 20638 9886 20690
rect 9938 20638 9940 20690
rect 9884 20244 9940 20638
rect 10444 20690 10500 20702
rect 10444 20638 10446 20690
rect 10498 20638 10500 20690
rect 9996 20580 10052 20590
rect 10220 20580 10276 20590
rect 9996 20486 10052 20524
rect 10108 20578 10276 20580
rect 10108 20526 10222 20578
rect 10274 20526 10276 20578
rect 10108 20524 10276 20526
rect 10108 20244 10164 20524
rect 10220 20514 10276 20524
rect 10444 20468 10500 20638
rect 10444 20402 10500 20412
rect 10556 20578 10612 20590
rect 10556 20526 10558 20578
rect 10610 20526 10612 20578
rect 9884 20178 9940 20188
rect 9996 20188 10164 20244
rect 10556 20356 10612 20526
rect 9996 20130 10052 20188
rect 9996 20078 9998 20130
rect 10050 20078 10052 20130
rect 9996 20066 10052 20078
rect 9772 20018 9828 20030
rect 9772 19966 9774 20018
rect 9826 19966 9828 20018
rect 9772 19460 9828 19966
rect 9884 19908 9940 19918
rect 9884 19814 9940 19852
rect 9948 19628 10212 19638
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 9948 19562 10212 19572
rect 9772 19404 9940 19460
rect 9548 19292 9716 19348
rect 9436 19124 9492 19134
rect 9436 19030 9492 19068
rect 9324 19012 9380 19022
rect 9212 18956 9324 19012
rect 9324 18918 9380 18956
rect 9548 18788 9604 19292
rect 9772 19124 9828 19134
rect 9772 19030 9828 19068
rect 9548 18732 9716 18788
rect 8988 18620 9604 18676
rect 8988 18452 9044 18462
rect 8988 18358 9044 18396
rect 9324 17892 9380 17902
rect 9324 17778 9380 17836
rect 9548 17890 9604 18620
rect 9548 17838 9550 17890
rect 9602 17838 9604 17890
rect 9548 17826 9604 17838
rect 9324 17726 9326 17778
rect 9378 17726 9380 17778
rect 9324 17714 9380 17726
rect 9660 17668 9716 18732
rect 9772 18452 9828 18462
rect 9772 18338 9828 18396
rect 9772 18286 9774 18338
rect 9826 18286 9828 18338
rect 9772 18274 9828 18286
rect 9884 18228 9940 19404
rect 10556 19236 10612 20300
rect 10668 19460 10724 21420
rect 10780 20578 10836 20590
rect 10780 20526 10782 20578
rect 10834 20526 10836 20578
rect 10780 20020 10836 20526
rect 11340 20132 11396 20142
rect 11340 20130 11508 20132
rect 11340 20078 11342 20130
rect 11394 20078 11508 20130
rect 11340 20076 11508 20078
rect 11340 20066 11396 20076
rect 10780 19954 10836 19964
rect 11228 20018 11284 20030
rect 11228 19966 11230 20018
rect 11282 19966 11284 20018
rect 11228 19908 11284 19966
rect 11228 19842 11284 19852
rect 10668 19394 10724 19404
rect 10668 19236 10724 19246
rect 10556 19234 10724 19236
rect 10556 19182 10670 19234
rect 10722 19182 10724 19234
rect 10556 19180 10724 19182
rect 10668 19170 10724 19180
rect 10892 19234 10948 19246
rect 10892 19182 10894 19234
rect 10946 19182 10948 19234
rect 10108 19124 10164 19134
rect 10108 19030 10164 19068
rect 10332 19124 10388 19134
rect 10892 19124 10948 19182
rect 10332 19122 10612 19124
rect 10332 19070 10334 19122
rect 10386 19070 10612 19122
rect 10332 19068 10612 19070
rect 9996 19010 10052 19022
rect 9996 18958 9998 19010
rect 10050 18958 10052 19010
rect 9996 18228 10052 18958
rect 10332 19012 10388 19068
rect 10332 18946 10388 18956
rect 9996 18172 10388 18228
rect 9884 18162 9940 18172
rect 9948 18060 10212 18070
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 9948 17994 10212 18004
rect 8764 17614 8766 17666
rect 8818 17614 8820 17666
rect 8764 17602 8820 17614
rect 9548 17612 9716 17668
rect 8540 17502 8542 17554
rect 8594 17502 8596 17554
rect 8540 17490 8596 17502
rect 7868 16996 7924 17006
rect 7868 16902 7924 16940
rect 8428 16996 8484 17006
rect 7644 16100 7700 16110
rect 7644 15428 7700 16044
rect 8092 15428 8148 15438
rect 7644 15426 8148 15428
rect 7644 15374 8094 15426
rect 8146 15374 8148 15426
rect 7644 15372 8148 15374
rect 7644 15314 7700 15372
rect 8092 15362 8148 15372
rect 8428 15426 8484 16940
rect 9548 16772 9604 17612
rect 9884 17444 9940 17454
rect 9884 17442 10052 17444
rect 9884 17390 9886 17442
rect 9938 17390 10052 17442
rect 9884 17388 10052 17390
rect 9884 17378 9940 17388
rect 9660 16996 9716 17006
rect 9660 16902 9716 16940
rect 9996 16772 10052 17388
rect 10108 16772 10164 16782
rect 9996 16770 10164 16772
rect 9996 16718 10110 16770
rect 10162 16718 10164 16770
rect 9996 16716 10164 16718
rect 9548 16210 9604 16716
rect 10108 16706 10164 16716
rect 10332 16770 10388 18172
rect 10332 16718 10334 16770
rect 10386 16718 10388 16770
rect 10332 16706 10388 16718
rect 10444 16660 10500 16670
rect 10444 16566 10500 16604
rect 9948 16492 10212 16502
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 9948 16426 10212 16436
rect 9548 16158 9550 16210
rect 9602 16158 9604 16210
rect 8764 16100 8820 16110
rect 8764 16006 8820 16044
rect 8428 15374 8430 15426
rect 8482 15374 8484 15426
rect 8428 15362 8484 15374
rect 7644 15262 7646 15314
rect 7698 15262 7700 15314
rect 7644 15250 7700 15262
rect 9548 15314 9604 16158
rect 9548 15262 9550 15314
rect 9602 15262 9604 15314
rect 9548 15148 9604 15262
rect 10332 15202 10388 15214
rect 10332 15150 10334 15202
rect 10386 15150 10388 15202
rect 7756 15092 7812 15102
rect 9548 15092 9716 15148
rect 7756 14530 7812 15036
rect 9660 15026 9716 15036
rect 9948 14924 10212 14934
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 9948 14858 10212 14868
rect 10332 14756 10388 15150
rect 9884 14700 10388 14756
rect 7756 14478 7758 14530
rect 7810 14478 7812 14530
rect 7756 14466 7812 14478
rect 8428 14532 8484 14542
rect 8428 14438 8484 14476
rect 8652 14308 8708 14318
rect 7756 13860 7812 13870
rect 7532 13858 7812 13860
rect 7532 13806 7758 13858
rect 7810 13806 7812 13858
rect 7532 13804 7812 13806
rect 7756 13794 7812 13804
rect 7980 13636 8036 13646
rect 7980 13542 8036 13580
rect 8316 13636 8372 13646
rect 8316 13542 8372 13580
rect 8652 13074 8708 14252
rect 9884 13970 9940 14700
rect 10556 14642 10612 19068
rect 10780 18450 10836 18462
rect 10780 18398 10782 18450
rect 10834 18398 10836 18450
rect 10780 17892 10836 18398
rect 10780 17826 10836 17836
rect 10892 17778 10948 19068
rect 11452 19124 11508 20076
rect 11452 19058 11508 19068
rect 11564 20018 11620 20030
rect 11564 19966 11566 20018
rect 11618 19966 11620 20018
rect 11228 19012 11284 19022
rect 11228 19010 11396 19012
rect 11228 18958 11230 19010
rect 11282 18958 11396 19010
rect 11228 18956 11396 18958
rect 11228 18946 11284 18956
rect 11116 18676 11172 18686
rect 11116 18582 11172 18620
rect 11340 18674 11396 18956
rect 11340 18622 11342 18674
rect 11394 18622 11396 18674
rect 11340 18610 11396 18622
rect 11564 18562 11620 19966
rect 11788 19684 11844 19694
rect 11788 19458 11844 19628
rect 11788 19406 11790 19458
rect 11842 19406 11844 19458
rect 11788 19394 11844 19406
rect 11900 19460 11956 19470
rect 11900 19366 11956 19404
rect 11900 19234 11956 19246
rect 11900 19182 11902 19234
rect 11954 19182 11956 19234
rect 11900 19124 11956 19182
rect 11900 19058 11956 19068
rect 11564 18510 11566 18562
rect 11618 18510 11620 18562
rect 11564 18498 11620 18510
rect 12012 18676 12068 22092
rect 13132 22082 13188 22092
rect 18508 22146 18788 22148
rect 18508 22094 18734 22146
rect 18786 22094 18788 22146
rect 18508 22092 18788 22094
rect 12860 21980 13124 21990
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 18508 21924 18564 22092
rect 18732 22082 18788 22092
rect 19180 22148 19236 22158
rect 19180 22054 19236 22092
rect 20188 22146 20244 22158
rect 20188 22094 20190 22146
rect 20242 22094 20244 22146
rect 12860 21914 13124 21924
rect 18396 21868 18564 21924
rect 18684 21980 18948 21990
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18684 21914 18948 21924
rect 15484 21756 15876 21812
rect 13020 21588 13076 21598
rect 13020 21494 13076 21532
rect 12572 21476 12628 21486
rect 13692 21476 13748 21486
rect 12572 21474 12740 21476
rect 12572 21422 12574 21474
rect 12626 21422 12740 21474
rect 12572 21420 12740 21422
rect 12572 21410 12628 21420
rect 12684 20132 12740 21420
rect 13692 21474 13972 21476
rect 13692 21422 13694 21474
rect 13746 21422 13972 21474
rect 13692 21420 13972 21422
rect 13692 21410 13748 21420
rect 12860 20412 13124 20422
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 12860 20346 13124 20356
rect 13916 20242 13972 21420
rect 13916 20190 13918 20242
rect 13970 20190 13972 20242
rect 13916 20178 13972 20190
rect 12908 20132 12964 20142
rect 13244 20132 13300 20142
rect 12684 20130 12964 20132
rect 12684 20078 12910 20130
rect 12962 20078 12964 20130
rect 12684 20076 12964 20078
rect 12908 19796 12964 20076
rect 13132 20076 13244 20132
rect 13132 20018 13188 20076
rect 13244 20066 13300 20076
rect 14140 20132 14196 20142
rect 14140 20038 14196 20076
rect 14924 20132 14980 20142
rect 14924 20038 14980 20076
rect 15148 20132 15204 20142
rect 13132 19966 13134 20018
rect 13186 19966 13188 20018
rect 13132 19954 13188 19966
rect 13580 20020 13636 20030
rect 13804 20020 13860 20030
rect 13580 20018 13972 20020
rect 13580 19966 13582 20018
rect 13634 19966 13806 20018
rect 13858 19966 13972 20018
rect 13580 19964 13972 19966
rect 13580 19954 13636 19964
rect 13804 19954 13860 19964
rect 13356 19908 13412 19918
rect 12908 19730 12964 19740
rect 13244 19906 13412 19908
rect 13244 19854 13358 19906
rect 13410 19854 13412 19906
rect 13244 19852 13412 19854
rect 13916 19908 13972 19964
rect 14252 20018 14308 20030
rect 14252 19966 14254 20018
rect 14306 19966 14308 20018
rect 13916 19852 14084 19908
rect 13244 19572 13300 19852
rect 13356 19842 13412 19852
rect 12572 19516 13300 19572
rect 13804 19796 13860 19806
rect 12572 19458 12628 19516
rect 12572 19406 12574 19458
rect 12626 19406 12628 19458
rect 12572 19394 12628 19406
rect 13804 19346 13860 19740
rect 13804 19294 13806 19346
rect 13858 19294 13860 19346
rect 13804 19282 13860 19294
rect 12348 19234 12404 19246
rect 12348 19182 12350 19234
rect 12402 19182 12404 19234
rect 12348 19012 12404 19182
rect 12348 18946 12404 18956
rect 13916 19236 13972 19246
rect 12860 18844 13124 18854
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 12860 18778 13124 18788
rect 12012 18450 12068 18620
rect 12012 18398 12014 18450
rect 12066 18398 12068 18450
rect 10892 17726 10894 17778
rect 10946 17726 10948 17778
rect 10892 17714 10948 17726
rect 11004 18226 11060 18238
rect 11004 18174 11006 18226
rect 11058 18174 11060 18226
rect 11004 17108 11060 18174
rect 11340 17892 11396 17902
rect 11340 17666 11396 17836
rect 12012 17778 12068 18398
rect 12236 18562 12292 18574
rect 12236 18510 12238 18562
rect 12290 18510 12292 18562
rect 12236 18452 12292 18510
rect 12236 18386 12292 18396
rect 12572 18562 12628 18574
rect 12572 18510 12574 18562
rect 12626 18510 12628 18562
rect 12572 18340 12628 18510
rect 12572 18274 12628 18284
rect 12908 18452 12964 18462
rect 12012 17726 12014 17778
rect 12066 17726 12068 17778
rect 12012 17714 12068 17726
rect 11340 17614 11342 17666
rect 11394 17614 11396 17666
rect 11340 17602 11396 17614
rect 12908 17556 12964 18396
rect 12908 17490 12964 17500
rect 11004 17042 11060 17052
rect 11900 17442 11956 17454
rect 11900 17390 11902 17442
rect 11954 17390 11956 17442
rect 11004 16882 11060 16894
rect 11004 16830 11006 16882
rect 11058 16830 11060 16882
rect 11004 16772 11060 16830
rect 11004 16706 11060 16716
rect 11788 16772 11844 16782
rect 11788 16678 11844 16716
rect 11900 16660 11956 17390
rect 13916 17332 13972 19180
rect 14028 18564 14084 19852
rect 14252 18674 14308 19966
rect 15148 19460 15204 20076
rect 15260 20018 15316 20030
rect 15260 19966 15262 20018
rect 15314 19966 15316 20018
rect 15260 19572 15316 19966
rect 15484 19572 15540 21756
rect 15708 21588 15764 21598
rect 15596 21532 15708 21588
rect 15596 20802 15652 21532
rect 15708 21522 15764 21532
rect 15820 21474 15876 21756
rect 17500 21700 17556 21710
rect 17500 21606 17556 21644
rect 16268 21588 16324 21598
rect 17388 21588 17444 21598
rect 16268 21494 16324 21532
rect 17164 21586 17444 21588
rect 17164 21534 17390 21586
rect 17442 21534 17444 21586
rect 17164 21532 17444 21534
rect 15820 21422 15822 21474
rect 15874 21422 15876 21474
rect 15820 21410 15876 21422
rect 16492 21364 16548 21374
rect 15772 21196 16036 21206
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 15772 21130 16036 21140
rect 15596 20750 15598 20802
rect 15650 20750 15652 20802
rect 15596 20738 15652 20750
rect 16380 20690 16436 20702
rect 16380 20638 16382 20690
rect 16434 20638 16436 20690
rect 16044 20018 16100 20030
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 16044 19796 16100 19966
rect 16380 19908 16436 20638
rect 16492 20130 16548 21308
rect 16492 20078 16494 20130
rect 16546 20078 16548 20130
rect 16492 20066 16548 20078
rect 16604 20132 16660 20142
rect 16604 20038 16660 20076
rect 16828 20020 16884 20030
rect 17164 20020 17220 21532
rect 17388 21522 17444 21532
rect 17948 21588 18004 21598
rect 17500 21364 17556 21374
rect 17500 21270 17556 21308
rect 16828 20018 17220 20020
rect 16828 19966 16830 20018
rect 16882 19966 17220 20018
rect 16828 19964 17220 19966
rect 17276 20132 17332 20142
rect 16492 19908 16548 19918
rect 16380 19906 16548 19908
rect 16380 19854 16494 19906
rect 16546 19854 16548 19906
rect 16380 19852 16548 19854
rect 16492 19842 16548 19852
rect 16716 19796 16772 19806
rect 16100 19740 16324 19796
rect 16044 19730 16100 19740
rect 15772 19628 16036 19638
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 15260 19516 15652 19572
rect 15772 19562 16036 19572
rect 15148 19404 15540 19460
rect 14364 19236 14420 19246
rect 14364 19142 14420 19180
rect 14588 19236 14644 19246
rect 14588 19142 14644 19180
rect 14812 19234 14868 19246
rect 14812 19182 14814 19234
rect 14866 19182 14868 19234
rect 14476 19012 14532 19022
rect 14476 18918 14532 18956
rect 14812 19012 14868 19182
rect 14812 18946 14868 18956
rect 14924 19234 14980 19246
rect 14924 19182 14926 19234
rect 14978 19182 14980 19234
rect 14252 18622 14254 18674
rect 14306 18622 14308 18674
rect 14252 18610 14308 18622
rect 14364 18676 14420 18686
rect 14364 18582 14420 18620
rect 14140 18564 14196 18574
rect 14028 18562 14196 18564
rect 14028 18510 14142 18562
rect 14194 18510 14196 18562
rect 14028 18508 14196 18510
rect 14140 18452 14196 18508
rect 14140 18386 14196 18396
rect 14812 18450 14868 18462
rect 14812 18398 14814 18450
rect 14866 18398 14868 18450
rect 14812 18340 14868 18398
rect 14812 18274 14868 18284
rect 14924 18228 14980 19182
rect 15148 18676 15204 19404
rect 15484 19346 15540 19404
rect 15484 19294 15486 19346
rect 15538 19294 15540 19346
rect 15484 19282 15540 19294
rect 15372 19236 15428 19246
rect 15372 19142 15428 19180
rect 15260 19012 15316 19022
rect 15316 18956 15428 19012
rect 15260 18946 15316 18956
rect 15148 18610 15204 18620
rect 15260 18562 15316 18574
rect 15260 18510 15262 18562
rect 15314 18510 15316 18562
rect 15148 18452 15204 18462
rect 15148 18358 15204 18396
rect 15260 18340 15316 18510
rect 15260 18274 15316 18284
rect 15036 18228 15092 18238
rect 14924 18226 15092 18228
rect 14924 18174 15038 18226
rect 15090 18174 15092 18226
rect 14924 18172 15092 18174
rect 14364 17892 14420 17902
rect 14924 17892 14980 18172
rect 15036 18162 15092 18172
rect 15372 18004 15428 18956
rect 14364 17890 14980 17892
rect 14364 17838 14366 17890
rect 14418 17838 14980 17890
rect 14364 17836 14980 17838
rect 15036 17948 15428 18004
rect 15484 18452 15540 18462
rect 14364 17826 14420 17836
rect 14476 17556 14532 17566
rect 14476 17554 14868 17556
rect 14476 17502 14478 17554
rect 14530 17502 14868 17554
rect 14476 17500 14868 17502
rect 14476 17490 14532 17500
rect 14364 17444 14420 17454
rect 12860 17276 13124 17286
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 13916 17266 13972 17276
rect 14252 17442 14420 17444
rect 14252 17390 14366 17442
rect 14418 17390 14420 17442
rect 14252 17388 14420 17390
rect 12860 17210 13124 17220
rect 14252 16996 14308 17388
rect 14364 17378 14420 17388
rect 13916 16994 14308 16996
rect 13916 16942 14254 16994
rect 14306 16942 14308 16994
rect 13916 16940 14308 16942
rect 13580 16772 13636 16782
rect 11900 15204 11956 16604
rect 13468 16660 13524 16670
rect 13468 15988 13524 16604
rect 13580 16322 13636 16716
rect 13916 16770 13972 16940
rect 14252 16930 14308 16940
rect 14364 16996 14420 17006
rect 14364 16994 14756 16996
rect 14364 16942 14366 16994
rect 14418 16942 14756 16994
rect 14364 16940 14756 16942
rect 14364 16930 14420 16940
rect 13916 16718 13918 16770
rect 13970 16718 13972 16770
rect 13916 16706 13972 16718
rect 13580 16270 13582 16322
rect 13634 16270 13636 16322
rect 13580 16258 13636 16270
rect 14476 16324 14532 16334
rect 13580 15988 13636 15998
rect 13468 15986 13636 15988
rect 13468 15934 13582 15986
rect 13634 15934 13636 15986
rect 13468 15932 13636 15934
rect 13580 15922 13636 15932
rect 13692 15988 13748 15998
rect 14140 15988 14196 15998
rect 13692 15986 14196 15988
rect 13692 15934 13694 15986
rect 13746 15934 14142 15986
rect 14194 15934 14196 15986
rect 13692 15932 14196 15934
rect 13692 15922 13748 15932
rect 14140 15922 14196 15932
rect 12860 15708 13124 15718
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 12860 15642 13124 15652
rect 14252 15540 14308 15550
rect 14140 15538 14308 15540
rect 14140 15486 14254 15538
rect 14306 15486 14308 15538
rect 14140 15484 14308 15486
rect 12236 15260 12516 15316
rect 12236 15148 12292 15260
rect 11900 15138 11956 15148
rect 10556 14590 10558 14642
rect 10610 14590 10612 14642
rect 10556 14578 10612 14590
rect 12124 15092 12292 15148
rect 12460 15202 12516 15260
rect 12460 15150 12462 15202
rect 12514 15150 12516 15202
rect 12460 15138 12516 15150
rect 12348 15092 12404 15102
rect 9884 13918 9886 13970
rect 9938 13918 9940 13970
rect 9884 13906 9940 13918
rect 9548 13746 9604 13758
rect 9548 13694 9550 13746
rect 9602 13694 9604 13746
rect 9548 13636 9604 13694
rect 11228 13748 11284 13758
rect 11564 13748 11620 13758
rect 11284 13746 11620 13748
rect 11284 13694 11566 13746
rect 11618 13694 11620 13746
rect 11284 13692 11620 13694
rect 11228 13654 11284 13692
rect 11564 13682 11620 13692
rect 9548 13570 9604 13580
rect 9948 13356 10212 13366
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 9948 13290 10212 13300
rect 8652 13022 8654 13074
rect 8706 13022 8708 13074
rect 8652 13010 8708 13022
rect 10780 13074 10836 13086
rect 10780 13022 10782 13074
rect 10834 13022 10836 13074
rect 7868 12964 7924 12974
rect 7868 11284 7924 12908
rect 10332 12290 10388 12302
rect 10332 12238 10334 12290
rect 10386 12238 10388 12290
rect 7868 11218 7924 11228
rect 8764 12066 8820 12078
rect 8764 12014 8766 12066
rect 8818 12014 8820 12066
rect 8764 10612 8820 12014
rect 9948 11788 10212 11798
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 9948 11722 10212 11732
rect 8764 10546 8820 10556
rect 9324 11284 9380 11294
rect 7420 9314 7476 9324
rect 7644 10498 7700 10510
rect 7644 10446 7646 10498
rect 7698 10446 7700 10498
rect 7196 9268 7252 9278
rect 7084 9212 7196 9268
rect 7084 9042 7140 9212
rect 7196 9202 7252 9212
rect 7308 9266 7364 9278
rect 7308 9214 7310 9266
rect 7362 9214 7364 9266
rect 7308 9156 7364 9214
rect 7308 9100 7588 9156
rect 7084 8990 7086 9042
rect 7138 8990 7140 9042
rect 7084 8978 7140 8990
rect 7532 8370 7588 9100
rect 7532 8318 7534 8370
rect 7586 8318 7588 8370
rect 7532 8306 7588 8318
rect 6860 8206 6862 8258
rect 6914 8206 6916 8258
rect 6636 7588 6692 7598
rect 6636 7494 6692 7532
rect 6412 7422 6414 7474
rect 6466 7422 6468 7474
rect 6412 7410 6468 7422
rect 5852 7198 5854 7250
rect 5906 7198 5908 7250
rect 4732 6638 4734 6690
rect 4786 6638 4788 6690
rect 4732 6626 4788 6638
rect 4396 6468 4452 6478
rect 4060 6466 4452 6468
rect 4060 6414 4398 6466
rect 4450 6414 4452 6466
rect 4060 6412 4452 6414
rect 4060 6018 4116 6412
rect 4396 6402 4452 6412
rect 4060 5966 4062 6018
rect 4114 5966 4116 6018
rect 4060 5954 4116 5966
rect 3388 5854 3390 5906
rect 3442 5854 3444 5906
rect 3388 5842 3444 5854
rect 5852 5796 5908 7198
rect 6188 5796 6244 5806
rect 5852 5794 6244 5796
rect 5852 5742 6190 5794
rect 6242 5742 6244 5794
rect 5852 5740 6244 5742
rect 6188 5730 6244 5740
rect 4124 5516 4388 5526
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4124 5450 4388 5460
rect 6860 5124 6916 8206
rect 7036 7868 7300 7878
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7036 7802 7300 7812
rect 7196 7588 7252 7598
rect 7196 7494 7252 7532
rect 7532 7476 7588 7486
rect 7644 7476 7700 10446
rect 8540 9828 8596 9838
rect 9212 9828 9268 9838
rect 9324 9828 9380 11228
rect 9772 10724 9828 10734
rect 9772 10630 9828 10668
rect 10220 10724 10276 10734
rect 10220 10630 10276 10668
rect 9948 10220 10212 10230
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 9948 10154 10212 10164
rect 10332 10052 10388 12238
rect 10668 12292 10724 12302
rect 10668 10724 10724 12236
rect 10780 12180 10836 13022
rect 10892 12180 10948 12190
rect 10780 12178 10948 12180
rect 10780 12126 10894 12178
rect 10946 12126 10948 12178
rect 10780 12124 10948 12126
rect 10892 12114 10948 12124
rect 11676 12180 11732 12190
rect 11676 12086 11732 12124
rect 12124 12068 12180 15092
rect 11788 12012 12180 12068
rect 12348 14306 12404 15036
rect 12908 14644 12964 14654
rect 12348 14254 12350 14306
rect 12402 14254 12404 14306
rect 12348 12068 12404 14254
rect 12684 14588 12908 14644
rect 12460 13748 12516 13758
rect 12460 12290 12516 13692
rect 12460 12238 12462 12290
rect 12514 12238 12516 12290
rect 12460 12226 12516 12238
rect 12684 12292 12740 14588
rect 12908 14550 12964 14588
rect 12860 14140 13124 14150
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 12860 14074 13124 14084
rect 14140 13748 14196 15484
rect 14252 15474 14308 15484
rect 14476 15428 14532 16268
rect 14588 16098 14644 16940
rect 14700 16882 14756 16940
rect 14700 16830 14702 16882
rect 14754 16830 14756 16882
rect 14700 16818 14756 16830
rect 14812 16994 14868 17500
rect 14812 16942 14814 16994
rect 14866 16942 14868 16994
rect 14812 16324 14868 16942
rect 15036 16436 15092 17948
rect 15484 16660 15540 18396
rect 15596 17892 15652 19516
rect 16268 18452 16324 19740
rect 16492 19684 16548 19694
rect 16268 18386 16324 18396
rect 16380 19010 16436 19022
rect 16380 18958 16382 19010
rect 16434 18958 16436 19010
rect 16156 18340 16212 18350
rect 15772 18060 16036 18070
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 15772 17994 16036 18004
rect 16156 17892 16212 18284
rect 16380 18228 16436 18958
rect 16380 18162 16436 18172
rect 15596 17836 15764 17892
rect 15708 16882 15764 17836
rect 15932 17836 16212 17892
rect 16492 17890 16548 19628
rect 16716 19458 16772 19740
rect 16828 19684 16884 19964
rect 16828 19618 16884 19628
rect 16716 19406 16718 19458
rect 16770 19406 16772 19458
rect 16716 19394 16772 19406
rect 16940 19236 16996 19246
rect 16940 19142 16996 19180
rect 17276 19234 17332 20076
rect 17948 20132 18004 21532
rect 18396 21588 18452 21868
rect 18396 21522 18452 21532
rect 18508 21700 18564 21710
rect 18508 20914 18564 21644
rect 20188 21588 20244 22094
rect 20860 22148 20916 22318
rect 21420 22370 21476 22382
rect 21420 22318 21422 22370
rect 21474 22318 21476 22370
rect 20860 22082 20916 22092
rect 21084 22146 21140 22158
rect 21084 22094 21086 22146
rect 21138 22094 21140 22146
rect 21084 21924 21140 22094
rect 21084 21858 21140 21868
rect 21420 21700 21476 22318
rect 24508 21980 24772 21990
rect 21420 21634 21476 21644
rect 23660 21924 23716 21934
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24508 21914 24772 21924
rect 20188 21522 20244 21532
rect 21196 21586 21252 21598
rect 21196 21534 21198 21586
rect 21250 21534 21252 21586
rect 18732 21476 18788 21486
rect 18732 21382 18788 21420
rect 20412 21476 20468 21486
rect 18508 20862 18510 20914
rect 18562 20862 18564 20914
rect 18508 20850 18564 20862
rect 19628 20914 19684 20926
rect 19628 20862 19630 20914
rect 19682 20862 19684 20914
rect 19516 20804 19572 20814
rect 19516 20710 19572 20748
rect 18684 20412 18948 20422
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18684 20346 18948 20356
rect 17948 20066 18004 20076
rect 18732 20132 18788 20142
rect 18732 20038 18788 20076
rect 19404 20132 19460 20142
rect 19404 20038 19460 20076
rect 18172 20018 18228 20030
rect 18172 19966 18174 20018
rect 18226 19966 18228 20018
rect 17948 19906 18004 19918
rect 17948 19854 17950 19906
rect 18002 19854 18004 19906
rect 17836 19796 17892 19806
rect 17836 19702 17892 19740
rect 17948 19346 18004 19854
rect 18172 19460 18228 19966
rect 18172 19394 18228 19404
rect 19628 20018 19684 20862
rect 20412 20914 20468 21420
rect 20412 20862 20414 20914
rect 20466 20862 20468 20914
rect 20412 20850 20468 20862
rect 20860 21474 20916 21486
rect 20860 21422 20862 21474
rect 20914 21422 20916 21474
rect 20860 20804 20916 21422
rect 19964 20692 20020 20702
rect 20300 20692 20356 20702
rect 19964 20690 20356 20692
rect 19964 20638 19966 20690
rect 20018 20638 20302 20690
rect 20354 20638 20356 20690
rect 19964 20636 20356 20638
rect 19964 20626 20020 20636
rect 20300 20626 20356 20636
rect 20636 20692 20692 20702
rect 20412 20580 20468 20590
rect 20412 20468 20468 20524
rect 20300 20412 20468 20468
rect 20524 20578 20580 20590
rect 20524 20526 20526 20578
rect 20578 20526 20580 20578
rect 19628 19966 19630 20018
rect 19682 19966 19684 20018
rect 17948 19294 17950 19346
rect 18002 19294 18004 19346
rect 17948 19282 18004 19294
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 17276 19170 17332 19182
rect 19628 19236 19684 19966
rect 19852 20130 19908 20142
rect 19852 20078 19854 20130
rect 19906 20078 19908 20130
rect 19852 19348 19908 20078
rect 19852 19282 19908 19292
rect 19964 20018 20020 20030
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19964 19796 20020 19966
rect 20300 19906 20356 20412
rect 20524 20356 20580 20526
rect 20300 19854 20302 19906
rect 20354 19854 20356 19906
rect 20300 19842 20356 19854
rect 20412 20300 20580 20356
rect 20412 20130 20468 20300
rect 20412 20078 20414 20130
rect 20466 20078 20468 20130
rect 19628 19170 19684 19180
rect 16604 19012 16660 19022
rect 16604 18918 16660 18956
rect 18684 18844 18948 18854
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18684 18778 18948 18788
rect 17388 18562 17444 18574
rect 17388 18510 17390 18562
rect 17442 18510 17444 18562
rect 17388 18452 17444 18510
rect 17388 18386 17444 18396
rect 17612 18450 17668 18462
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 16492 17838 16494 17890
rect 16546 17838 16548 17890
rect 15932 17778 15988 17836
rect 15932 17726 15934 17778
rect 15986 17726 15988 17778
rect 15932 17714 15988 17726
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16818 15764 16830
rect 16044 16660 16100 17836
rect 16492 17826 16548 17838
rect 16828 18340 16884 18350
rect 16156 17668 16212 17678
rect 16156 17666 16772 17668
rect 16156 17614 16158 17666
rect 16210 17614 16772 17666
rect 16156 17612 16772 17614
rect 16156 17602 16212 17612
rect 16268 17332 16324 17342
rect 16156 17106 16212 17118
rect 16156 17054 16158 17106
rect 16210 17054 16212 17106
rect 16156 16996 16212 17054
rect 16156 16930 16212 16940
rect 16268 16994 16324 17276
rect 16268 16942 16270 16994
rect 16322 16942 16324 16994
rect 16268 16930 16324 16942
rect 16492 16996 16548 17006
rect 16044 16604 16212 16660
rect 15036 16380 15204 16436
rect 14812 16258 14868 16268
rect 14588 16046 14590 16098
rect 14642 16046 14644 16098
rect 14588 16034 14644 16046
rect 14924 16100 14980 16110
rect 14700 15988 14756 15998
rect 14700 15764 14756 15932
rect 14364 15314 14420 15326
rect 14364 15262 14366 15314
rect 14418 15262 14420 15314
rect 14364 15204 14420 15262
rect 14364 15138 14420 15148
rect 14476 14420 14532 15372
rect 14588 15708 14756 15764
rect 14588 15314 14644 15708
rect 14924 15652 14980 16044
rect 15036 16098 15092 16110
rect 15036 16046 15038 16098
rect 15090 16046 15092 16098
rect 15036 15988 15092 16046
rect 15036 15922 15092 15932
rect 14588 15262 14590 15314
rect 14642 15262 14644 15314
rect 14588 15250 14644 15262
rect 14700 15314 14756 15326
rect 14700 15262 14702 15314
rect 14754 15262 14756 15314
rect 14588 14756 14644 14766
rect 14700 14756 14756 15262
rect 14588 14754 14756 14756
rect 14588 14702 14590 14754
rect 14642 14702 14756 14754
rect 14588 14700 14756 14702
rect 14588 14690 14644 14700
rect 14476 14418 14644 14420
rect 14476 14366 14478 14418
rect 14530 14366 14644 14418
rect 14476 14364 14644 14366
rect 14476 14354 14532 14364
rect 14140 13682 14196 13692
rect 14252 13074 14308 13086
rect 14252 13022 14254 13074
rect 14306 13022 14308 13074
rect 12860 12572 13124 12582
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 12860 12506 13124 12516
rect 14252 12404 14308 13022
rect 14252 12338 14308 12348
rect 12684 12226 12740 12236
rect 14252 12068 14308 12078
rect 12348 12012 12516 12068
rect 11228 11954 11284 11966
rect 11228 11902 11230 11954
rect 11282 11902 11284 11954
rect 11228 11620 11284 11902
rect 11228 11554 11284 11564
rect 11452 11396 11508 11406
rect 11452 11302 11508 11340
rect 10668 10658 10724 10668
rect 11340 11284 11396 11294
rect 10444 10612 10500 10622
rect 10444 10518 10500 10556
rect 11340 10610 11396 11228
rect 11340 10558 11342 10610
rect 11394 10558 11396 10610
rect 11340 10546 11396 10558
rect 8540 9826 8708 9828
rect 8540 9774 8542 9826
rect 8594 9774 8708 9826
rect 8540 9772 8708 9774
rect 8540 9762 8596 9772
rect 8652 9380 8708 9772
rect 9212 9826 9380 9828
rect 9212 9774 9214 9826
rect 9266 9774 9380 9826
rect 9212 9772 9380 9774
rect 9996 9996 10332 10052
rect 9212 9762 9268 9772
rect 9884 9714 9940 9726
rect 9884 9662 9886 9714
rect 9938 9662 9940 9714
rect 8764 9604 8820 9614
rect 9884 9604 9940 9662
rect 8764 9602 9940 9604
rect 8764 9550 8766 9602
rect 8818 9550 9940 9602
rect 8764 9548 9940 9550
rect 8764 9538 8820 9548
rect 8652 9324 9716 9380
rect 9660 9266 9716 9324
rect 9660 9214 9662 9266
rect 9714 9214 9716 9266
rect 9660 9202 9716 9214
rect 9996 9042 10052 9996
rect 10332 9958 10388 9996
rect 10780 10386 10836 10398
rect 10780 10334 10782 10386
rect 10834 10334 10836 10386
rect 9996 8990 9998 9042
rect 10050 8990 10052 9042
rect 9996 8978 10052 8990
rect 10332 9154 10388 9166
rect 10332 9102 10334 9154
rect 10386 9102 10388 9154
rect 9948 8652 10212 8662
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 9948 8586 10212 8596
rect 9660 8370 9716 8382
rect 9660 8318 9662 8370
rect 9714 8318 9716 8370
rect 7532 7474 7700 7476
rect 7532 7422 7534 7474
rect 7586 7422 7700 7474
rect 7532 7420 7700 7422
rect 7756 7586 7812 7598
rect 7756 7534 7758 7586
rect 7810 7534 7812 7586
rect 7756 7476 7812 7534
rect 8316 7588 8372 7598
rect 8316 7494 8372 7532
rect 9212 7588 9268 7598
rect 7532 7410 7588 7420
rect 7756 7410 7812 7420
rect 9212 6916 9268 7532
rect 9660 7476 9716 8318
rect 10108 8372 10164 8382
rect 10332 8372 10388 9102
rect 10780 9154 10836 10334
rect 10780 9102 10782 9154
rect 10834 9102 10836 9154
rect 10780 9090 10836 9102
rect 11340 8930 11396 8942
rect 11340 8878 11342 8930
rect 11394 8878 11396 8930
rect 11340 8428 11396 8878
rect 10108 8370 10332 8372
rect 10108 8318 10110 8370
rect 10162 8318 10332 8370
rect 10108 8316 10332 8318
rect 10108 8306 10164 8316
rect 10332 8306 10388 8316
rect 10892 8372 11396 8428
rect 10444 8258 10500 8270
rect 10444 8206 10446 8258
rect 10498 8206 10500 8258
rect 10444 7812 10500 8206
rect 9660 7410 9716 7420
rect 10332 7476 10388 7486
rect 10332 7382 10388 7420
rect 9996 7252 10052 7262
rect 9772 7250 10052 7252
rect 9772 7198 9998 7250
rect 10050 7198 10052 7250
rect 9772 7196 10052 7198
rect 9212 6914 9716 6916
rect 9212 6862 9214 6914
rect 9266 6862 9716 6914
rect 9212 6860 9716 6862
rect 9212 6850 9268 6860
rect 8316 6692 8372 6702
rect 8316 6598 8372 6636
rect 8876 6692 8932 6702
rect 8876 6598 8932 6636
rect 7980 6468 8036 6478
rect 7756 6466 8036 6468
rect 7756 6414 7982 6466
rect 8034 6414 8036 6466
rect 7756 6412 8036 6414
rect 7036 6300 7300 6310
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7036 6234 7300 6244
rect 7756 5234 7812 6412
rect 7980 6402 8036 6412
rect 7756 5182 7758 5234
rect 7810 5182 7812 5234
rect 7756 5170 7812 5182
rect 9660 5236 9716 6860
rect 9772 6578 9828 7196
rect 9996 7186 10052 7196
rect 9948 7084 10212 7094
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 9948 7018 10212 7028
rect 10444 6804 10500 7756
rect 10556 7700 10612 7710
rect 10892 7700 10948 8372
rect 11788 8370 11844 12012
rect 12348 11172 12404 11182
rect 12124 11170 12404 11172
rect 12124 11118 12350 11170
rect 12402 11118 12404 11170
rect 12124 11116 12404 11118
rect 12124 10722 12180 11116
rect 12348 11106 12404 11116
rect 12124 10670 12126 10722
rect 12178 10670 12180 10722
rect 12124 10658 12180 10670
rect 12012 10052 12068 10062
rect 12012 9938 12068 9996
rect 12012 9886 12014 9938
rect 12066 9886 12068 9938
rect 12012 9874 12068 9886
rect 11788 8318 11790 8370
rect 11842 8318 11844 8370
rect 11788 8306 11844 8318
rect 11900 9044 11956 9054
rect 12460 9044 12516 12012
rect 13916 12012 14252 12068
rect 13916 11618 13972 12012
rect 13916 11566 13918 11618
rect 13970 11566 13972 11618
rect 13916 11554 13972 11566
rect 12684 11284 12740 11294
rect 12684 11190 12740 11228
rect 13580 11284 13636 11294
rect 13580 11190 13636 11228
rect 12860 11004 13124 11014
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 12860 10938 13124 10948
rect 14252 10498 14308 12012
rect 14588 12066 14644 14364
rect 14924 13858 14980 15596
rect 15148 15540 15204 16380
rect 15484 16212 15540 16604
rect 15772 16492 16036 16502
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 15772 16426 16036 16436
rect 16156 16324 16212 16604
rect 15820 16268 16212 16324
rect 15484 16156 15764 16212
rect 15484 15986 15540 15998
rect 15484 15934 15486 15986
rect 15538 15934 15540 15986
rect 15484 15652 15540 15934
rect 15596 15988 15652 15998
rect 15596 15894 15652 15932
rect 15708 15876 15764 16156
rect 15820 16098 15876 16268
rect 15820 16046 15822 16098
rect 15874 16046 15876 16098
rect 15820 16034 15876 16046
rect 15708 15820 15988 15876
rect 15484 15596 15652 15652
rect 15036 15428 15092 15438
rect 15148 15428 15204 15484
rect 15596 15538 15652 15596
rect 15596 15486 15598 15538
rect 15650 15486 15652 15538
rect 15596 15474 15652 15486
rect 15036 15426 15204 15428
rect 15036 15374 15038 15426
rect 15090 15374 15204 15426
rect 15036 15372 15204 15374
rect 15484 15428 15540 15438
rect 15036 15362 15092 15372
rect 15484 15334 15540 15372
rect 15596 15316 15652 15326
rect 15260 15204 15316 15214
rect 15260 15092 15428 15148
rect 15372 14642 15428 15092
rect 15596 14754 15652 15260
rect 15708 15314 15764 15326
rect 15708 15262 15710 15314
rect 15762 15262 15764 15314
rect 15708 15092 15764 15262
rect 15932 15148 15988 15820
rect 16044 15540 16100 16268
rect 16492 16098 16548 16940
rect 16492 16046 16494 16098
rect 16546 16046 16548 16098
rect 16492 16034 16548 16046
rect 16156 15876 16212 15886
rect 16156 15874 16436 15876
rect 16156 15822 16158 15874
rect 16210 15822 16436 15874
rect 16156 15820 16436 15822
rect 16156 15810 16212 15820
rect 16268 15540 16324 15550
rect 16044 15538 16324 15540
rect 16044 15486 16270 15538
rect 16322 15486 16324 15538
rect 16044 15484 16324 15486
rect 16268 15474 16324 15484
rect 15932 15092 16324 15148
rect 15708 15026 15764 15036
rect 15772 14924 16036 14934
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 15772 14858 16036 14868
rect 15596 14702 15598 14754
rect 15650 14702 15652 14754
rect 15596 14690 15652 14702
rect 15372 14590 15374 14642
rect 15426 14590 15428 14642
rect 15372 14578 15428 14590
rect 16268 14532 16324 15092
rect 16380 15092 16436 15820
rect 16604 15428 16660 15438
rect 16492 15316 16548 15354
rect 16492 15250 16548 15260
rect 16380 15026 16436 15036
rect 16492 14980 16548 14990
rect 16492 14644 16548 14924
rect 16380 14532 16436 14542
rect 16268 14530 16436 14532
rect 16268 14478 16382 14530
rect 16434 14478 16436 14530
rect 16268 14476 16436 14478
rect 16380 14466 16436 14476
rect 15932 14308 15988 14318
rect 15932 14306 16212 14308
rect 15932 14254 15934 14306
rect 15986 14254 16212 14306
rect 15932 14252 16212 14254
rect 15932 14242 15988 14252
rect 14924 13806 14926 13858
rect 14978 13806 14980 13858
rect 14588 12014 14590 12066
rect 14642 12014 14644 12066
rect 14588 12002 14644 12014
rect 14812 12180 14868 12190
rect 14700 11844 14756 11854
rect 14476 11620 14532 11630
rect 14476 11282 14532 11564
rect 14476 11230 14478 11282
rect 14530 11230 14532 11282
rect 14476 11218 14532 11230
rect 14700 11394 14756 11788
rect 14700 11342 14702 11394
rect 14754 11342 14756 11394
rect 14252 10446 14254 10498
rect 14306 10446 14308 10498
rect 14252 10434 14308 10446
rect 14700 9716 14756 11342
rect 14812 10836 14868 12124
rect 14924 11396 14980 13806
rect 15772 13356 16036 13366
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 15772 13290 16036 13300
rect 15484 12404 15540 12414
rect 15484 12310 15540 12348
rect 15596 12292 15652 12302
rect 15036 12178 15092 12190
rect 15036 12126 15038 12178
rect 15090 12126 15092 12178
rect 15036 12068 15092 12126
rect 15036 12002 15092 12012
rect 15260 12178 15316 12190
rect 15260 12126 15262 12178
rect 15314 12126 15316 12178
rect 14924 11330 14980 11340
rect 14924 10836 14980 10846
rect 14812 10834 14980 10836
rect 14812 10782 14926 10834
rect 14978 10782 14980 10834
rect 14812 10780 14980 10782
rect 14924 10770 14980 10780
rect 15260 10724 15316 12126
rect 15596 12178 15652 12236
rect 15596 12126 15598 12178
rect 15650 12126 15652 12178
rect 15372 12068 15428 12078
rect 15372 11974 15428 12012
rect 15596 11844 15652 12126
rect 16156 12178 16212 14252
rect 16492 14196 16548 14588
rect 16604 14530 16660 15372
rect 16716 15092 16772 17612
rect 16828 17666 16884 18284
rect 17612 18228 17668 18398
rect 19180 18452 19236 18462
rect 19180 18450 19348 18452
rect 19180 18398 19182 18450
rect 19234 18398 19348 18450
rect 19180 18396 19348 18398
rect 19180 18386 19236 18396
rect 17612 18162 17668 18172
rect 16828 17614 16830 17666
rect 16882 17614 16884 17666
rect 16828 17602 16884 17614
rect 17164 17668 17220 17678
rect 17164 17574 17220 17612
rect 18060 17668 18116 17678
rect 18060 17574 18116 17612
rect 19180 17668 19236 17678
rect 19180 17574 19236 17612
rect 16940 17556 16996 17566
rect 16940 17462 16996 17500
rect 18284 17442 18340 17454
rect 18284 17390 18286 17442
rect 18338 17390 18340 17442
rect 17388 16882 17444 16894
rect 17388 16830 17390 16882
rect 17442 16830 17444 16882
rect 16716 15026 16772 15036
rect 17276 16212 17332 16222
rect 17276 16098 17332 16156
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 14532 17332 16046
rect 17388 15652 17444 16830
rect 18060 15988 18116 15998
rect 18060 15894 18116 15932
rect 17388 15586 17444 15596
rect 17388 15428 17444 15438
rect 17388 15334 17444 15372
rect 17612 15316 17668 15326
rect 17612 15222 17668 15260
rect 18284 15148 18340 17390
rect 18684 17276 18948 17286
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18684 17210 18948 17220
rect 19292 16548 19348 18396
rect 19964 18450 20020 19740
rect 20412 19458 20468 20078
rect 20412 19406 20414 19458
rect 20466 19406 20468 19458
rect 20412 19394 20468 19406
rect 20524 20132 20580 20142
rect 20076 19348 20132 19358
rect 20076 19254 20132 19292
rect 20524 19348 20580 20076
rect 20636 20130 20692 20636
rect 20860 20244 20916 20748
rect 20860 20178 20916 20188
rect 20636 20078 20638 20130
rect 20690 20078 20692 20130
rect 20636 20066 20692 20078
rect 21196 20132 21252 21534
rect 23548 21588 23604 21598
rect 21980 21474 22036 21486
rect 21980 21422 21982 21474
rect 22034 21422 22036 21474
rect 21596 21196 21860 21206
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21596 21130 21860 21140
rect 21980 21028 22036 21422
rect 21868 20972 22036 21028
rect 21756 20692 21812 20702
rect 21756 20598 21812 20636
rect 21532 20578 21588 20590
rect 21532 20526 21534 20578
rect 21586 20526 21588 20578
rect 21196 20066 21252 20076
rect 21308 20130 21364 20142
rect 21308 20078 21310 20130
rect 21362 20078 21364 20130
rect 21084 20020 21140 20030
rect 21084 19926 21140 19964
rect 20860 19458 20916 19470
rect 20860 19406 20862 19458
rect 20914 19406 20916 19458
rect 20524 19346 20692 19348
rect 20524 19294 20526 19346
rect 20578 19294 20692 19346
rect 20524 19292 20692 19294
rect 20524 19282 20580 19292
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19292 16482 19348 16492
rect 19404 18338 19460 18350
rect 19404 18286 19406 18338
rect 19458 18286 19460 18338
rect 18684 15708 18948 15718
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18684 15642 18948 15652
rect 19404 15316 19460 18286
rect 19516 18228 19572 18238
rect 19964 18228 20020 18398
rect 20076 19012 20132 19022
rect 20076 18450 20132 18956
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 20076 18386 20132 18398
rect 20636 18452 20692 19292
rect 20412 18340 20468 18350
rect 20412 18246 20468 18284
rect 19516 18226 19684 18228
rect 19516 18174 19518 18226
rect 19570 18174 19684 18226
rect 19516 18172 19684 18174
rect 19964 18172 20244 18228
rect 19516 18162 19572 18172
rect 19516 17444 19572 17454
rect 19516 17350 19572 17388
rect 19628 16100 19684 18172
rect 20188 17890 20244 18172
rect 20188 17838 20190 17890
rect 20242 17838 20244 17890
rect 20188 17826 20244 17838
rect 20300 18226 20356 18238
rect 20300 18174 20302 18226
rect 20354 18174 20356 18226
rect 20300 17668 20356 18174
rect 20524 18228 20580 18238
rect 20524 17892 20580 18172
rect 20188 16548 20244 16558
rect 20188 16210 20244 16492
rect 20188 16158 20190 16210
rect 20242 16158 20244 16210
rect 20188 16146 20244 16158
rect 19628 16034 19684 16044
rect 20076 15988 20132 15998
rect 20076 15426 20132 15932
rect 20076 15374 20078 15426
rect 20130 15374 20132 15426
rect 20076 15362 20132 15374
rect 19404 15250 19460 15260
rect 20188 15316 20244 15326
rect 20300 15316 20356 17612
rect 20188 15314 20356 15316
rect 20188 15262 20190 15314
rect 20242 15262 20356 15314
rect 20188 15260 20356 15262
rect 20412 17890 20580 17892
rect 20412 17838 20526 17890
rect 20578 17838 20580 17890
rect 20412 17836 20580 17838
rect 20412 15314 20468 17836
rect 20524 17826 20580 17836
rect 20636 16994 20692 18396
rect 20748 18338 20804 18350
rect 20748 18286 20750 18338
rect 20802 18286 20804 18338
rect 20748 17780 20804 18286
rect 20748 17686 20804 17724
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16212 20692 16942
rect 20412 15262 20414 15314
rect 20466 15262 20468 15314
rect 20188 15250 20244 15260
rect 20412 15250 20468 15262
rect 20524 15316 20580 15326
rect 20524 15222 20580 15260
rect 18284 15092 18452 15148
rect 17500 14532 17556 14542
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16604 14466 16660 14478
rect 16940 14530 17556 14532
rect 16940 14478 17502 14530
rect 17554 14478 17556 14530
rect 16940 14476 17556 14478
rect 16156 12126 16158 12178
rect 16210 12126 16212 12178
rect 15596 11778 15652 11788
rect 15772 11788 16036 11798
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 15772 11722 16036 11732
rect 15484 11396 15540 11406
rect 15484 11302 15540 11340
rect 15932 10836 15988 10846
rect 16156 10836 16212 12126
rect 15932 10834 16212 10836
rect 15932 10782 15934 10834
rect 15986 10782 16212 10834
rect 15932 10780 16212 10782
rect 16268 14140 16548 14196
rect 16716 14418 16772 14430
rect 16716 14366 16718 14418
rect 16770 14366 16772 14418
rect 16268 10836 16324 14140
rect 16716 13076 16772 14366
rect 16716 13010 16772 13020
rect 16380 12852 16436 12862
rect 16380 12850 16772 12852
rect 16380 12798 16382 12850
rect 16434 12798 16772 12850
rect 16380 12796 16772 12798
rect 16380 12786 16436 12796
rect 16716 12402 16772 12796
rect 16716 12350 16718 12402
rect 16770 12350 16772 12402
rect 16716 12338 16772 12350
rect 16380 12292 16436 12302
rect 16380 12198 16436 12236
rect 16940 12180 16996 14476
rect 17500 14466 17556 14476
rect 18284 14418 18340 14430
rect 18284 14366 18286 14418
rect 18338 14366 18340 14418
rect 17164 14306 17220 14318
rect 17164 14254 17166 14306
rect 17218 14254 17220 14306
rect 17164 14196 17220 14254
rect 17164 14140 18004 14196
rect 17388 13972 17444 13982
rect 17388 13878 17444 13916
rect 17948 13858 18004 14140
rect 18284 13970 18340 14366
rect 18284 13918 18286 13970
rect 18338 13918 18340 13970
rect 18284 13906 18340 13918
rect 17948 13806 17950 13858
rect 18002 13806 18004 13858
rect 17948 13794 18004 13806
rect 17500 13634 17556 13646
rect 17500 13582 17502 13634
rect 17554 13582 17556 13634
rect 16940 12114 16996 12124
rect 17164 12962 17220 12974
rect 17164 12910 17166 12962
rect 17218 12910 17220 12962
rect 16828 12068 16884 12078
rect 16828 11974 16884 12012
rect 17164 11284 17220 12910
rect 17500 12404 17556 13582
rect 18284 13076 18340 13086
rect 18284 12982 18340 13020
rect 18396 12852 18452 15092
rect 20412 14644 20468 14654
rect 20300 14642 20468 14644
rect 20300 14590 20414 14642
rect 20466 14590 20468 14642
rect 20300 14588 20468 14590
rect 18684 14140 18948 14150
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18684 14074 18948 14084
rect 19628 13858 19684 13870
rect 19628 13806 19630 13858
rect 19682 13806 19684 13858
rect 18956 12964 19012 12974
rect 18956 12962 19124 12964
rect 18956 12910 18958 12962
rect 19010 12910 19124 12962
rect 18956 12908 19124 12910
rect 18956 12898 19012 12908
rect 17500 12338 17556 12348
rect 18284 12796 18396 12852
rect 17500 11284 17556 11294
rect 17164 11282 17556 11284
rect 17164 11230 17502 11282
rect 17554 11230 17556 11282
rect 17164 11228 17556 11230
rect 16492 10836 16548 10846
rect 16268 10834 16548 10836
rect 16268 10782 16494 10834
rect 16546 10782 16548 10834
rect 16268 10780 16548 10782
rect 15932 10770 15988 10780
rect 16492 10770 16548 10780
rect 15260 10668 15876 10724
rect 15036 9826 15092 9838
rect 15036 9774 15038 9826
rect 15090 9774 15092 9826
rect 14812 9716 14868 9726
rect 14700 9714 14868 9716
rect 14700 9662 14814 9714
rect 14866 9662 14868 9714
rect 14700 9660 14868 9662
rect 12860 9436 13124 9446
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 12860 9370 13124 9380
rect 14812 9380 14868 9660
rect 14812 9314 14868 9324
rect 14924 9602 14980 9614
rect 14924 9550 14926 9602
rect 14978 9550 14980 9602
rect 14700 9156 14756 9166
rect 14924 9156 14980 9550
rect 14700 9154 14980 9156
rect 14700 9102 14702 9154
rect 14754 9102 14980 9154
rect 14700 9100 14980 9102
rect 14700 9090 14756 9100
rect 11900 9042 12516 9044
rect 11900 8990 11902 9042
rect 11954 8990 12516 9042
rect 11900 8988 12516 8990
rect 12572 9044 12628 9054
rect 10612 7644 10948 7700
rect 11004 8146 11060 8158
rect 11004 8094 11006 8146
rect 11058 8094 11060 8146
rect 10556 7586 10612 7644
rect 10556 7534 10558 7586
rect 10610 7534 10612 7586
rect 10556 7522 10612 7534
rect 11004 7364 11060 8094
rect 11564 8148 11620 8158
rect 11900 8148 11956 8988
rect 12572 8930 12628 8988
rect 12572 8878 12574 8930
rect 12626 8878 12628 8930
rect 12572 8866 12628 8878
rect 15036 8428 15092 9774
rect 15260 9826 15316 10668
rect 15820 10612 15876 10668
rect 16380 10612 16436 10622
rect 15820 10610 16436 10612
rect 15820 10558 16382 10610
rect 16434 10558 16436 10610
rect 15820 10556 16436 10558
rect 15484 10500 15540 10510
rect 15484 10498 15652 10500
rect 15484 10446 15486 10498
rect 15538 10446 15652 10498
rect 15484 10444 15652 10446
rect 15484 10434 15540 10444
rect 15260 9774 15262 9826
rect 15314 9774 15316 9826
rect 15260 9762 15316 9774
rect 15596 10388 15652 10444
rect 16268 10388 16324 10398
rect 15596 10386 16324 10388
rect 15596 10334 16270 10386
rect 16322 10334 16324 10386
rect 15596 10332 16324 10334
rect 15372 9044 15428 9054
rect 15036 8372 15316 8428
rect 15260 8370 15316 8372
rect 15260 8318 15262 8370
rect 15314 8318 15316 8370
rect 15260 8306 15316 8318
rect 15372 8370 15428 8988
rect 15484 9042 15540 9054
rect 15484 8990 15486 9042
rect 15538 8990 15540 9042
rect 15484 8932 15540 8990
rect 15484 8866 15540 8876
rect 15372 8318 15374 8370
rect 15426 8318 15428 8370
rect 15372 8306 15428 8318
rect 11564 8146 11956 8148
rect 11564 8094 11566 8146
rect 11618 8094 11956 8146
rect 11564 8092 11956 8094
rect 11564 8082 11620 8092
rect 12124 8036 12180 8046
rect 12124 8034 12628 8036
rect 12124 7982 12126 8034
rect 12178 7982 12628 8034
rect 12124 7980 12628 7982
rect 12124 7970 12180 7980
rect 11116 7588 11172 7598
rect 12012 7588 12068 7598
rect 11172 7532 11396 7588
rect 11116 7494 11172 7532
rect 11004 7298 11060 7308
rect 10108 6748 10500 6804
rect 9996 6692 10052 6702
rect 10108 6692 10164 6748
rect 9996 6690 10164 6692
rect 9996 6638 9998 6690
rect 10050 6638 10164 6690
rect 9996 6636 10164 6638
rect 9996 6626 10052 6636
rect 9772 6526 9774 6578
rect 9826 6526 9828 6578
rect 9772 6514 9828 6526
rect 11340 5794 11396 7532
rect 12012 7474 12068 7532
rect 12572 7586 12628 7980
rect 12860 7868 13124 7878
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 12860 7802 13124 7812
rect 12572 7534 12574 7586
rect 12626 7534 12628 7586
rect 12572 7522 12628 7534
rect 12796 7588 12852 7598
rect 12012 7422 12014 7474
rect 12066 7422 12068 7474
rect 12012 7410 12068 7422
rect 12796 7474 12852 7532
rect 15596 7588 15652 10332
rect 16268 10322 16324 10332
rect 15772 10220 16036 10230
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 15772 10154 16036 10164
rect 16380 10052 16436 10556
rect 16044 9996 16436 10052
rect 17388 10610 17444 11228
rect 17500 11218 17556 11228
rect 17388 10558 17390 10610
rect 17442 10558 17444 10610
rect 17388 10164 17444 10558
rect 16044 9266 16100 9996
rect 16044 9214 16046 9266
rect 16098 9214 16100 9266
rect 16044 9202 16100 9214
rect 16380 9268 16436 9278
rect 16380 9174 16436 9212
rect 15820 9044 15876 9054
rect 15820 8950 15876 8988
rect 16268 9042 16324 9054
rect 16268 8990 16270 9042
rect 16322 8990 16324 9042
rect 16156 8930 16212 8942
rect 16156 8878 16158 8930
rect 16210 8878 16212 8930
rect 15772 8652 16036 8662
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 15772 8586 16036 8596
rect 16156 8484 16212 8878
rect 15708 8428 16212 8484
rect 15708 8370 15764 8428
rect 15708 8318 15710 8370
rect 15762 8318 15764 8370
rect 15708 8306 15764 8318
rect 15820 8036 15876 8046
rect 15820 8034 16100 8036
rect 15820 7982 15822 8034
rect 15874 7982 16100 8034
rect 15820 7980 16100 7982
rect 15820 7970 15876 7980
rect 15596 7522 15652 7532
rect 16044 7586 16100 7980
rect 16044 7534 16046 7586
rect 16098 7534 16100 7586
rect 16044 7522 16100 7534
rect 12796 7422 12798 7474
rect 12850 7422 12852 7474
rect 12796 7410 12852 7422
rect 13916 7364 13972 7374
rect 13916 7270 13972 7308
rect 16268 7364 16324 8990
rect 17388 9042 17444 10108
rect 18172 10498 18228 10510
rect 18172 10446 18174 10498
rect 18226 10446 18228 10498
rect 18172 10050 18228 10446
rect 18172 9998 18174 10050
rect 18226 9998 18228 10050
rect 18172 9986 18228 9998
rect 18172 9716 18228 9726
rect 18172 9154 18228 9660
rect 18172 9102 18174 9154
rect 18226 9102 18228 9154
rect 18172 9090 18228 9102
rect 18284 9714 18340 12796
rect 18396 12786 18452 12796
rect 18684 12572 18948 12582
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18684 12506 18948 12516
rect 19068 12404 19124 12908
rect 19180 12962 19236 12974
rect 19180 12910 19182 12962
rect 19234 12910 19236 12962
rect 19180 12628 19236 12910
rect 19180 12572 19460 12628
rect 19292 12404 19348 12414
rect 19068 12348 19292 12404
rect 19292 12310 19348 12348
rect 19180 12180 19236 12190
rect 19404 12180 19460 12572
rect 19628 12404 19684 13806
rect 19964 13748 20020 13758
rect 19964 13654 20020 13692
rect 20300 13748 20356 14588
rect 20412 14578 20468 14588
rect 20300 13682 20356 13692
rect 20412 13748 20468 13758
rect 20636 13748 20692 16156
rect 20412 13746 20692 13748
rect 20412 13694 20414 13746
rect 20466 13694 20692 13746
rect 20412 13692 20692 13694
rect 20748 17444 20804 17454
rect 20860 17444 20916 19406
rect 21308 19236 21364 20078
rect 21532 20020 21588 20526
rect 21868 20580 21924 20972
rect 21868 20514 21924 20524
rect 21980 20802 22036 20814
rect 21980 20750 21982 20802
rect 22034 20750 22036 20802
rect 21868 20244 21924 20254
rect 21868 20130 21924 20188
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 20066 21924 20078
rect 21532 19954 21588 19964
rect 21644 20018 21700 20030
rect 21644 19966 21646 20018
rect 21698 19966 21700 20018
rect 21644 19796 21700 19966
rect 21980 19906 22036 20750
rect 22428 20804 22484 20814
rect 22428 20710 22484 20748
rect 23212 20804 23268 20814
rect 23212 20710 23268 20748
rect 23548 20802 23604 21532
rect 23548 20750 23550 20802
rect 23602 20750 23604 20802
rect 23548 20738 23604 20750
rect 23212 20244 23268 20254
rect 21980 19854 21982 19906
rect 22034 19854 22036 19906
rect 21980 19842 22036 19854
rect 22092 20130 22148 20142
rect 22092 20078 22094 20130
rect 22146 20078 22148 20130
rect 21644 19730 21700 19740
rect 21596 19628 21860 19638
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21596 19562 21860 19572
rect 21420 19460 21476 19470
rect 21420 19346 21476 19404
rect 21644 19460 21700 19470
rect 21644 19366 21700 19404
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 21420 19282 21476 19294
rect 21532 19348 21588 19358
rect 21308 19170 21364 19180
rect 21420 19124 21476 19134
rect 21532 19124 21588 19292
rect 22092 19348 22148 20078
rect 22092 19282 22148 19292
rect 22428 20130 22484 20142
rect 22428 20078 22430 20130
rect 22482 20078 22484 20130
rect 21420 19122 21588 19124
rect 21420 19070 21422 19122
rect 21474 19070 21588 19122
rect 21420 19068 21588 19070
rect 21980 19122 22036 19134
rect 21980 19070 21982 19122
rect 22034 19070 22036 19122
rect 21420 19058 21476 19068
rect 21532 18228 21588 18238
rect 20804 17388 20916 17444
rect 21420 18172 21532 18228
rect 20412 13412 20468 13692
rect 20412 13346 20468 13356
rect 20524 13524 20580 13534
rect 20188 13076 20244 13086
rect 20524 13076 20580 13468
rect 20748 13188 20804 17388
rect 21308 16548 21364 16558
rect 21308 16210 21364 16492
rect 21420 16324 21476 18172
rect 21532 18162 21588 18172
rect 21868 18228 21924 18238
rect 21980 18228 22036 19070
rect 22092 19012 22148 19022
rect 22092 18918 22148 18956
rect 22204 19010 22260 19022
rect 22204 18958 22206 19010
rect 22258 18958 22260 19010
rect 21924 18172 22036 18228
rect 21868 18162 21924 18172
rect 22204 18116 22260 18958
rect 21596 18060 21860 18070
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21596 17994 21860 18004
rect 21980 18060 22260 18116
rect 21980 17780 22036 18060
rect 21980 17686 22036 17724
rect 22316 17668 22372 17678
rect 22428 17668 22484 20078
rect 22764 20018 22820 20030
rect 22764 19966 22766 20018
rect 22818 19966 22820 20018
rect 22764 18676 22820 19966
rect 23212 20018 23268 20188
rect 23212 19966 23214 20018
rect 23266 19966 23268 20018
rect 23212 19954 23268 19966
rect 23660 20018 23716 21868
rect 24108 21476 24164 21486
rect 23996 21474 24164 21476
rect 23996 21422 24110 21474
rect 24162 21422 24164 21474
rect 23996 21420 24164 21422
rect 23996 20804 24052 21420
rect 24108 21410 24164 21420
rect 23996 20738 24052 20748
rect 24108 20692 24164 20702
rect 24108 20690 24948 20692
rect 24108 20638 24110 20690
rect 24162 20638 24948 20690
rect 24108 20636 24948 20638
rect 24108 20626 24164 20636
rect 24508 20412 24772 20422
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24508 20346 24772 20356
rect 23660 19966 23662 20018
rect 23714 19966 23716 20018
rect 23660 19954 23716 19966
rect 24108 19908 24164 19918
rect 23996 19906 24164 19908
rect 23996 19854 24110 19906
rect 24162 19854 24164 19906
rect 23996 19852 24164 19854
rect 22876 19348 22932 19358
rect 22876 19254 22932 19292
rect 22988 19236 23044 19246
rect 22988 19142 23044 19180
rect 22764 18610 22820 18620
rect 23660 19122 23716 19134
rect 23660 19070 23662 19122
rect 23714 19070 23716 19122
rect 23548 18452 23604 18462
rect 23548 18358 23604 18396
rect 22876 18340 22932 18350
rect 22876 18246 22932 18284
rect 22316 17666 22484 17668
rect 22316 17614 22318 17666
rect 22370 17614 22484 17666
rect 22316 17612 22484 17614
rect 23100 17892 23156 17902
rect 22316 17602 22372 17612
rect 22764 17556 22820 17566
rect 22652 17554 22820 17556
rect 22652 17502 22766 17554
rect 22818 17502 22820 17554
rect 22652 17500 22820 17502
rect 21980 17444 22036 17454
rect 21596 16492 21860 16502
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21596 16426 21860 16436
rect 21868 16324 21924 16334
rect 21420 16322 21924 16324
rect 21420 16270 21870 16322
rect 21922 16270 21924 16322
rect 21420 16268 21924 16270
rect 21868 16258 21924 16268
rect 21308 16158 21310 16210
rect 21362 16158 21364 16210
rect 21308 15316 21364 16158
rect 21308 15250 21364 15260
rect 21532 16100 21588 16110
rect 21532 15148 21588 16044
rect 21980 15538 22036 17388
rect 21980 15486 21982 15538
rect 22034 15486 22036 15538
rect 21980 15474 22036 15486
rect 22316 16884 22372 16894
rect 20188 13074 20580 13076
rect 20188 13022 20190 13074
rect 20242 13022 20580 13074
rect 20188 13020 20580 13022
rect 20188 13010 20244 13020
rect 20524 12962 20580 13020
rect 20524 12910 20526 12962
rect 20578 12910 20580 12962
rect 20524 12898 20580 12910
rect 20636 13132 20804 13188
rect 20972 15092 21588 15148
rect 21756 15426 21812 15438
rect 21756 15374 21758 15426
rect 21810 15374 21812 15426
rect 21644 15092 21700 15102
rect 20972 13188 21028 15092
rect 21756 15092 21812 15374
rect 21980 15316 22036 15326
rect 21868 15092 21924 15102
rect 21756 15036 21868 15092
rect 21644 14998 21700 15036
rect 21868 15026 21924 15036
rect 21596 14924 21860 14934
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21596 14858 21860 14868
rect 21980 14642 22036 15260
rect 22316 15314 22372 16828
rect 22652 16772 22708 17500
rect 22764 17490 22820 17500
rect 23100 17106 23156 17836
rect 23660 17220 23716 19070
rect 23884 17444 23940 17454
rect 23884 17350 23940 17388
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 23100 17042 23156 17054
rect 23548 17164 23716 17220
rect 23436 16996 23492 17006
rect 23324 16884 23380 16894
rect 22540 16716 22708 16772
rect 23212 16828 23324 16884
rect 22540 15986 22596 16716
rect 22540 15934 22542 15986
rect 22594 15934 22596 15986
rect 22540 15922 22596 15934
rect 23100 16098 23156 16110
rect 23100 16046 23102 16098
rect 23154 16046 23156 16098
rect 22316 15262 22318 15314
rect 22370 15262 22372 15314
rect 22316 15250 22372 15262
rect 22428 15484 22708 15540
rect 21980 14590 21982 14642
rect 22034 14590 22036 14642
rect 21980 14578 22036 14590
rect 22316 14530 22372 14542
rect 22316 14478 22318 14530
rect 22370 14478 22372 14530
rect 21420 14306 21476 14318
rect 21420 14254 21422 14306
rect 21474 14254 21476 14306
rect 21084 13634 21140 13646
rect 21084 13582 21086 13634
rect 21138 13582 21140 13634
rect 21084 13300 21140 13582
rect 21420 13412 21476 14254
rect 22316 13972 22372 14478
rect 22316 13906 22372 13916
rect 21084 13244 21364 13300
rect 20972 13132 21252 13188
rect 20636 12404 20692 13132
rect 20748 12964 20804 12974
rect 20748 12850 20804 12908
rect 20748 12798 20750 12850
rect 20802 12798 20804 12850
rect 20748 12786 20804 12798
rect 19628 12338 19684 12348
rect 20412 12348 20692 12404
rect 20860 12404 20916 12414
rect 19740 12290 19796 12302
rect 19740 12238 19742 12290
rect 19794 12238 19796 12290
rect 19740 12180 19796 12238
rect 19180 12178 19796 12180
rect 19180 12126 19182 12178
rect 19234 12126 19796 12178
rect 19180 12124 19796 12126
rect 19180 12114 19236 12124
rect 19292 11956 19348 11966
rect 19180 11954 19348 11956
rect 19180 11902 19294 11954
rect 19346 11902 19348 11954
rect 19180 11900 19348 11902
rect 18684 11004 18948 11014
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18684 10938 18948 10948
rect 19180 9938 19236 11900
rect 19292 11890 19348 11900
rect 19740 11844 19796 12124
rect 19740 11778 19796 11788
rect 20076 12178 20132 12190
rect 20076 12126 20078 12178
rect 20130 12126 20132 12178
rect 20076 11396 20132 12126
rect 20300 12178 20356 12190
rect 20300 12126 20302 12178
rect 20354 12126 20356 12178
rect 20300 11844 20356 12126
rect 20300 11778 20356 11788
rect 20076 11330 20132 11340
rect 19628 10612 19684 10622
rect 19180 9886 19182 9938
rect 19234 9886 19236 9938
rect 19180 9874 19236 9886
rect 19516 10388 19572 10398
rect 19516 9826 19572 10332
rect 19516 9774 19518 9826
rect 19570 9774 19572 9826
rect 19516 9762 19572 9774
rect 18284 9662 18286 9714
rect 18338 9662 18340 9714
rect 17388 8990 17390 9042
rect 17442 8990 17444 9042
rect 16268 7298 16324 7308
rect 16828 8932 16884 8942
rect 16828 7474 16884 8876
rect 17388 8932 17444 8990
rect 17388 8866 17444 8876
rect 16828 7422 16830 7474
rect 16882 7422 16884 7474
rect 11676 7250 11732 7262
rect 11676 7198 11678 7250
rect 11730 7198 11732 7250
rect 11676 6692 11732 7198
rect 15772 7084 16036 7094
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 15772 7018 16036 7028
rect 11788 6692 11844 6702
rect 11676 6690 11844 6692
rect 11676 6638 11790 6690
rect 11842 6638 11844 6690
rect 11676 6636 11844 6638
rect 16828 6692 16884 7422
rect 17052 6692 17108 6702
rect 16828 6690 17108 6692
rect 16828 6638 17054 6690
rect 17106 6638 17108 6690
rect 16828 6636 17108 6638
rect 11788 6626 11844 6636
rect 12124 6468 12180 6478
rect 12124 6374 12180 6412
rect 13468 6468 13524 6478
rect 12860 6300 13124 6310
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 12860 6234 13124 6244
rect 13468 6018 13524 6412
rect 13468 5966 13470 6018
rect 13522 5966 13524 6018
rect 13468 5954 13524 5966
rect 14252 5908 14308 5918
rect 14252 5814 14308 5852
rect 17052 5908 17108 6636
rect 18284 6692 18340 9662
rect 18508 9716 18564 9726
rect 18844 9716 18900 9726
rect 18508 9714 18900 9716
rect 18508 9662 18510 9714
rect 18562 9662 18846 9714
rect 18898 9662 18900 9714
rect 18508 9660 18900 9662
rect 18508 9650 18564 9660
rect 18844 9650 18900 9660
rect 18684 9436 18948 9446
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18684 9370 18948 9380
rect 19628 8258 19684 10556
rect 20300 10498 20356 10510
rect 20300 10446 20302 10498
rect 20354 10446 20356 10498
rect 20300 10388 20356 10446
rect 20300 10322 20356 10332
rect 20300 9940 20356 9950
rect 20412 9940 20468 12348
rect 20860 12290 20916 12348
rect 20860 12238 20862 12290
rect 20914 12238 20916 12290
rect 20636 12178 20692 12190
rect 20636 12126 20638 12178
rect 20690 12126 20692 12178
rect 20636 11284 20692 12126
rect 20860 11956 20916 12238
rect 21196 12292 21252 13132
rect 21308 13186 21364 13244
rect 21308 13134 21310 13186
rect 21362 13134 21364 13186
rect 21308 13122 21364 13134
rect 21308 12962 21364 12974
rect 21308 12910 21310 12962
rect 21362 12910 21364 12962
rect 21308 12852 21364 12910
rect 21308 12786 21364 12796
rect 21420 12404 21476 13356
rect 21596 13356 21860 13366
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21596 13290 21860 13300
rect 21644 12852 21700 12862
rect 22204 12852 22260 12862
rect 21644 12850 22148 12852
rect 21644 12798 21646 12850
rect 21698 12798 22148 12850
rect 21644 12796 22148 12798
rect 21644 12786 21700 12796
rect 21532 12404 21588 12414
rect 21420 12348 21532 12404
rect 21532 12338 21588 12348
rect 22092 12292 22148 12796
rect 22204 12758 22260 12796
rect 22204 12292 22260 12302
rect 21196 12236 21476 12292
rect 22092 12290 22260 12292
rect 22092 12238 22206 12290
rect 22258 12238 22260 12290
rect 22092 12236 22260 12238
rect 20972 12068 21028 12078
rect 21308 12068 21364 12078
rect 20972 12066 21364 12068
rect 20972 12014 20974 12066
rect 21026 12014 21310 12066
rect 21362 12014 21364 12066
rect 20972 12012 21364 12014
rect 20972 12002 21028 12012
rect 21308 12002 21364 12012
rect 20860 11890 20916 11900
rect 20636 10388 20692 11228
rect 21084 11844 21140 11854
rect 21420 11844 21476 12236
rect 22204 12226 22260 12236
rect 21756 12178 21812 12190
rect 21756 12126 21758 12178
rect 21810 12126 21812 12178
rect 21756 12068 21812 12126
rect 21980 12068 22036 12078
rect 21756 12012 21980 12068
rect 20972 10500 21028 10510
rect 20636 10322 20692 10332
rect 20748 10444 20972 10500
rect 20300 9938 20468 9940
rect 20300 9886 20302 9938
rect 20354 9886 20468 9938
rect 20300 9884 20468 9886
rect 20188 9716 20244 9726
rect 20188 9622 20244 9660
rect 20300 9156 20356 9884
rect 20524 9828 20580 9838
rect 20188 9100 20356 9156
rect 20412 9826 20580 9828
rect 20412 9774 20526 9826
rect 20578 9774 20580 9826
rect 20412 9772 20580 9774
rect 19628 8206 19630 8258
rect 19682 8206 19684 8258
rect 18684 7868 18948 7878
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18684 7802 18948 7812
rect 19628 7700 19684 8206
rect 19852 8932 19908 8942
rect 19852 8258 19908 8876
rect 20188 8820 20244 9100
rect 20300 8932 20356 8942
rect 20300 8838 20356 8876
rect 20188 8754 20244 8764
rect 20300 8484 20356 8494
rect 20412 8484 20468 9772
rect 20524 9762 20580 9772
rect 20748 9826 20804 10444
rect 20972 10434 21028 10444
rect 20748 9774 20750 9826
rect 20802 9774 20804 9826
rect 20748 9762 20804 9774
rect 20972 10052 21028 10062
rect 20636 9492 20692 9502
rect 20636 8932 20692 9436
rect 20748 9268 20804 9278
rect 20748 9042 20804 9212
rect 20972 9266 21028 9996
rect 20972 9214 20974 9266
rect 21026 9214 21028 9266
rect 20972 9202 21028 9214
rect 20748 8990 20750 9042
rect 20802 8990 20804 9042
rect 20748 8978 20804 8990
rect 20636 8866 20692 8876
rect 21084 8708 21140 11788
rect 21196 11788 21476 11844
rect 21596 11788 21860 11798
rect 21196 11618 21252 11788
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21596 11722 21860 11732
rect 21980 11620 22036 12012
rect 21196 11566 21198 11618
rect 21250 11566 21252 11618
rect 21196 11554 21252 11566
rect 21868 11564 22036 11620
rect 22092 11956 22148 11966
rect 21420 11396 21476 11406
rect 21196 11340 21420 11396
rect 21196 9266 21252 11340
rect 21420 11302 21476 11340
rect 21868 11394 21924 11564
rect 21868 11342 21870 11394
rect 21922 11342 21924 11394
rect 21868 11330 21924 11342
rect 22092 11394 22148 11900
rect 22092 11342 22094 11394
rect 22146 11342 22148 11394
rect 22092 11330 22148 11342
rect 21980 11284 22036 11294
rect 21980 11190 22036 11228
rect 21420 10610 21476 10622
rect 21420 10558 21422 10610
rect 21474 10558 21476 10610
rect 21196 9214 21198 9266
rect 21250 9214 21252 9266
rect 21196 9202 21252 9214
rect 21308 10164 21364 10174
rect 21308 9826 21364 10108
rect 21308 9774 21310 9826
rect 21362 9774 21364 9826
rect 21308 8820 21364 9774
rect 21420 9156 21476 10558
rect 21644 10612 21700 10622
rect 21644 10518 21700 10556
rect 21980 10610 22036 10622
rect 21980 10558 21982 10610
rect 22034 10558 22036 10610
rect 21532 10500 21588 10510
rect 21532 10406 21588 10444
rect 21596 10220 21860 10230
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21596 10154 21860 10164
rect 21868 9380 21924 9390
rect 21980 9380 22036 10558
rect 22428 10276 22484 15484
rect 22652 15426 22708 15484
rect 22652 15374 22654 15426
rect 22706 15374 22708 15426
rect 22652 15362 22708 15374
rect 22540 15314 22596 15326
rect 22540 15262 22542 15314
rect 22594 15262 22596 15314
rect 22540 15148 22596 15262
rect 23100 15148 23156 16046
rect 23212 15874 23268 16828
rect 23324 16818 23380 16828
rect 23436 16882 23492 16940
rect 23436 16830 23438 16882
rect 23490 16830 23492 16882
rect 23436 16818 23492 16830
rect 23548 16324 23604 17164
rect 23660 16884 23716 16894
rect 23660 16790 23716 16828
rect 23884 16884 23940 16894
rect 23884 16790 23940 16828
rect 23212 15822 23214 15874
rect 23266 15822 23268 15874
rect 23212 15810 23268 15822
rect 23436 16268 23604 16324
rect 23436 15876 23492 16268
rect 23548 16100 23604 16110
rect 23548 16098 23716 16100
rect 23548 16046 23550 16098
rect 23602 16046 23716 16098
rect 23548 16044 23716 16046
rect 23548 16034 23604 16044
rect 23436 15820 23604 15876
rect 23548 15314 23604 15820
rect 23548 15262 23550 15314
rect 23602 15262 23604 15314
rect 23548 15250 23604 15262
rect 22540 15092 22820 15148
rect 23100 15092 23380 15148
rect 23660 15092 23716 16044
rect 23996 15988 24052 19852
rect 24108 19842 24164 19852
rect 24108 19010 24164 19022
rect 24108 18958 24110 19010
rect 24162 18958 24164 19010
rect 24108 18676 24164 18958
rect 24508 18844 24772 18854
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24508 18778 24772 18788
rect 24108 18610 24164 18620
rect 24108 18452 24164 18462
rect 24108 18358 24164 18396
rect 24108 17666 24164 17678
rect 24108 17614 24110 17666
rect 24162 17614 24164 17666
rect 24108 16884 24164 17614
rect 24508 17276 24772 17286
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24508 17210 24772 17220
rect 24108 16818 24164 16828
rect 24220 16882 24276 16894
rect 24220 16830 24222 16882
rect 24274 16830 24276 16882
rect 24108 15988 24164 15998
rect 23996 15986 24164 15988
rect 23996 15934 24110 15986
rect 24162 15934 24164 15986
rect 23996 15932 24164 15934
rect 24108 15922 24164 15932
rect 24220 15652 24276 16830
rect 23996 15596 24276 15652
rect 23996 15538 24052 15596
rect 23996 15486 23998 15538
rect 24050 15486 24052 15538
rect 23996 15474 24052 15486
rect 24108 15426 24164 15438
rect 24108 15374 24110 15426
rect 24162 15374 24164 15426
rect 24108 15148 24164 15374
rect 22764 14642 22820 15092
rect 22764 14590 22766 14642
rect 22818 14590 22820 14642
rect 22764 14578 22820 14590
rect 23212 13634 23268 13646
rect 23212 13582 23214 13634
rect 23266 13582 23268 13634
rect 23212 13300 23268 13582
rect 22876 13244 23268 13300
rect 22876 12964 22932 13244
rect 22988 12964 23044 12974
rect 22876 12962 23044 12964
rect 22876 12910 22990 12962
rect 23042 12910 23044 12962
rect 22876 12908 23044 12910
rect 22540 12738 22596 12750
rect 22540 12686 22542 12738
rect 22594 12686 22596 12738
rect 22540 11732 22596 12686
rect 22764 12404 22820 12414
rect 22764 12310 22820 12348
rect 22988 12068 23044 12908
rect 23212 12964 23268 12974
rect 23212 12870 23268 12908
rect 23324 12740 23380 15092
rect 23436 15036 23716 15092
rect 23884 15092 23940 15102
rect 23436 14868 23492 15036
rect 23660 14868 23716 14878
rect 23436 14812 23660 14868
rect 23660 14802 23716 14812
rect 23436 14644 23492 14654
rect 23492 14588 23548 14644
rect 23436 14578 23548 14588
rect 23492 14532 23548 14578
rect 23660 14642 23716 14654
rect 23660 14590 23662 14642
rect 23714 14590 23716 14642
rect 23660 14532 23716 14590
rect 23492 14476 23716 14532
rect 23884 14418 23940 15036
rect 23884 14366 23886 14418
rect 23938 14366 23940 14418
rect 23884 14354 23940 14366
rect 23996 15092 24164 15148
rect 23100 12684 23380 12740
rect 23660 14308 23716 14318
rect 23100 12290 23156 12684
rect 23100 12238 23102 12290
rect 23154 12238 23156 12290
rect 23100 12226 23156 12238
rect 22988 12002 23044 12012
rect 23548 12178 23604 12190
rect 23548 12126 23550 12178
rect 23602 12126 23604 12178
rect 22540 11676 23268 11732
rect 23100 11394 23156 11406
rect 23100 11342 23102 11394
rect 23154 11342 23156 11394
rect 22540 11282 22596 11294
rect 22540 11230 22542 11282
rect 22594 11230 22596 11282
rect 22540 10724 22596 11230
rect 22652 10724 22708 10734
rect 22540 10722 22708 10724
rect 22540 10670 22654 10722
rect 22706 10670 22708 10722
rect 22540 10668 22708 10670
rect 22652 10658 22708 10668
rect 23100 10388 23156 11342
rect 23212 10610 23268 11676
rect 23548 11620 23604 12126
rect 23436 11564 23604 11620
rect 23212 10558 23214 10610
rect 23266 10558 23268 10610
rect 23212 10546 23268 10558
rect 23324 11284 23380 11294
rect 23324 10500 23380 11228
rect 23436 11172 23492 11564
rect 23660 11508 23716 14252
rect 23884 13972 23940 13982
rect 23884 13878 23940 13916
rect 23884 13076 23940 13086
rect 23996 13076 24052 15092
rect 24220 14530 24276 15596
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 24220 14466 24276 14478
rect 24332 15988 24388 15998
rect 24332 14756 24388 15932
rect 24508 15708 24772 15718
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24508 15642 24772 15652
rect 24332 14308 24388 14700
rect 24108 14252 24388 14308
rect 24108 13746 24164 14252
rect 24508 14140 24772 14150
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24508 14074 24772 14084
rect 24108 13694 24110 13746
rect 24162 13694 24164 13746
rect 24108 13682 24164 13694
rect 24220 13748 24276 13758
rect 24220 13524 24276 13692
rect 23884 13074 24052 13076
rect 23884 13022 23886 13074
rect 23938 13022 24052 13074
rect 23884 13020 24052 13022
rect 24108 13468 24276 13524
rect 23884 13010 23940 13020
rect 23996 12180 24052 12190
rect 24108 12180 24164 13468
rect 24220 12852 24276 12862
rect 24276 12796 24388 12852
rect 24220 12786 24276 12796
rect 23996 12178 24164 12180
rect 23996 12126 23998 12178
rect 24050 12126 24164 12178
rect 23996 12124 24164 12126
rect 24220 12628 24276 12638
rect 23996 12114 24052 12124
rect 23772 11508 23828 11518
rect 23660 11506 23828 11508
rect 23660 11454 23774 11506
rect 23826 11454 23828 11506
rect 23660 11452 23828 11454
rect 23772 11442 23828 11452
rect 23548 11396 23604 11406
rect 23548 11302 23604 11340
rect 24108 11284 24164 11294
rect 23996 11282 24164 11284
rect 23996 11230 24110 11282
rect 24162 11230 24164 11282
rect 23996 11228 24164 11230
rect 23436 11116 23604 11172
rect 23436 10500 23492 10510
rect 23324 10498 23492 10500
rect 23324 10446 23438 10498
rect 23490 10446 23492 10498
rect 23324 10444 23492 10446
rect 23436 10434 23492 10444
rect 23100 10332 23268 10388
rect 22428 10220 23156 10276
rect 22764 9940 22820 9950
rect 21924 9324 22036 9380
rect 22092 9714 22148 9726
rect 22092 9662 22094 9714
rect 22146 9662 22148 9714
rect 21420 9090 21476 9100
rect 21756 9156 21812 9166
rect 21644 9044 21700 9054
rect 21644 8950 21700 8988
rect 21756 8932 21812 9100
rect 21868 9154 21924 9324
rect 21868 9102 21870 9154
rect 21922 9102 21924 9154
rect 21868 9090 21924 9102
rect 21980 9042 22036 9054
rect 21980 8990 21982 9042
rect 22034 8990 22036 9042
rect 21980 8932 22036 8990
rect 21756 8876 22036 8932
rect 21308 8764 21476 8820
rect 21196 8708 21252 8718
rect 21084 8652 21196 8708
rect 21196 8642 21252 8652
rect 20300 8482 21364 8484
rect 20300 8430 20302 8482
rect 20354 8430 21364 8482
rect 20300 8428 21364 8430
rect 20300 8418 20356 8428
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8194 19908 8206
rect 19740 8146 19796 8158
rect 19740 8094 19742 8146
rect 19794 8094 19796 8146
rect 19740 7924 19796 8094
rect 19740 7868 19908 7924
rect 19740 7700 19796 7710
rect 19628 7698 19796 7700
rect 19628 7646 19742 7698
rect 19794 7646 19796 7698
rect 19628 7644 19796 7646
rect 18340 6636 18452 6692
rect 18284 6626 18340 6636
rect 17836 6578 17892 6590
rect 17836 6526 17838 6578
rect 17890 6526 17892 6578
rect 17836 6132 17892 6526
rect 17836 6066 17892 6076
rect 18396 6018 18452 6636
rect 18684 6300 18948 6310
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18684 6234 18948 6244
rect 18508 6132 18564 6142
rect 18508 6038 18564 6076
rect 18732 6132 18788 6142
rect 18396 5966 18398 6018
rect 18450 5966 18452 6018
rect 18396 5954 18452 5966
rect 17052 5842 17108 5852
rect 18732 5906 18788 6076
rect 18732 5854 18734 5906
rect 18786 5854 18788 5906
rect 18732 5842 18788 5854
rect 19740 6132 19796 7644
rect 19740 5906 19796 6076
rect 19740 5854 19742 5906
rect 19794 5854 19796 5906
rect 19740 5842 19796 5854
rect 19852 5908 19908 7868
rect 21308 7586 21364 8428
rect 21308 7534 21310 7586
rect 21362 7534 21364 7586
rect 21308 7522 21364 7534
rect 20076 7476 20132 7486
rect 19964 6804 20020 6814
rect 20076 6804 20132 7420
rect 19964 6802 20132 6804
rect 19964 6750 19966 6802
rect 20018 6750 20132 6802
rect 19964 6748 20132 6750
rect 20748 6802 20804 6814
rect 20748 6750 20750 6802
rect 20802 6750 20804 6802
rect 19964 6738 20020 6748
rect 20636 6692 20692 6702
rect 20412 6580 20468 6590
rect 20412 6578 20580 6580
rect 20412 6526 20414 6578
rect 20466 6526 20580 6578
rect 20412 6524 20580 6526
rect 20412 6514 20468 6524
rect 19964 5908 20020 5918
rect 19852 5852 19964 5908
rect 19964 5842 20020 5852
rect 20412 5908 20468 5918
rect 20412 5814 20468 5852
rect 11340 5742 11342 5794
rect 11394 5742 11396 5794
rect 11340 5730 11396 5742
rect 20524 5794 20580 6524
rect 20636 6578 20692 6636
rect 20636 6526 20638 6578
rect 20690 6526 20692 6578
rect 20636 6514 20692 6526
rect 20748 6580 20804 6750
rect 21420 6690 21476 8764
rect 21596 8652 21860 8662
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21596 8586 21860 8596
rect 21644 8484 21700 8494
rect 21980 8428 22036 8876
rect 21644 8390 21700 8428
rect 21868 8372 22036 8428
rect 22092 8482 22148 9662
rect 22764 9268 22820 9884
rect 22764 9174 22820 9212
rect 22092 8430 22094 8482
rect 22146 8430 22148 8482
rect 22092 8418 22148 8430
rect 22204 8930 22260 8942
rect 22204 8878 22206 8930
rect 22258 8878 22260 8930
rect 21756 8258 21812 8270
rect 21756 8206 21758 8258
rect 21810 8206 21812 8258
rect 21532 7700 21588 7710
rect 21532 7606 21588 7644
rect 21644 7364 21700 7374
rect 21756 7364 21812 8206
rect 21868 7924 21924 8372
rect 21980 8260 22036 8270
rect 21980 8166 22036 8204
rect 21868 7868 22036 7924
rect 21644 7362 21812 7364
rect 21644 7310 21646 7362
rect 21698 7310 21812 7362
rect 21644 7308 21812 7310
rect 21644 7298 21700 7308
rect 21596 7084 21860 7094
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21596 7018 21860 7028
rect 21420 6638 21422 6690
rect 21474 6638 21476 6690
rect 21420 6626 21476 6638
rect 20748 6514 20804 6524
rect 21980 5908 22036 7868
rect 22204 7476 22260 8878
rect 22764 8484 22820 8494
rect 22540 8258 22596 8270
rect 22540 8206 22542 8258
rect 22594 8206 22596 8258
rect 22540 7700 22596 8206
rect 22764 8146 22820 8428
rect 23100 8370 23156 10220
rect 23100 8318 23102 8370
rect 23154 8318 23156 8370
rect 23100 8306 23156 8318
rect 23212 8148 23268 10332
rect 23548 10052 23604 11116
rect 23548 9986 23604 9996
rect 23548 9380 23604 9390
rect 23436 9042 23492 9054
rect 23436 8990 23438 9042
rect 23490 8990 23492 9042
rect 23436 8484 23492 8990
rect 23436 8418 23492 8428
rect 23548 8370 23604 9324
rect 23884 9044 23940 9054
rect 23884 8950 23940 8988
rect 23548 8318 23550 8370
rect 23602 8318 23604 8370
rect 23548 8306 23604 8318
rect 23772 8260 23828 8270
rect 23772 8258 23940 8260
rect 23772 8206 23774 8258
rect 23826 8206 23940 8258
rect 23772 8204 23940 8206
rect 23772 8194 23828 8204
rect 22764 8094 22766 8146
rect 22818 8094 22820 8146
rect 22764 8082 22820 8094
rect 22876 8092 23268 8148
rect 22652 7700 22708 7710
rect 22540 7644 22652 7700
rect 22652 7606 22708 7644
rect 22876 7586 22932 8092
rect 22876 7534 22878 7586
rect 22930 7534 22932 7586
rect 22876 7522 22932 7534
rect 22204 7410 22260 7420
rect 23324 7476 23380 7486
rect 23324 7382 23380 7420
rect 23660 7364 23716 7374
rect 23548 7362 23716 7364
rect 23548 7310 23662 7362
rect 23714 7310 23716 7362
rect 23548 7308 23716 7310
rect 23212 6804 23268 6814
rect 22092 6580 22148 6590
rect 22092 6486 22148 6524
rect 22764 6132 22820 6142
rect 23212 6132 23268 6748
rect 22764 6130 23268 6132
rect 22764 6078 22766 6130
rect 22818 6078 23268 6130
rect 22764 6076 23268 6078
rect 22764 6066 22820 6076
rect 21980 5842 22036 5852
rect 22428 6018 22484 6030
rect 22428 5966 22430 6018
rect 22482 5966 22484 6018
rect 22428 5908 22484 5966
rect 22428 5842 22484 5852
rect 23212 5906 23268 6076
rect 23212 5854 23214 5906
rect 23266 5854 23268 5906
rect 23212 5842 23268 5854
rect 20524 5742 20526 5794
rect 20578 5742 20580 5794
rect 20524 5730 20580 5742
rect 9948 5516 10212 5526
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 9948 5450 10212 5460
rect 15772 5516 16036 5526
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 15772 5450 16036 5460
rect 21596 5516 21860 5526
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21596 5450 21860 5460
rect 9884 5236 9940 5246
rect 9660 5234 9940 5236
rect 9660 5182 9886 5234
rect 9938 5182 9940 5234
rect 9660 5180 9940 5182
rect 9884 5170 9940 5180
rect 6972 5124 7028 5134
rect 6860 5122 7028 5124
rect 6860 5070 6974 5122
rect 7026 5070 7028 5122
rect 6860 5068 7028 5070
rect 6972 5058 7028 5068
rect 7036 4732 7300 4742
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7036 4666 7300 4676
rect 12860 4732 13124 4742
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 12860 4666 13124 4676
rect 18684 4732 18948 4742
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18684 4666 18948 4676
rect 4124 3948 4388 3958
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4124 3882 4388 3892
rect 9948 3948 10212 3958
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 9948 3882 10212 3892
rect 15772 3948 16036 3958
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 15772 3882 16036 3892
rect 21596 3948 21860 3958
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21596 3882 21860 3892
rect 23436 3444 23492 3482
rect 23548 3444 23604 7308
rect 23660 7298 23716 7308
rect 23660 5908 23716 5918
rect 23660 5906 23828 5908
rect 23660 5854 23662 5906
rect 23714 5854 23828 5906
rect 23660 5852 23828 5854
rect 23660 5842 23716 5852
rect 23660 5236 23716 5246
rect 23660 5142 23716 5180
rect 23772 4564 23828 5852
rect 23884 5010 23940 8204
rect 23996 6020 24052 11228
rect 24108 11218 24164 11228
rect 24220 11060 24276 12572
rect 24108 11004 24276 11060
rect 24332 11956 24388 12796
rect 24508 12572 24772 12582
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24508 12506 24772 12516
rect 24108 9154 24164 11004
rect 24220 10836 24276 10846
rect 24332 10836 24388 11900
rect 24892 11396 24948 20636
rect 24892 11330 24948 11340
rect 24508 11004 24772 11014
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24508 10938 24772 10948
rect 24220 10834 24388 10836
rect 24220 10782 24222 10834
rect 24274 10782 24388 10834
rect 24220 10780 24388 10782
rect 24220 10770 24276 10780
rect 24108 9102 24110 9154
rect 24162 9102 24164 9154
rect 24108 9090 24164 9102
rect 24220 9938 24276 9950
rect 24220 9886 24222 9938
rect 24274 9886 24276 9938
rect 24220 9044 24276 9886
rect 24508 9436 24772 9446
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24508 9370 24772 9380
rect 24220 8978 24276 8988
rect 24508 7868 24772 7878
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24508 7802 24772 7812
rect 24220 6804 24276 6814
rect 24220 6710 24276 6748
rect 24508 6300 24772 6310
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24508 6234 24772 6244
rect 24108 6020 24164 6030
rect 23996 6018 24164 6020
rect 23996 5966 24110 6018
rect 24162 5966 24164 6018
rect 23996 5964 24164 5966
rect 24108 5954 24164 5964
rect 24220 5908 24276 5918
rect 24220 5236 24276 5852
rect 24220 5122 24276 5180
rect 24220 5070 24222 5122
rect 24274 5070 24276 5122
rect 24220 5058 24276 5070
rect 23884 4958 23886 5010
rect 23938 4958 23940 5010
rect 23884 4946 23940 4958
rect 24508 4732 24772 4742
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24508 4666 24772 4676
rect 23884 4564 23940 4574
rect 23772 4562 23940 4564
rect 23772 4510 23886 4562
rect 23938 4510 23940 4562
rect 23772 4508 23940 4510
rect 23884 4498 23940 4508
rect 24220 4338 24276 4350
rect 24220 4286 24222 4338
rect 24274 4286 24276 4338
rect 23660 4228 23716 4238
rect 24220 4228 24276 4286
rect 23660 4226 24276 4228
rect 23660 4174 23662 4226
rect 23714 4174 24276 4226
rect 23660 4172 24276 4174
rect 23660 4162 23716 4172
rect 24220 3892 24276 4172
rect 24220 3826 24276 3836
rect 23660 3444 23716 3454
rect 23548 3442 23716 3444
rect 23548 3390 23662 3442
rect 23714 3390 23716 3442
rect 23548 3388 23716 3390
rect 23436 3378 23492 3388
rect 23660 3378 23716 3388
rect 23884 3444 23940 3454
rect 23996 3444 24052 3482
rect 23940 3442 24052 3444
rect 23940 3390 23998 3442
rect 24050 3390 24052 3442
rect 23940 3388 24052 3390
rect 23884 3378 23940 3388
rect 7036 3164 7300 3174
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7036 3098 7300 3108
rect 12860 3164 13124 3174
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 12860 3098 13124 3108
rect 18684 3164 18948 3174
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18684 3098 18948 3108
rect 23996 1876 24052 3388
rect 24508 3164 24772 3174
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24508 3098 24772 3108
rect 23996 1810 24052 1820
<< via2 >>
rect 4124 22762 4180 22764
rect 4124 22710 4126 22762
rect 4126 22710 4178 22762
rect 4178 22710 4180 22762
rect 4124 22708 4180 22710
rect 4228 22762 4284 22764
rect 4228 22710 4230 22762
rect 4230 22710 4282 22762
rect 4282 22710 4284 22762
rect 4228 22708 4284 22710
rect 4332 22762 4388 22764
rect 4332 22710 4334 22762
rect 4334 22710 4386 22762
rect 4386 22710 4388 22762
rect 4332 22708 4388 22710
rect 2268 21308 2324 21364
rect 4124 21194 4180 21196
rect 4124 21142 4126 21194
rect 4126 21142 4178 21194
rect 4178 21142 4180 21194
rect 4124 21140 4180 21142
rect 4228 21194 4284 21196
rect 4228 21142 4230 21194
rect 4230 21142 4282 21194
rect 4282 21142 4284 21194
rect 4228 21140 4284 21142
rect 4332 21194 4388 21196
rect 4332 21142 4334 21194
rect 4334 21142 4386 21194
rect 4386 21142 4388 21194
rect 4332 21140 4388 21142
rect 1932 18508 1988 18564
rect 4124 19626 4180 19628
rect 4124 19574 4126 19626
rect 4126 19574 4178 19626
rect 4178 19574 4180 19626
rect 4124 19572 4180 19574
rect 4228 19626 4284 19628
rect 4228 19574 4230 19626
rect 4230 19574 4282 19626
rect 4282 19574 4284 19626
rect 4228 19572 4284 19574
rect 4332 19626 4388 19628
rect 4332 19574 4334 19626
rect 4334 19574 4386 19626
rect 4386 19574 4388 19626
rect 4332 19572 4388 19574
rect 2940 18508 2996 18564
rect 2492 17836 2548 17892
rect 3612 18396 3668 18452
rect 3164 18172 3220 18228
rect 2044 16268 2100 16324
rect 3836 18284 3892 18340
rect 4396 18396 4452 18452
rect 4284 18284 4340 18340
rect 4124 18058 4180 18060
rect 4124 18006 4126 18058
rect 4126 18006 4178 18058
rect 4178 18006 4180 18058
rect 4124 18004 4180 18006
rect 4228 18058 4284 18060
rect 4228 18006 4230 18058
rect 4230 18006 4282 18058
rect 4282 18006 4284 18058
rect 4228 18004 4284 18006
rect 4332 18058 4388 18060
rect 4332 18006 4334 18058
rect 4334 18006 4386 18058
rect 4386 18006 4388 18058
rect 4332 18004 4388 18006
rect 3948 17500 4004 17556
rect 4284 17836 4340 17892
rect 3164 16994 3220 16996
rect 3164 16942 3166 16994
rect 3166 16942 3218 16994
rect 3218 16942 3220 16994
rect 3164 16940 3220 16942
rect 2492 16322 2548 16324
rect 2492 16270 2494 16322
rect 2494 16270 2546 16322
rect 2546 16270 2548 16322
rect 2492 16268 2548 16270
rect 2380 16044 2436 16100
rect 2044 15260 2100 15316
rect 1820 15036 1876 15092
rect 2492 15820 2548 15876
rect 2380 15260 2436 15316
rect 1932 14530 1988 14532
rect 1932 14478 1934 14530
rect 1934 14478 1986 14530
rect 1986 14478 1988 14530
rect 1932 14476 1988 14478
rect 2716 15372 2772 15428
rect 2604 14924 2660 14980
rect 4620 18508 4676 18564
rect 3724 16940 3780 16996
rect 3388 16268 3444 16324
rect 4396 17106 4452 17108
rect 4396 17054 4398 17106
rect 4398 17054 4450 17106
rect 4450 17054 4452 17106
rect 4396 17052 4452 17054
rect 9948 22762 10004 22764
rect 9948 22710 9950 22762
rect 9950 22710 10002 22762
rect 10002 22710 10004 22762
rect 9948 22708 10004 22710
rect 10052 22762 10108 22764
rect 10052 22710 10054 22762
rect 10054 22710 10106 22762
rect 10106 22710 10108 22762
rect 10052 22708 10108 22710
rect 10156 22762 10212 22764
rect 10156 22710 10158 22762
rect 10158 22710 10210 22762
rect 10210 22710 10212 22762
rect 10156 22708 10212 22710
rect 20300 23996 20356 24052
rect 15772 22762 15828 22764
rect 15772 22710 15774 22762
rect 15774 22710 15826 22762
rect 15826 22710 15828 22762
rect 15772 22708 15828 22710
rect 15876 22762 15932 22764
rect 15876 22710 15878 22762
rect 15878 22710 15930 22762
rect 15930 22710 15932 22762
rect 15876 22708 15932 22710
rect 15980 22762 16036 22764
rect 15980 22710 15982 22762
rect 15982 22710 16034 22762
rect 16034 22710 16036 22762
rect 15980 22708 16036 22710
rect 21596 22762 21652 22764
rect 21596 22710 21598 22762
rect 21598 22710 21650 22762
rect 21650 22710 21652 22762
rect 21596 22708 21652 22710
rect 21700 22762 21756 22764
rect 21700 22710 21702 22762
rect 21702 22710 21754 22762
rect 21754 22710 21756 22762
rect 21700 22708 21756 22710
rect 21804 22762 21860 22764
rect 21804 22710 21806 22762
rect 21806 22710 21858 22762
rect 21858 22710 21860 22762
rect 21804 22708 21860 22710
rect 21308 22540 21364 22596
rect 22428 22594 22484 22596
rect 22428 22542 22430 22594
rect 22430 22542 22482 22594
rect 22482 22542 22484 22594
rect 22428 22540 22484 22542
rect 7036 21978 7092 21980
rect 7036 21926 7038 21978
rect 7038 21926 7090 21978
rect 7090 21926 7092 21978
rect 7036 21924 7092 21926
rect 7140 21978 7196 21980
rect 7140 21926 7142 21978
rect 7142 21926 7194 21978
rect 7194 21926 7196 21978
rect 7140 21924 7196 21926
rect 7244 21978 7300 21980
rect 7244 21926 7246 21978
rect 7246 21926 7298 21978
rect 7298 21926 7300 21978
rect 7244 21924 7300 21926
rect 7644 21756 7700 21812
rect 5068 21308 5124 21364
rect 5404 19852 5460 19908
rect 5180 18620 5236 18676
rect 4956 18450 5012 18452
rect 4956 18398 4958 18450
rect 4958 18398 5010 18450
rect 5010 18398 5012 18450
rect 4956 18396 5012 18398
rect 4844 18226 4900 18228
rect 4844 18174 4846 18226
rect 4846 18174 4898 18226
rect 4898 18174 4900 18226
rect 4844 18172 4900 18174
rect 5516 18172 5572 18228
rect 5628 18396 5684 18452
rect 4124 16490 4180 16492
rect 4124 16438 4126 16490
rect 4126 16438 4178 16490
rect 4178 16438 4180 16490
rect 4124 16436 4180 16438
rect 4228 16490 4284 16492
rect 4228 16438 4230 16490
rect 4230 16438 4282 16490
rect 4282 16438 4284 16490
rect 4228 16436 4284 16438
rect 4332 16490 4388 16492
rect 4332 16438 4334 16490
rect 4334 16438 4386 16490
rect 4386 16438 4388 16490
rect 4332 16436 4388 16438
rect 3612 15874 3668 15876
rect 3612 15822 3614 15874
rect 3614 15822 3666 15874
rect 3666 15822 3668 15874
rect 3612 15820 3668 15822
rect 3164 15314 3220 15316
rect 3164 15262 3166 15314
rect 3166 15262 3218 15314
rect 3218 15262 3220 15314
rect 3164 15260 3220 15262
rect 4060 15260 4116 15316
rect 4956 17052 5012 17108
rect 8204 21810 8260 21812
rect 8204 21758 8206 21810
rect 8206 21758 8258 21810
rect 8258 21758 8260 21810
rect 8204 21756 8260 21758
rect 7036 20410 7092 20412
rect 7036 20358 7038 20410
rect 7038 20358 7090 20410
rect 7090 20358 7092 20410
rect 7036 20356 7092 20358
rect 7140 20410 7196 20412
rect 7140 20358 7142 20410
rect 7142 20358 7194 20410
rect 7194 20358 7196 20410
rect 7140 20356 7196 20358
rect 7244 20410 7300 20412
rect 7244 20358 7246 20410
rect 7246 20358 7298 20410
rect 7298 20358 7300 20410
rect 7244 20356 7300 20358
rect 7868 20748 7924 20804
rect 7756 20578 7812 20580
rect 7756 20526 7758 20578
rect 7758 20526 7810 20578
rect 7810 20526 7812 20578
rect 7756 20524 7812 20526
rect 7644 20300 7700 20356
rect 6748 20242 6804 20244
rect 6748 20190 6750 20242
rect 6750 20190 6802 20242
rect 6802 20190 6804 20242
rect 6748 20188 6804 20190
rect 9660 21308 9716 21364
rect 8652 20802 8708 20804
rect 8652 20750 8654 20802
rect 8654 20750 8706 20802
rect 8706 20750 8708 20802
rect 8652 20748 8708 20750
rect 8428 20412 8484 20468
rect 8092 20188 8148 20244
rect 8316 20300 8372 20356
rect 7980 20018 8036 20020
rect 7980 19966 7982 20018
rect 7982 19966 8034 20018
rect 8034 19966 8036 20018
rect 7980 19964 8036 19966
rect 6636 19906 6692 19908
rect 6636 19854 6638 19906
rect 6638 19854 6690 19906
rect 6690 19854 6692 19906
rect 6636 19852 6692 19854
rect 6412 18284 6468 18340
rect 6748 18620 6804 18676
rect 7036 18842 7092 18844
rect 7036 18790 7038 18842
rect 7038 18790 7090 18842
rect 7090 18790 7092 18842
rect 7036 18788 7092 18790
rect 7140 18842 7196 18844
rect 7140 18790 7142 18842
rect 7142 18790 7194 18842
rect 7194 18790 7196 18842
rect 7140 18788 7196 18790
rect 7244 18842 7300 18844
rect 7244 18790 7246 18842
rect 7246 18790 7298 18842
rect 7298 18790 7300 18842
rect 7244 18788 7300 18790
rect 7308 18396 7364 18452
rect 7036 17274 7092 17276
rect 7036 17222 7038 17274
rect 7038 17222 7090 17274
rect 7090 17222 7092 17274
rect 7036 17220 7092 17222
rect 7140 17274 7196 17276
rect 7140 17222 7142 17274
rect 7142 17222 7194 17274
rect 7194 17222 7196 17274
rect 7140 17220 7196 17222
rect 7244 17274 7300 17276
rect 7244 17222 7246 17274
rect 7246 17222 7298 17274
rect 7298 17222 7300 17274
rect 7244 17220 7300 17222
rect 5740 16828 5796 16884
rect 5180 16268 5236 16324
rect 4732 15820 4788 15876
rect 4620 15372 4676 15428
rect 4396 15314 4452 15316
rect 4396 15262 4398 15314
rect 4398 15262 4450 15314
rect 4450 15262 4452 15314
rect 4396 15260 4452 15262
rect 3052 15036 3108 15092
rect 3164 14924 3220 14980
rect 2940 14476 2996 14532
rect 2716 13580 2772 13636
rect 4124 14922 4180 14924
rect 4124 14870 4126 14922
rect 4126 14870 4178 14922
rect 4178 14870 4180 14922
rect 4124 14868 4180 14870
rect 4228 14922 4284 14924
rect 4228 14870 4230 14922
rect 4230 14870 4282 14922
rect 4282 14870 4284 14922
rect 4228 14868 4284 14870
rect 4332 14922 4388 14924
rect 4332 14870 4334 14922
rect 4334 14870 4386 14922
rect 4386 14870 4388 14922
rect 4332 14868 4388 14870
rect 4396 14306 4452 14308
rect 4396 14254 4398 14306
rect 4398 14254 4450 14306
rect 4450 14254 4452 14306
rect 4396 14252 4452 14254
rect 5516 15820 5572 15876
rect 5404 15426 5460 15428
rect 5404 15374 5406 15426
rect 5406 15374 5458 15426
rect 5458 15374 5460 15426
rect 5404 15372 5460 15374
rect 5740 16658 5796 16660
rect 5740 16606 5742 16658
rect 5742 16606 5794 16658
rect 5794 16606 5796 16658
rect 5740 16604 5796 16606
rect 6748 16828 6804 16884
rect 6076 16322 6132 16324
rect 6076 16270 6078 16322
rect 6078 16270 6130 16322
rect 6130 16270 6132 16322
rect 6076 16268 6132 16270
rect 6300 16604 6356 16660
rect 5852 16098 5908 16100
rect 5852 16046 5854 16098
rect 5854 16046 5906 16098
rect 5906 16046 5908 16098
rect 5852 16044 5908 16046
rect 6524 16098 6580 16100
rect 6524 16046 6526 16098
rect 6526 16046 6578 16098
rect 6578 16046 6580 16098
rect 6524 16044 6580 16046
rect 5628 15036 5684 15092
rect 6412 14476 6468 14532
rect 4956 13916 5012 13972
rect 5292 13522 5348 13524
rect 5292 13470 5294 13522
rect 5294 13470 5346 13522
rect 5346 13470 5348 13522
rect 5292 13468 5348 13470
rect 6188 13804 6244 13860
rect 7308 15820 7364 15876
rect 7036 15706 7092 15708
rect 7036 15654 7038 15706
rect 7038 15654 7090 15706
rect 7090 15654 7092 15706
rect 7036 15652 7092 15654
rect 7140 15706 7196 15708
rect 7140 15654 7142 15706
rect 7142 15654 7194 15706
rect 7194 15654 7196 15706
rect 7140 15652 7196 15654
rect 7244 15706 7300 15708
rect 7244 15654 7246 15706
rect 7246 15654 7298 15706
rect 7298 15654 7300 15706
rect 7244 15652 7300 15654
rect 6636 15314 6692 15316
rect 6636 15262 6638 15314
rect 6638 15262 6690 15314
rect 6690 15262 6692 15314
rect 6636 15260 6692 15262
rect 6412 13746 6468 13748
rect 6412 13694 6414 13746
rect 6414 13694 6466 13746
rect 6466 13694 6468 13746
rect 6412 13692 6468 13694
rect 4124 13354 4180 13356
rect 4124 13302 4126 13354
rect 4126 13302 4178 13354
rect 4178 13302 4180 13354
rect 4124 13300 4180 13302
rect 4228 13354 4284 13356
rect 4228 13302 4230 13354
rect 4230 13302 4282 13354
rect 4282 13302 4284 13354
rect 4228 13300 4284 13302
rect 4332 13354 4388 13356
rect 4332 13302 4334 13354
rect 4334 13302 4386 13354
rect 4386 13302 4388 13354
rect 4332 13300 4388 13302
rect 6076 13468 6132 13524
rect 4124 11786 4180 11788
rect 4124 11734 4126 11786
rect 4126 11734 4178 11786
rect 4178 11734 4180 11786
rect 4124 11732 4180 11734
rect 4228 11786 4284 11788
rect 4228 11734 4230 11786
rect 4230 11734 4282 11786
rect 4282 11734 4284 11786
rect 4228 11732 4284 11734
rect 4332 11786 4388 11788
rect 4332 11734 4334 11786
rect 4334 11734 4386 11786
rect 4386 11734 4388 11786
rect 4332 11732 4388 11734
rect 3388 11452 3444 11508
rect 2044 10556 2100 10612
rect 3500 10668 3556 10724
rect 3276 10556 3332 10612
rect 3164 8818 3220 8820
rect 3164 8766 3166 8818
rect 3166 8766 3218 8818
rect 3218 8766 3220 8818
rect 3164 8764 3220 8766
rect 4124 10218 4180 10220
rect 4124 10166 4126 10218
rect 4126 10166 4178 10218
rect 4178 10166 4180 10218
rect 4124 10164 4180 10166
rect 4228 10218 4284 10220
rect 4228 10166 4230 10218
rect 4230 10166 4282 10218
rect 4282 10166 4284 10218
rect 4228 10164 4284 10166
rect 4332 10218 4388 10220
rect 4332 10166 4334 10218
rect 4334 10166 4386 10218
rect 4386 10166 4388 10218
rect 4332 10164 4388 10166
rect 3724 8316 3780 8372
rect 4620 10668 4676 10724
rect 4124 8650 4180 8652
rect 4124 8598 4126 8650
rect 4126 8598 4178 8650
rect 4178 8598 4180 8650
rect 4124 8596 4180 8598
rect 4228 8650 4284 8652
rect 4228 8598 4230 8650
rect 4230 8598 4282 8650
rect 4282 8598 4284 8650
rect 4228 8596 4284 8598
rect 4332 8650 4388 8652
rect 4332 8598 4334 8650
rect 4334 8598 4386 8650
rect 4386 8598 4388 8650
rect 4332 8596 4388 8598
rect 5964 12908 6020 12964
rect 7084 14530 7140 14532
rect 7084 14478 7086 14530
rect 7086 14478 7138 14530
rect 7138 14478 7140 14530
rect 7084 14476 7140 14478
rect 7036 14138 7092 14140
rect 7036 14086 7038 14138
rect 7038 14086 7090 14138
rect 7090 14086 7092 14138
rect 7036 14084 7092 14086
rect 7140 14138 7196 14140
rect 7140 14086 7142 14138
rect 7142 14086 7194 14138
rect 7194 14086 7196 14138
rect 7140 14084 7196 14086
rect 7244 14138 7300 14140
rect 7244 14086 7246 14138
rect 7246 14086 7298 14138
rect 7298 14086 7300 14138
rect 7244 14084 7300 14086
rect 6860 13858 6916 13860
rect 6860 13806 6862 13858
rect 6862 13806 6914 13858
rect 6914 13806 6916 13858
rect 6860 13804 6916 13806
rect 7084 13692 7140 13748
rect 6972 13580 7028 13636
rect 4844 11676 4900 11732
rect 4844 10610 4900 10612
rect 4844 10558 4846 10610
rect 4846 10558 4898 10610
rect 4898 10558 4900 10610
rect 4844 10556 4900 10558
rect 5964 11676 6020 11732
rect 5516 11452 5572 11508
rect 7036 12570 7092 12572
rect 7036 12518 7038 12570
rect 7038 12518 7090 12570
rect 7090 12518 7092 12570
rect 7036 12516 7092 12518
rect 7140 12570 7196 12572
rect 7140 12518 7142 12570
rect 7142 12518 7194 12570
rect 7194 12518 7196 12570
rect 7140 12516 7196 12518
rect 7244 12570 7300 12572
rect 7244 12518 7246 12570
rect 7246 12518 7298 12570
rect 7298 12518 7300 12570
rect 7244 12516 7300 12518
rect 6860 11452 6916 11508
rect 6860 11228 6916 11284
rect 4844 8764 4900 8820
rect 4956 7586 5012 7588
rect 4956 7534 4958 7586
rect 4958 7534 5010 7586
rect 5010 7534 5012 7586
rect 4956 7532 5012 7534
rect 4844 7474 4900 7476
rect 4844 7422 4846 7474
rect 4846 7422 4898 7474
rect 4898 7422 4900 7474
rect 4844 7420 4900 7422
rect 6412 8316 6468 8372
rect 5628 7420 5684 7476
rect 5852 7532 5908 7588
rect 4732 7196 4788 7252
rect 4124 7082 4180 7084
rect 4124 7030 4126 7082
rect 4126 7030 4178 7082
rect 4178 7030 4180 7082
rect 4124 7028 4180 7030
rect 4228 7082 4284 7084
rect 4228 7030 4230 7082
rect 4230 7030 4282 7082
rect 4282 7030 4284 7082
rect 4228 7028 4284 7030
rect 4332 7082 4388 7084
rect 4332 7030 4334 7082
rect 4334 7030 4386 7082
rect 4386 7030 4388 7082
rect 4332 7028 4388 7030
rect 5516 7250 5572 7252
rect 5516 7198 5518 7250
rect 5518 7198 5570 7250
rect 5570 7198 5572 7250
rect 5516 7196 5572 7198
rect 7036 11002 7092 11004
rect 7036 10950 7038 11002
rect 7038 10950 7090 11002
rect 7090 10950 7092 11002
rect 7036 10948 7092 10950
rect 7140 11002 7196 11004
rect 7140 10950 7142 11002
rect 7142 10950 7194 11002
rect 7194 10950 7196 11002
rect 7140 10948 7196 10950
rect 7244 11002 7300 11004
rect 7244 10950 7246 11002
rect 7246 10950 7298 11002
rect 7298 10950 7300 11002
rect 7244 10948 7300 10950
rect 7036 9434 7092 9436
rect 7036 9382 7038 9434
rect 7038 9382 7090 9434
rect 7090 9382 7092 9434
rect 7036 9380 7092 9382
rect 7140 9434 7196 9436
rect 7140 9382 7142 9434
rect 7142 9382 7194 9434
rect 7194 9382 7196 9434
rect 7140 9380 7196 9382
rect 7244 9434 7300 9436
rect 7244 9382 7246 9434
rect 7246 9382 7298 9434
rect 7298 9382 7300 9434
rect 7244 9380 7300 9382
rect 8316 19852 8372 19908
rect 8652 19122 8708 19124
rect 8652 19070 8654 19122
rect 8654 19070 8706 19122
rect 8706 19070 8708 19122
rect 8652 19068 8708 19070
rect 7756 18562 7812 18564
rect 7756 18510 7758 18562
rect 7758 18510 7810 18562
rect 7810 18510 7812 18562
rect 7756 18508 7812 18510
rect 8540 18172 8596 18228
rect 9548 19964 9604 20020
rect 9948 21194 10004 21196
rect 9948 21142 9950 21194
rect 9950 21142 10002 21194
rect 10002 21142 10004 21194
rect 9948 21140 10004 21142
rect 10052 21194 10108 21196
rect 10052 21142 10054 21194
rect 10054 21142 10106 21194
rect 10106 21142 10108 21194
rect 10052 21140 10108 21142
rect 10156 21194 10212 21196
rect 10156 21142 10158 21194
rect 10158 21142 10210 21194
rect 10210 21142 10212 21194
rect 10156 21140 10212 21142
rect 9996 20578 10052 20580
rect 9996 20526 9998 20578
rect 9998 20526 10050 20578
rect 10050 20526 10052 20578
rect 9996 20524 10052 20526
rect 10444 20412 10500 20468
rect 9884 20188 9940 20244
rect 10556 20300 10612 20356
rect 9884 19906 9940 19908
rect 9884 19854 9886 19906
rect 9886 19854 9938 19906
rect 9938 19854 9940 19906
rect 9884 19852 9940 19854
rect 9948 19626 10004 19628
rect 9948 19574 9950 19626
rect 9950 19574 10002 19626
rect 10002 19574 10004 19626
rect 9948 19572 10004 19574
rect 10052 19626 10108 19628
rect 10052 19574 10054 19626
rect 10054 19574 10106 19626
rect 10106 19574 10108 19626
rect 10052 19572 10108 19574
rect 10156 19626 10212 19628
rect 10156 19574 10158 19626
rect 10158 19574 10210 19626
rect 10210 19574 10212 19626
rect 10156 19572 10212 19574
rect 9436 19122 9492 19124
rect 9436 19070 9438 19122
rect 9438 19070 9490 19122
rect 9490 19070 9492 19122
rect 9436 19068 9492 19070
rect 9324 19010 9380 19012
rect 9324 18958 9326 19010
rect 9326 18958 9378 19010
rect 9378 18958 9380 19010
rect 9324 18956 9380 18958
rect 9772 19122 9828 19124
rect 9772 19070 9774 19122
rect 9774 19070 9826 19122
rect 9826 19070 9828 19122
rect 9772 19068 9828 19070
rect 8988 18450 9044 18452
rect 8988 18398 8990 18450
rect 8990 18398 9042 18450
rect 9042 18398 9044 18450
rect 8988 18396 9044 18398
rect 9324 17836 9380 17892
rect 9772 18396 9828 18452
rect 10780 19964 10836 20020
rect 11228 19852 11284 19908
rect 10668 19404 10724 19460
rect 10108 19122 10164 19124
rect 10108 19070 10110 19122
rect 10110 19070 10162 19122
rect 10162 19070 10164 19122
rect 10108 19068 10164 19070
rect 9884 18172 9940 18228
rect 10332 18956 10388 19012
rect 9948 18058 10004 18060
rect 9948 18006 9950 18058
rect 9950 18006 10002 18058
rect 10002 18006 10004 18058
rect 9948 18004 10004 18006
rect 10052 18058 10108 18060
rect 10052 18006 10054 18058
rect 10054 18006 10106 18058
rect 10106 18006 10108 18058
rect 10052 18004 10108 18006
rect 10156 18058 10212 18060
rect 10156 18006 10158 18058
rect 10158 18006 10210 18058
rect 10210 18006 10212 18058
rect 10156 18004 10212 18006
rect 7868 16994 7924 16996
rect 7868 16942 7870 16994
rect 7870 16942 7922 16994
rect 7922 16942 7924 16994
rect 7868 16940 7924 16942
rect 8428 16940 8484 16996
rect 7644 16044 7700 16100
rect 9660 16994 9716 16996
rect 9660 16942 9662 16994
rect 9662 16942 9714 16994
rect 9714 16942 9716 16994
rect 9660 16940 9716 16942
rect 9548 16716 9604 16772
rect 10444 16658 10500 16660
rect 10444 16606 10446 16658
rect 10446 16606 10498 16658
rect 10498 16606 10500 16658
rect 10444 16604 10500 16606
rect 9948 16490 10004 16492
rect 9948 16438 9950 16490
rect 9950 16438 10002 16490
rect 10002 16438 10004 16490
rect 9948 16436 10004 16438
rect 10052 16490 10108 16492
rect 10052 16438 10054 16490
rect 10054 16438 10106 16490
rect 10106 16438 10108 16490
rect 10052 16436 10108 16438
rect 10156 16490 10212 16492
rect 10156 16438 10158 16490
rect 10158 16438 10210 16490
rect 10210 16438 10212 16490
rect 10156 16436 10212 16438
rect 8764 16098 8820 16100
rect 8764 16046 8766 16098
rect 8766 16046 8818 16098
rect 8818 16046 8820 16098
rect 8764 16044 8820 16046
rect 7756 15036 7812 15092
rect 9660 15036 9716 15092
rect 9948 14922 10004 14924
rect 9948 14870 9950 14922
rect 9950 14870 10002 14922
rect 10002 14870 10004 14922
rect 9948 14868 10004 14870
rect 10052 14922 10108 14924
rect 10052 14870 10054 14922
rect 10054 14870 10106 14922
rect 10106 14870 10108 14922
rect 10052 14868 10108 14870
rect 10156 14922 10212 14924
rect 10156 14870 10158 14922
rect 10158 14870 10210 14922
rect 10210 14870 10212 14922
rect 10156 14868 10212 14870
rect 8428 14530 8484 14532
rect 8428 14478 8430 14530
rect 8430 14478 8482 14530
rect 8482 14478 8484 14530
rect 8428 14476 8484 14478
rect 8652 14252 8708 14308
rect 7980 13634 8036 13636
rect 7980 13582 7982 13634
rect 7982 13582 8034 13634
rect 8034 13582 8036 13634
rect 7980 13580 8036 13582
rect 8316 13634 8372 13636
rect 8316 13582 8318 13634
rect 8318 13582 8370 13634
rect 8370 13582 8372 13634
rect 8316 13580 8372 13582
rect 10892 19068 10948 19124
rect 10780 17836 10836 17892
rect 11452 19068 11508 19124
rect 11116 18674 11172 18676
rect 11116 18622 11118 18674
rect 11118 18622 11170 18674
rect 11170 18622 11172 18674
rect 11116 18620 11172 18622
rect 11788 19628 11844 19684
rect 11900 19458 11956 19460
rect 11900 19406 11902 19458
rect 11902 19406 11954 19458
rect 11954 19406 11956 19458
rect 11900 19404 11956 19406
rect 11900 19068 11956 19124
rect 12860 21978 12916 21980
rect 12860 21926 12862 21978
rect 12862 21926 12914 21978
rect 12914 21926 12916 21978
rect 12860 21924 12916 21926
rect 12964 21978 13020 21980
rect 12964 21926 12966 21978
rect 12966 21926 13018 21978
rect 13018 21926 13020 21978
rect 12964 21924 13020 21926
rect 13068 21978 13124 21980
rect 13068 21926 13070 21978
rect 13070 21926 13122 21978
rect 13122 21926 13124 21978
rect 13068 21924 13124 21926
rect 19180 22146 19236 22148
rect 19180 22094 19182 22146
rect 19182 22094 19234 22146
rect 19234 22094 19236 22146
rect 19180 22092 19236 22094
rect 18684 21978 18740 21980
rect 18684 21926 18686 21978
rect 18686 21926 18738 21978
rect 18738 21926 18740 21978
rect 18684 21924 18740 21926
rect 18788 21978 18844 21980
rect 18788 21926 18790 21978
rect 18790 21926 18842 21978
rect 18842 21926 18844 21978
rect 18788 21924 18844 21926
rect 18892 21978 18948 21980
rect 18892 21926 18894 21978
rect 18894 21926 18946 21978
rect 18946 21926 18948 21978
rect 18892 21924 18948 21926
rect 13020 21586 13076 21588
rect 13020 21534 13022 21586
rect 13022 21534 13074 21586
rect 13074 21534 13076 21586
rect 13020 21532 13076 21534
rect 12860 20410 12916 20412
rect 12860 20358 12862 20410
rect 12862 20358 12914 20410
rect 12914 20358 12916 20410
rect 12860 20356 12916 20358
rect 12964 20410 13020 20412
rect 12964 20358 12966 20410
rect 12966 20358 13018 20410
rect 13018 20358 13020 20410
rect 12964 20356 13020 20358
rect 13068 20410 13124 20412
rect 13068 20358 13070 20410
rect 13070 20358 13122 20410
rect 13122 20358 13124 20410
rect 13068 20356 13124 20358
rect 13244 20076 13300 20132
rect 14140 20130 14196 20132
rect 14140 20078 14142 20130
rect 14142 20078 14194 20130
rect 14194 20078 14196 20130
rect 14140 20076 14196 20078
rect 14924 20130 14980 20132
rect 14924 20078 14926 20130
rect 14926 20078 14978 20130
rect 14978 20078 14980 20130
rect 14924 20076 14980 20078
rect 15148 20076 15204 20132
rect 12908 19740 12964 19796
rect 13804 19740 13860 19796
rect 12348 18956 12404 19012
rect 13916 19234 13972 19236
rect 13916 19182 13918 19234
rect 13918 19182 13970 19234
rect 13970 19182 13972 19234
rect 13916 19180 13972 19182
rect 12860 18842 12916 18844
rect 12860 18790 12862 18842
rect 12862 18790 12914 18842
rect 12914 18790 12916 18842
rect 12860 18788 12916 18790
rect 12964 18842 13020 18844
rect 12964 18790 12966 18842
rect 12966 18790 13018 18842
rect 13018 18790 13020 18842
rect 12964 18788 13020 18790
rect 13068 18842 13124 18844
rect 13068 18790 13070 18842
rect 13070 18790 13122 18842
rect 13122 18790 13124 18842
rect 13068 18788 13124 18790
rect 12012 18620 12068 18676
rect 11340 17836 11396 17892
rect 12236 18396 12292 18452
rect 12572 18284 12628 18340
rect 12908 18450 12964 18452
rect 12908 18398 12910 18450
rect 12910 18398 12962 18450
rect 12962 18398 12964 18450
rect 12908 18396 12964 18398
rect 12908 17500 12964 17556
rect 11004 17052 11060 17108
rect 11004 16716 11060 16772
rect 11788 16770 11844 16772
rect 11788 16718 11790 16770
rect 11790 16718 11842 16770
rect 11842 16718 11844 16770
rect 11788 16716 11844 16718
rect 15708 21532 15764 21588
rect 17500 21698 17556 21700
rect 17500 21646 17502 21698
rect 17502 21646 17554 21698
rect 17554 21646 17556 21698
rect 17500 21644 17556 21646
rect 16268 21586 16324 21588
rect 16268 21534 16270 21586
rect 16270 21534 16322 21586
rect 16322 21534 16324 21586
rect 16268 21532 16324 21534
rect 16492 21308 16548 21364
rect 15772 21194 15828 21196
rect 15772 21142 15774 21194
rect 15774 21142 15826 21194
rect 15826 21142 15828 21194
rect 15772 21140 15828 21142
rect 15876 21194 15932 21196
rect 15876 21142 15878 21194
rect 15878 21142 15930 21194
rect 15930 21142 15932 21194
rect 15876 21140 15932 21142
rect 15980 21194 16036 21196
rect 15980 21142 15982 21194
rect 15982 21142 16034 21194
rect 16034 21142 16036 21194
rect 15980 21140 16036 21142
rect 16604 20130 16660 20132
rect 16604 20078 16606 20130
rect 16606 20078 16658 20130
rect 16658 20078 16660 20130
rect 16604 20076 16660 20078
rect 17948 21586 18004 21588
rect 17948 21534 17950 21586
rect 17950 21534 18002 21586
rect 18002 21534 18004 21586
rect 17948 21532 18004 21534
rect 17500 21362 17556 21364
rect 17500 21310 17502 21362
rect 17502 21310 17554 21362
rect 17554 21310 17556 21362
rect 17500 21308 17556 21310
rect 17276 20076 17332 20132
rect 16044 19740 16100 19796
rect 15772 19626 15828 19628
rect 15772 19574 15774 19626
rect 15774 19574 15826 19626
rect 15826 19574 15828 19626
rect 15772 19572 15828 19574
rect 15876 19626 15932 19628
rect 15876 19574 15878 19626
rect 15878 19574 15930 19626
rect 15930 19574 15932 19626
rect 15876 19572 15932 19574
rect 15980 19626 16036 19628
rect 15980 19574 15982 19626
rect 15982 19574 16034 19626
rect 16034 19574 16036 19626
rect 15980 19572 16036 19574
rect 14364 19234 14420 19236
rect 14364 19182 14366 19234
rect 14366 19182 14418 19234
rect 14418 19182 14420 19234
rect 14364 19180 14420 19182
rect 14588 19234 14644 19236
rect 14588 19182 14590 19234
rect 14590 19182 14642 19234
rect 14642 19182 14644 19234
rect 14588 19180 14644 19182
rect 14476 19010 14532 19012
rect 14476 18958 14478 19010
rect 14478 18958 14530 19010
rect 14530 18958 14532 19010
rect 14476 18956 14532 18958
rect 14812 18956 14868 19012
rect 14364 18674 14420 18676
rect 14364 18622 14366 18674
rect 14366 18622 14418 18674
rect 14418 18622 14420 18674
rect 14364 18620 14420 18622
rect 14140 18396 14196 18452
rect 14812 18284 14868 18340
rect 15372 19234 15428 19236
rect 15372 19182 15374 19234
rect 15374 19182 15426 19234
rect 15426 19182 15428 19234
rect 15372 19180 15428 19182
rect 15260 18956 15316 19012
rect 15148 18620 15204 18676
rect 15148 18450 15204 18452
rect 15148 18398 15150 18450
rect 15150 18398 15202 18450
rect 15202 18398 15204 18450
rect 15148 18396 15204 18398
rect 15260 18284 15316 18340
rect 15484 18396 15540 18452
rect 12860 17274 12916 17276
rect 12860 17222 12862 17274
rect 12862 17222 12914 17274
rect 12914 17222 12916 17274
rect 12860 17220 12916 17222
rect 12964 17274 13020 17276
rect 12964 17222 12966 17274
rect 12966 17222 13018 17274
rect 13018 17222 13020 17274
rect 12964 17220 13020 17222
rect 13068 17274 13124 17276
rect 13068 17222 13070 17274
rect 13070 17222 13122 17274
rect 13122 17222 13124 17274
rect 13916 17276 13972 17332
rect 13068 17220 13124 17222
rect 13580 16716 13636 16772
rect 11900 16604 11956 16660
rect 13468 16604 13524 16660
rect 14476 16268 14532 16324
rect 12860 15706 12916 15708
rect 12860 15654 12862 15706
rect 12862 15654 12914 15706
rect 12914 15654 12916 15706
rect 12860 15652 12916 15654
rect 12964 15706 13020 15708
rect 12964 15654 12966 15706
rect 12966 15654 13018 15706
rect 13018 15654 13020 15706
rect 12964 15652 13020 15654
rect 13068 15706 13124 15708
rect 13068 15654 13070 15706
rect 13070 15654 13122 15706
rect 13122 15654 13124 15706
rect 13068 15652 13124 15654
rect 11900 15148 11956 15204
rect 11228 13746 11284 13748
rect 11228 13694 11230 13746
rect 11230 13694 11282 13746
rect 11282 13694 11284 13746
rect 11228 13692 11284 13694
rect 9548 13580 9604 13636
rect 9948 13354 10004 13356
rect 9948 13302 9950 13354
rect 9950 13302 10002 13354
rect 10002 13302 10004 13354
rect 9948 13300 10004 13302
rect 10052 13354 10108 13356
rect 10052 13302 10054 13354
rect 10054 13302 10106 13354
rect 10106 13302 10108 13354
rect 10052 13300 10108 13302
rect 10156 13354 10212 13356
rect 10156 13302 10158 13354
rect 10158 13302 10210 13354
rect 10210 13302 10212 13354
rect 10156 13300 10212 13302
rect 7868 12962 7924 12964
rect 7868 12910 7870 12962
rect 7870 12910 7922 12962
rect 7922 12910 7924 12962
rect 7868 12908 7924 12910
rect 7868 11228 7924 11284
rect 9948 11786 10004 11788
rect 9948 11734 9950 11786
rect 9950 11734 10002 11786
rect 10002 11734 10004 11786
rect 9948 11732 10004 11734
rect 10052 11786 10108 11788
rect 10052 11734 10054 11786
rect 10054 11734 10106 11786
rect 10106 11734 10108 11786
rect 10052 11732 10108 11734
rect 10156 11786 10212 11788
rect 10156 11734 10158 11786
rect 10158 11734 10210 11786
rect 10210 11734 10212 11786
rect 10156 11732 10212 11734
rect 8764 10556 8820 10612
rect 9324 11282 9380 11284
rect 9324 11230 9326 11282
rect 9326 11230 9378 11282
rect 9378 11230 9380 11282
rect 9324 11228 9380 11230
rect 7420 9324 7476 9380
rect 7196 9212 7252 9268
rect 6636 7586 6692 7588
rect 6636 7534 6638 7586
rect 6638 7534 6690 7586
rect 6690 7534 6692 7586
rect 6636 7532 6692 7534
rect 4124 5514 4180 5516
rect 4124 5462 4126 5514
rect 4126 5462 4178 5514
rect 4178 5462 4180 5514
rect 4124 5460 4180 5462
rect 4228 5514 4284 5516
rect 4228 5462 4230 5514
rect 4230 5462 4282 5514
rect 4282 5462 4284 5514
rect 4228 5460 4284 5462
rect 4332 5514 4388 5516
rect 4332 5462 4334 5514
rect 4334 5462 4386 5514
rect 4386 5462 4388 5514
rect 4332 5460 4388 5462
rect 7036 7866 7092 7868
rect 7036 7814 7038 7866
rect 7038 7814 7090 7866
rect 7090 7814 7092 7866
rect 7036 7812 7092 7814
rect 7140 7866 7196 7868
rect 7140 7814 7142 7866
rect 7142 7814 7194 7866
rect 7194 7814 7196 7866
rect 7140 7812 7196 7814
rect 7244 7866 7300 7868
rect 7244 7814 7246 7866
rect 7246 7814 7298 7866
rect 7298 7814 7300 7866
rect 7244 7812 7300 7814
rect 7196 7586 7252 7588
rect 7196 7534 7198 7586
rect 7198 7534 7250 7586
rect 7250 7534 7252 7586
rect 7196 7532 7252 7534
rect 9772 10722 9828 10724
rect 9772 10670 9774 10722
rect 9774 10670 9826 10722
rect 9826 10670 9828 10722
rect 9772 10668 9828 10670
rect 10220 10722 10276 10724
rect 10220 10670 10222 10722
rect 10222 10670 10274 10722
rect 10274 10670 10276 10722
rect 10220 10668 10276 10670
rect 9948 10218 10004 10220
rect 9948 10166 9950 10218
rect 9950 10166 10002 10218
rect 10002 10166 10004 10218
rect 9948 10164 10004 10166
rect 10052 10218 10108 10220
rect 10052 10166 10054 10218
rect 10054 10166 10106 10218
rect 10106 10166 10108 10218
rect 10052 10164 10108 10166
rect 10156 10218 10212 10220
rect 10156 10166 10158 10218
rect 10158 10166 10210 10218
rect 10210 10166 10212 10218
rect 10156 10164 10212 10166
rect 10668 12290 10724 12292
rect 10668 12238 10670 12290
rect 10670 12238 10722 12290
rect 10722 12238 10724 12290
rect 10668 12236 10724 12238
rect 11676 12178 11732 12180
rect 11676 12126 11678 12178
rect 11678 12126 11730 12178
rect 11730 12126 11732 12178
rect 11676 12124 11732 12126
rect 12348 15036 12404 15092
rect 12908 14642 12964 14644
rect 12908 14590 12910 14642
rect 12910 14590 12962 14642
rect 12962 14590 12964 14642
rect 12908 14588 12964 14590
rect 12460 13692 12516 13748
rect 12860 14138 12916 14140
rect 12860 14086 12862 14138
rect 12862 14086 12914 14138
rect 12914 14086 12916 14138
rect 12860 14084 12916 14086
rect 12964 14138 13020 14140
rect 12964 14086 12966 14138
rect 12966 14086 13018 14138
rect 13018 14086 13020 14138
rect 12964 14084 13020 14086
rect 13068 14138 13124 14140
rect 13068 14086 13070 14138
rect 13070 14086 13122 14138
rect 13122 14086 13124 14138
rect 13068 14084 13124 14086
rect 16716 19740 16772 19796
rect 16492 19628 16548 19684
rect 16268 18396 16324 18452
rect 16156 18284 16212 18340
rect 15772 18058 15828 18060
rect 15772 18006 15774 18058
rect 15774 18006 15826 18058
rect 15826 18006 15828 18058
rect 15772 18004 15828 18006
rect 15876 18058 15932 18060
rect 15876 18006 15878 18058
rect 15878 18006 15930 18058
rect 15930 18006 15932 18058
rect 15876 18004 15932 18006
rect 15980 18058 16036 18060
rect 15980 18006 15982 18058
rect 15982 18006 16034 18058
rect 16034 18006 16036 18058
rect 15980 18004 16036 18006
rect 16380 18172 16436 18228
rect 16828 19628 16884 19684
rect 16940 19234 16996 19236
rect 16940 19182 16942 19234
rect 16942 19182 16994 19234
rect 16994 19182 16996 19234
rect 16940 19180 16996 19182
rect 18396 21532 18452 21588
rect 18508 21644 18564 21700
rect 20860 22092 20916 22148
rect 21084 21868 21140 21924
rect 24508 21978 24564 21980
rect 21420 21644 21476 21700
rect 23660 21868 23716 21924
rect 24508 21926 24510 21978
rect 24510 21926 24562 21978
rect 24562 21926 24564 21978
rect 24508 21924 24564 21926
rect 24612 21978 24668 21980
rect 24612 21926 24614 21978
rect 24614 21926 24666 21978
rect 24666 21926 24668 21978
rect 24612 21924 24668 21926
rect 24716 21978 24772 21980
rect 24716 21926 24718 21978
rect 24718 21926 24770 21978
rect 24770 21926 24772 21978
rect 24716 21924 24772 21926
rect 20188 21532 20244 21588
rect 18732 21474 18788 21476
rect 18732 21422 18734 21474
rect 18734 21422 18786 21474
rect 18786 21422 18788 21474
rect 18732 21420 18788 21422
rect 20412 21420 20468 21476
rect 19516 20802 19572 20804
rect 19516 20750 19518 20802
rect 19518 20750 19570 20802
rect 19570 20750 19572 20802
rect 19516 20748 19572 20750
rect 18684 20410 18740 20412
rect 18684 20358 18686 20410
rect 18686 20358 18738 20410
rect 18738 20358 18740 20410
rect 18684 20356 18740 20358
rect 18788 20410 18844 20412
rect 18788 20358 18790 20410
rect 18790 20358 18842 20410
rect 18842 20358 18844 20410
rect 18788 20356 18844 20358
rect 18892 20410 18948 20412
rect 18892 20358 18894 20410
rect 18894 20358 18946 20410
rect 18946 20358 18948 20410
rect 18892 20356 18948 20358
rect 17948 20076 18004 20132
rect 18732 20130 18788 20132
rect 18732 20078 18734 20130
rect 18734 20078 18786 20130
rect 18786 20078 18788 20130
rect 18732 20076 18788 20078
rect 19404 20130 19460 20132
rect 19404 20078 19406 20130
rect 19406 20078 19458 20130
rect 19458 20078 19460 20130
rect 19404 20076 19460 20078
rect 17836 19794 17892 19796
rect 17836 19742 17838 19794
rect 17838 19742 17890 19794
rect 17890 19742 17892 19794
rect 17836 19740 17892 19742
rect 18172 19404 18228 19460
rect 20860 20748 20916 20804
rect 20636 20636 20692 20692
rect 20412 20524 20468 20580
rect 19852 19292 19908 19348
rect 19964 19740 20020 19796
rect 19628 19180 19684 19236
rect 16604 19010 16660 19012
rect 16604 18958 16606 19010
rect 16606 18958 16658 19010
rect 16658 18958 16660 19010
rect 16604 18956 16660 18958
rect 18684 18842 18740 18844
rect 18684 18790 18686 18842
rect 18686 18790 18738 18842
rect 18738 18790 18740 18842
rect 18684 18788 18740 18790
rect 18788 18842 18844 18844
rect 18788 18790 18790 18842
rect 18790 18790 18842 18842
rect 18842 18790 18844 18842
rect 18788 18788 18844 18790
rect 18892 18842 18948 18844
rect 18892 18790 18894 18842
rect 18894 18790 18946 18842
rect 18946 18790 18948 18842
rect 18892 18788 18948 18790
rect 17388 18396 17444 18452
rect 15484 16604 15540 16660
rect 16828 18284 16884 18340
rect 16268 17276 16324 17332
rect 16156 16940 16212 16996
rect 16492 16940 16548 16996
rect 14812 16268 14868 16324
rect 14924 16044 14980 16100
rect 14700 15932 14756 15988
rect 14476 15372 14532 15428
rect 14364 15148 14420 15204
rect 15036 15932 15092 15988
rect 14924 15596 14980 15652
rect 14140 13692 14196 13748
rect 12860 12570 12916 12572
rect 12860 12518 12862 12570
rect 12862 12518 12914 12570
rect 12914 12518 12916 12570
rect 12860 12516 12916 12518
rect 12964 12570 13020 12572
rect 12964 12518 12966 12570
rect 12966 12518 13018 12570
rect 13018 12518 13020 12570
rect 12964 12516 13020 12518
rect 13068 12570 13124 12572
rect 13068 12518 13070 12570
rect 13070 12518 13122 12570
rect 13122 12518 13124 12570
rect 13068 12516 13124 12518
rect 14252 12348 14308 12404
rect 12684 12236 12740 12292
rect 11228 11564 11284 11620
rect 11452 11394 11508 11396
rect 11452 11342 11454 11394
rect 11454 11342 11506 11394
rect 11506 11342 11508 11394
rect 11452 11340 11508 11342
rect 10668 10668 10724 10724
rect 11340 11228 11396 11284
rect 10444 10610 10500 10612
rect 10444 10558 10446 10610
rect 10446 10558 10498 10610
rect 10498 10558 10500 10610
rect 10444 10556 10500 10558
rect 10332 9996 10388 10052
rect 9948 8650 10004 8652
rect 9948 8598 9950 8650
rect 9950 8598 10002 8650
rect 10002 8598 10004 8650
rect 9948 8596 10004 8598
rect 10052 8650 10108 8652
rect 10052 8598 10054 8650
rect 10054 8598 10106 8650
rect 10106 8598 10108 8650
rect 10052 8596 10108 8598
rect 10156 8650 10212 8652
rect 10156 8598 10158 8650
rect 10158 8598 10210 8650
rect 10210 8598 10212 8650
rect 10156 8596 10212 8598
rect 8316 7586 8372 7588
rect 8316 7534 8318 7586
rect 8318 7534 8370 7586
rect 8370 7534 8372 7586
rect 8316 7532 8372 7534
rect 9212 7532 9268 7588
rect 7756 7420 7812 7476
rect 10332 8316 10388 8372
rect 10444 7756 10500 7812
rect 9660 7420 9716 7476
rect 10332 7474 10388 7476
rect 10332 7422 10334 7474
rect 10334 7422 10386 7474
rect 10386 7422 10388 7474
rect 10332 7420 10388 7422
rect 8316 6690 8372 6692
rect 8316 6638 8318 6690
rect 8318 6638 8370 6690
rect 8370 6638 8372 6690
rect 8316 6636 8372 6638
rect 8876 6690 8932 6692
rect 8876 6638 8878 6690
rect 8878 6638 8930 6690
rect 8930 6638 8932 6690
rect 8876 6636 8932 6638
rect 7036 6298 7092 6300
rect 7036 6246 7038 6298
rect 7038 6246 7090 6298
rect 7090 6246 7092 6298
rect 7036 6244 7092 6246
rect 7140 6298 7196 6300
rect 7140 6246 7142 6298
rect 7142 6246 7194 6298
rect 7194 6246 7196 6298
rect 7140 6244 7196 6246
rect 7244 6298 7300 6300
rect 7244 6246 7246 6298
rect 7246 6246 7298 6298
rect 7298 6246 7300 6298
rect 7244 6244 7300 6246
rect 9948 7082 10004 7084
rect 9948 7030 9950 7082
rect 9950 7030 10002 7082
rect 10002 7030 10004 7082
rect 9948 7028 10004 7030
rect 10052 7082 10108 7084
rect 10052 7030 10054 7082
rect 10054 7030 10106 7082
rect 10106 7030 10108 7082
rect 10052 7028 10108 7030
rect 10156 7082 10212 7084
rect 10156 7030 10158 7082
rect 10158 7030 10210 7082
rect 10210 7030 10212 7082
rect 10156 7028 10212 7030
rect 12012 9996 12068 10052
rect 14252 12012 14308 12068
rect 12684 11282 12740 11284
rect 12684 11230 12686 11282
rect 12686 11230 12738 11282
rect 12738 11230 12740 11282
rect 12684 11228 12740 11230
rect 13580 11282 13636 11284
rect 13580 11230 13582 11282
rect 13582 11230 13634 11282
rect 13634 11230 13636 11282
rect 13580 11228 13636 11230
rect 12860 11002 12916 11004
rect 12860 10950 12862 11002
rect 12862 10950 12914 11002
rect 12914 10950 12916 11002
rect 12860 10948 12916 10950
rect 12964 11002 13020 11004
rect 12964 10950 12966 11002
rect 12966 10950 13018 11002
rect 13018 10950 13020 11002
rect 12964 10948 13020 10950
rect 13068 11002 13124 11004
rect 13068 10950 13070 11002
rect 13070 10950 13122 11002
rect 13122 10950 13124 11002
rect 13068 10948 13124 10950
rect 15772 16490 15828 16492
rect 15772 16438 15774 16490
rect 15774 16438 15826 16490
rect 15826 16438 15828 16490
rect 15772 16436 15828 16438
rect 15876 16490 15932 16492
rect 15876 16438 15878 16490
rect 15878 16438 15930 16490
rect 15930 16438 15932 16490
rect 15876 16436 15932 16438
rect 15980 16490 16036 16492
rect 15980 16438 15982 16490
rect 15982 16438 16034 16490
rect 16034 16438 16036 16490
rect 15980 16436 16036 16438
rect 15596 15986 15652 15988
rect 15596 15934 15598 15986
rect 15598 15934 15650 15986
rect 15650 15934 15652 15986
rect 15596 15932 15652 15934
rect 15148 15484 15204 15540
rect 15484 15426 15540 15428
rect 15484 15374 15486 15426
rect 15486 15374 15538 15426
rect 15538 15374 15540 15426
rect 15484 15372 15540 15374
rect 15596 15260 15652 15316
rect 15260 15148 15316 15204
rect 15708 15036 15764 15092
rect 15772 14922 15828 14924
rect 15772 14870 15774 14922
rect 15774 14870 15826 14922
rect 15826 14870 15828 14922
rect 15772 14868 15828 14870
rect 15876 14922 15932 14924
rect 15876 14870 15878 14922
rect 15878 14870 15930 14922
rect 15930 14870 15932 14922
rect 15876 14868 15932 14870
rect 15980 14922 16036 14924
rect 15980 14870 15982 14922
rect 15982 14870 16034 14922
rect 16034 14870 16036 14922
rect 15980 14868 16036 14870
rect 16604 15372 16660 15428
rect 16492 15314 16548 15316
rect 16492 15262 16494 15314
rect 16494 15262 16546 15314
rect 16546 15262 16548 15314
rect 16492 15260 16548 15262
rect 16380 15036 16436 15092
rect 16492 14924 16548 14980
rect 16492 14588 16548 14644
rect 14812 12124 14868 12180
rect 14700 11788 14756 11844
rect 14476 11564 14532 11620
rect 15772 13354 15828 13356
rect 15772 13302 15774 13354
rect 15774 13302 15826 13354
rect 15826 13302 15828 13354
rect 15772 13300 15828 13302
rect 15876 13354 15932 13356
rect 15876 13302 15878 13354
rect 15878 13302 15930 13354
rect 15930 13302 15932 13354
rect 15876 13300 15932 13302
rect 15980 13354 16036 13356
rect 15980 13302 15982 13354
rect 15982 13302 16034 13354
rect 16034 13302 16036 13354
rect 15980 13300 16036 13302
rect 15484 12402 15540 12404
rect 15484 12350 15486 12402
rect 15486 12350 15538 12402
rect 15538 12350 15540 12402
rect 15484 12348 15540 12350
rect 15596 12236 15652 12292
rect 15036 12012 15092 12068
rect 14924 11340 14980 11396
rect 15372 12066 15428 12068
rect 15372 12014 15374 12066
rect 15374 12014 15426 12066
rect 15426 12014 15428 12066
rect 15372 12012 15428 12014
rect 15596 11788 15652 11844
rect 17612 18172 17668 18228
rect 17164 17666 17220 17668
rect 17164 17614 17166 17666
rect 17166 17614 17218 17666
rect 17218 17614 17220 17666
rect 17164 17612 17220 17614
rect 18060 17666 18116 17668
rect 18060 17614 18062 17666
rect 18062 17614 18114 17666
rect 18114 17614 18116 17666
rect 18060 17612 18116 17614
rect 19180 17666 19236 17668
rect 19180 17614 19182 17666
rect 19182 17614 19234 17666
rect 19234 17614 19236 17666
rect 19180 17612 19236 17614
rect 16940 17554 16996 17556
rect 16940 17502 16942 17554
rect 16942 17502 16994 17554
rect 16994 17502 16996 17554
rect 16940 17500 16996 17502
rect 16716 15036 16772 15092
rect 17276 16156 17332 16212
rect 18060 15986 18116 15988
rect 18060 15934 18062 15986
rect 18062 15934 18114 15986
rect 18114 15934 18116 15986
rect 18060 15932 18116 15934
rect 17388 15596 17444 15652
rect 17388 15426 17444 15428
rect 17388 15374 17390 15426
rect 17390 15374 17442 15426
rect 17442 15374 17444 15426
rect 17388 15372 17444 15374
rect 17612 15314 17668 15316
rect 17612 15262 17614 15314
rect 17614 15262 17666 15314
rect 17666 15262 17668 15314
rect 17612 15260 17668 15262
rect 18684 17274 18740 17276
rect 18684 17222 18686 17274
rect 18686 17222 18738 17274
rect 18738 17222 18740 17274
rect 18684 17220 18740 17222
rect 18788 17274 18844 17276
rect 18788 17222 18790 17274
rect 18790 17222 18842 17274
rect 18842 17222 18844 17274
rect 18788 17220 18844 17222
rect 18892 17274 18948 17276
rect 18892 17222 18894 17274
rect 18894 17222 18946 17274
rect 18946 17222 18948 17274
rect 18892 17220 18948 17222
rect 20524 20076 20580 20132
rect 20076 19346 20132 19348
rect 20076 19294 20078 19346
rect 20078 19294 20130 19346
rect 20130 19294 20132 19346
rect 20076 19292 20132 19294
rect 20860 20188 20916 20244
rect 23548 21532 23604 21588
rect 21596 21194 21652 21196
rect 21596 21142 21598 21194
rect 21598 21142 21650 21194
rect 21650 21142 21652 21194
rect 21596 21140 21652 21142
rect 21700 21194 21756 21196
rect 21700 21142 21702 21194
rect 21702 21142 21754 21194
rect 21754 21142 21756 21194
rect 21700 21140 21756 21142
rect 21804 21194 21860 21196
rect 21804 21142 21806 21194
rect 21806 21142 21858 21194
rect 21858 21142 21860 21194
rect 21804 21140 21860 21142
rect 21756 20690 21812 20692
rect 21756 20638 21758 20690
rect 21758 20638 21810 20690
rect 21810 20638 21812 20690
rect 21756 20636 21812 20638
rect 21196 20076 21252 20132
rect 21084 20018 21140 20020
rect 21084 19966 21086 20018
rect 21086 19966 21138 20018
rect 21138 19966 21140 20018
rect 21084 19964 21140 19966
rect 19292 16492 19348 16548
rect 18684 15706 18740 15708
rect 18684 15654 18686 15706
rect 18686 15654 18738 15706
rect 18738 15654 18740 15706
rect 18684 15652 18740 15654
rect 18788 15706 18844 15708
rect 18788 15654 18790 15706
rect 18790 15654 18842 15706
rect 18842 15654 18844 15706
rect 18788 15652 18844 15654
rect 18892 15706 18948 15708
rect 18892 15654 18894 15706
rect 18894 15654 18946 15706
rect 18946 15654 18948 15706
rect 18892 15652 18948 15654
rect 20076 18956 20132 19012
rect 20636 18396 20692 18452
rect 20412 18338 20468 18340
rect 20412 18286 20414 18338
rect 20414 18286 20466 18338
rect 20466 18286 20468 18338
rect 20412 18284 20468 18286
rect 19516 17442 19572 17444
rect 19516 17390 19518 17442
rect 19518 17390 19570 17442
rect 19570 17390 19572 17442
rect 19516 17388 19572 17390
rect 20524 18172 20580 18228
rect 20300 17612 20356 17668
rect 20188 16492 20244 16548
rect 19628 16044 19684 16100
rect 20076 15932 20132 15988
rect 19404 15260 19460 15316
rect 20748 17778 20804 17780
rect 20748 17726 20750 17778
rect 20750 17726 20802 17778
rect 20802 17726 20804 17778
rect 20748 17724 20804 17726
rect 20636 16210 20692 16212
rect 20636 16158 20638 16210
rect 20638 16158 20690 16210
rect 20690 16158 20692 16210
rect 20636 16156 20692 16158
rect 20524 15314 20580 15316
rect 20524 15262 20526 15314
rect 20526 15262 20578 15314
rect 20578 15262 20580 15314
rect 20524 15260 20580 15262
rect 15772 11786 15828 11788
rect 15772 11734 15774 11786
rect 15774 11734 15826 11786
rect 15826 11734 15828 11786
rect 15772 11732 15828 11734
rect 15876 11786 15932 11788
rect 15876 11734 15878 11786
rect 15878 11734 15930 11786
rect 15930 11734 15932 11786
rect 15876 11732 15932 11734
rect 15980 11786 16036 11788
rect 15980 11734 15982 11786
rect 15982 11734 16034 11786
rect 16034 11734 16036 11786
rect 15980 11732 16036 11734
rect 15484 11394 15540 11396
rect 15484 11342 15486 11394
rect 15486 11342 15538 11394
rect 15538 11342 15540 11394
rect 15484 11340 15540 11342
rect 16716 13020 16772 13076
rect 16380 12290 16436 12292
rect 16380 12238 16382 12290
rect 16382 12238 16434 12290
rect 16434 12238 16436 12290
rect 16380 12236 16436 12238
rect 17388 13970 17444 13972
rect 17388 13918 17390 13970
rect 17390 13918 17442 13970
rect 17442 13918 17444 13970
rect 17388 13916 17444 13918
rect 16940 12124 16996 12180
rect 16828 12066 16884 12068
rect 16828 12014 16830 12066
rect 16830 12014 16882 12066
rect 16882 12014 16884 12066
rect 16828 12012 16884 12014
rect 18284 13074 18340 13076
rect 18284 13022 18286 13074
rect 18286 13022 18338 13074
rect 18338 13022 18340 13074
rect 18284 13020 18340 13022
rect 18684 14138 18740 14140
rect 18684 14086 18686 14138
rect 18686 14086 18738 14138
rect 18738 14086 18740 14138
rect 18684 14084 18740 14086
rect 18788 14138 18844 14140
rect 18788 14086 18790 14138
rect 18790 14086 18842 14138
rect 18842 14086 18844 14138
rect 18788 14084 18844 14086
rect 18892 14138 18948 14140
rect 18892 14086 18894 14138
rect 18894 14086 18946 14138
rect 18946 14086 18948 14138
rect 18892 14084 18948 14086
rect 17500 12348 17556 12404
rect 18396 12796 18452 12852
rect 12860 9434 12916 9436
rect 12860 9382 12862 9434
rect 12862 9382 12914 9434
rect 12914 9382 12916 9434
rect 12860 9380 12916 9382
rect 12964 9434 13020 9436
rect 12964 9382 12966 9434
rect 12966 9382 13018 9434
rect 13018 9382 13020 9434
rect 12964 9380 13020 9382
rect 13068 9434 13124 9436
rect 13068 9382 13070 9434
rect 13070 9382 13122 9434
rect 13122 9382 13124 9434
rect 13068 9380 13124 9382
rect 14812 9324 14868 9380
rect 12572 8988 12628 9044
rect 10556 7644 10612 7700
rect 15372 8988 15428 9044
rect 15484 8876 15540 8932
rect 11116 7586 11172 7588
rect 11116 7534 11118 7586
rect 11118 7534 11170 7586
rect 11170 7534 11172 7586
rect 11116 7532 11172 7534
rect 11004 7308 11060 7364
rect 12012 7532 12068 7588
rect 12860 7866 12916 7868
rect 12860 7814 12862 7866
rect 12862 7814 12914 7866
rect 12914 7814 12916 7866
rect 12860 7812 12916 7814
rect 12964 7866 13020 7868
rect 12964 7814 12966 7866
rect 12966 7814 13018 7866
rect 13018 7814 13020 7866
rect 12964 7812 13020 7814
rect 13068 7866 13124 7868
rect 13068 7814 13070 7866
rect 13070 7814 13122 7866
rect 13122 7814 13124 7866
rect 13068 7812 13124 7814
rect 12796 7532 12852 7588
rect 15772 10218 15828 10220
rect 15772 10166 15774 10218
rect 15774 10166 15826 10218
rect 15826 10166 15828 10218
rect 15772 10164 15828 10166
rect 15876 10218 15932 10220
rect 15876 10166 15878 10218
rect 15878 10166 15930 10218
rect 15930 10166 15932 10218
rect 15876 10164 15932 10166
rect 15980 10218 16036 10220
rect 15980 10166 15982 10218
rect 15982 10166 16034 10218
rect 16034 10166 16036 10218
rect 15980 10164 16036 10166
rect 17388 10108 17444 10164
rect 16380 9266 16436 9268
rect 16380 9214 16382 9266
rect 16382 9214 16434 9266
rect 16434 9214 16436 9266
rect 16380 9212 16436 9214
rect 15820 9042 15876 9044
rect 15820 8990 15822 9042
rect 15822 8990 15874 9042
rect 15874 8990 15876 9042
rect 15820 8988 15876 8990
rect 15772 8650 15828 8652
rect 15772 8598 15774 8650
rect 15774 8598 15826 8650
rect 15826 8598 15828 8650
rect 15772 8596 15828 8598
rect 15876 8650 15932 8652
rect 15876 8598 15878 8650
rect 15878 8598 15930 8650
rect 15930 8598 15932 8650
rect 15876 8596 15932 8598
rect 15980 8650 16036 8652
rect 15980 8598 15982 8650
rect 15982 8598 16034 8650
rect 16034 8598 16036 8650
rect 15980 8596 16036 8598
rect 15596 7532 15652 7588
rect 13916 7362 13972 7364
rect 13916 7310 13918 7362
rect 13918 7310 13970 7362
rect 13970 7310 13972 7362
rect 13916 7308 13972 7310
rect 18172 9660 18228 9716
rect 18684 12570 18740 12572
rect 18684 12518 18686 12570
rect 18686 12518 18738 12570
rect 18738 12518 18740 12570
rect 18684 12516 18740 12518
rect 18788 12570 18844 12572
rect 18788 12518 18790 12570
rect 18790 12518 18842 12570
rect 18842 12518 18844 12570
rect 18788 12516 18844 12518
rect 18892 12570 18948 12572
rect 18892 12518 18894 12570
rect 18894 12518 18946 12570
rect 18946 12518 18948 12570
rect 18892 12516 18948 12518
rect 19292 12402 19348 12404
rect 19292 12350 19294 12402
rect 19294 12350 19346 12402
rect 19346 12350 19348 12402
rect 19292 12348 19348 12350
rect 19964 13746 20020 13748
rect 19964 13694 19966 13746
rect 19966 13694 20018 13746
rect 20018 13694 20020 13746
rect 19964 13692 20020 13694
rect 20300 13692 20356 13748
rect 21868 20524 21924 20580
rect 21868 20188 21924 20244
rect 21532 19964 21588 20020
rect 22428 20802 22484 20804
rect 22428 20750 22430 20802
rect 22430 20750 22482 20802
rect 22482 20750 22484 20802
rect 22428 20748 22484 20750
rect 23212 20802 23268 20804
rect 23212 20750 23214 20802
rect 23214 20750 23266 20802
rect 23266 20750 23268 20802
rect 23212 20748 23268 20750
rect 23212 20188 23268 20244
rect 21644 19740 21700 19796
rect 21596 19626 21652 19628
rect 21596 19574 21598 19626
rect 21598 19574 21650 19626
rect 21650 19574 21652 19626
rect 21596 19572 21652 19574
rect 21700 19626 21756 19628
rect 21700 19574 21702 19626
rect 21702 19574 21754 19626
rect 21754 19574 21756 19626
rect 21700 19572 21756 19574
rect 21804 19626 21860 19628
rect 21804 19574 21806 19626
rect 21806 19574 21858 19626
rect 21858 19574 21860 19626
rect 21804 19572 21860 19574
rect 21420 19404 21476 19460
rect 21644 19458 21700 19460
rect 21644 19406 21646 19458
rect 21646 19406 21698 19458
rect 21698 19406 21700 19458
rect 21644 19404 21700 19406
rect 21532 19292 21588 19348
rect 21308 19180 21364 19236
rect 22092 19292 22148 19348
rect 20748 17388 20804 17444
rect 21532 18172 21588 18228
rect 20412 13356 20468 13412
rect 20524 13468 20580 13524
rect 21308 16492 21364 16548
rect 22092 19010 22148 19012
rect 22092 18958 22094 19010
rect 22094 18958 22146 19010
rect 22146 18958 22148 19010
rect 22092 18956 22148 18958
rect 21868 18172 21924 18228
rect 21596 18058 21652 18060
rect 21596 18006 21598 18058
rect 21598 18006 21650 18058
rect 21650 18006 21652 18058
rect 21596 18004 21652 18006
rect 21700 18058 21756 18060
rect 21700 18006 21702 18058
rect 21702 18006 21754 18058
rect 21754 18006 21756 18058
rect 21700 18004 21756 18006
rect 21804 18058 21860 18060
rect 21804 18006 21806 18058
rect 21806 18006 21858 18058
rect 21858 18006 21860 18058
rect 21804 18004 21860 18006
rect 21980 17778 22036 17780
rect 21980 17726 21982 17778
rect 21982 17726 22034 17778
rect 22034 17726 22036 17778
rect 21980 17724 22036 17726
rect 23996 20748 24052 20804
rect 24508 20410 24564 20412
rect 24508 20358 24510 20410
rect 24510 20358 24562 20410
rect 24562 20358 24564 20410
rect 24508 20356 24564 20358
rect 24612 20410 24668 20412
rect 24612 20358 24614 20410
rect 24614 20358 24666 20410
rect 24666 20358 24668 20410
rect 24612 20356 24668 20358
rect 24716 20410 24772 20412
rect 24716 20358 24718 20410
rect 24718 20358 24770 20410
rect 24770 20358 24772 20410
rect 24716 20356 24772 20358
rect 22876 19346 22932 19348
rect 22876 19294 22878 19346
rect 22878 19294 22930 19346
rect 22930 19294 22932 19346
rect 22876 19292 22932 19294
rect 22988 19234 23044 19236
rect 22988 19182 22990 19234
rect 22990 19182 23042 19234
rect 23042 19182 23044 19234
rect 22988 19180 23044 19182
rect 22764 18620 22820 18676
rect 23548 18450 23604 18452
rect 23548 18398 23550 18450
rect 23550 18398 23602 18450
rect 23602 18398 23604 18450
rect 23548 18396 23604 18398
rect 22876 18338 22932 18340
rect 22876 18286 22878 18338
rect 22878 18286 22930 18338
rect 22930 18286 22932 18338
rect 22876 18284 22932 18286
rect 23100 17836 23156 17892
rect 21980 17388 22036 17444
rect 21596 16490 21652 16492
rect 21596 16438 21598 16490
rect 21598 16438 21650 16490
rect 21650 16438 21652 16490
rect 21596 16436 21652 16438
rect 21700 16490 21756 16492
rect 21700 16438 21702 16490
rect 21702 16438 21754 16490
rect 21754 16438 21756 16490
rect 21700 16436 21756 16438
rect 21804 16490 21860 16492
rect 21804 16438 21806 16490
rect 21806 16438 21858 16490
rect 21858 16438 21860 16490
rect 21804 16436 21860 16438
rect 21308 15260 21364 15316
rect 21532 16098 21588 16100
rect 21532 16046 21534 16098
rect 21534 16046 21586 16098
rect 21586 16046 21588 16098
rect 21532 16044 21588 16046
rect 22316 16828 22372 16884
rect 21644 15090 21700 15092
rect 21644 15038 21646 15090
rect 21646 15038 21698 15090
rect 21698 15038 21700 15090
rect 21644 15036 21700 15038
rect 21980 15260 22036 15316
rect 21868 15036 21924 15092
rect 21596 14922 21652 14924
rect 21596 14870 21598 14922
rect 21598 14870 21650 14922
rect 21650 14870 21652 14922
rect 21596 14868 21652 14870
rect 21700 14922 21756 14924
rect 21700 14870 21702 14922
rect 21702 14870 21754 14922
rect 21754 14870 21756 14922
rect 21700 14868 21756 14870
rect 21804 14922 21860 14924
rect 21804 14870 21806 14922
rect 21806 14870 21858 14922
rect 21858 14870 21860 14922
rect 21804 14868 21860 14870
rect 23884 17442 23940 17444
rect 23884 17390 23886 17442
rect 23886 17390 23938 17442
rect 23938 17390 23940 17442
rect 23884 17388 23940 17390
rect 23436 16940 23492 16996
rect 23324 16828 23380 16884
rect 22316 13916 22372 13972
rect 21420 13356 21476 13412
rect 20748 12908 20804 12964
rect 19628 12348 19684 12404
rect 20860 12348 20916 12404
rect 18684 11002 18740 11004
rect 18684 10950 18686 11002
rect 18686 10950 18738 11002
rect 18738 10950 18740 11002
rect 18684 10948 18740 10950
rect 18788 11002 18844 11004
rect 18788 10950 18790 11002
rect 18790 10950 18842 11002
rect 18842 10950 18844 11002
rect 18788 10948 18844 10950
rect 18892 11002 18948 11004
rect 18892 10950 18894 11002
rect 18894 10950 18946 11002
rect 18946 10950 18948 11002
rect 18892 10948 18948 10950
rect 19740 11788 19796 11844
rect 20300 11788 20356 11844
rect 20076 11340 20132 11396
rect 19628 10556 19684 10612
rect 19516 10332 19572 10388
rect 16268 7308 16324 7364
rect 16828 8876 16884 8932
rect 17388 8876 17444 8932
rect 15772 7082 15828 7084
rect 15772 7030 15774 7082
rect 15774 7030 15826 7082
rect 15826 7030 15828 7082
rect 15772 7028 15828 7030
rect 15876 7082 15932 7084
rect 15876 7030 15878 7082
rect 15878 7030 15930 7082
rect 15930 7030 15932 7082
rect 15876 7028 15932 7030
rect 15980 7082 16036 7084
rect 15980 7030 15982 7082
rect 15982 7030 16034 7082
rect 16034 7030 16036 7082
rect 15980 7028 16036 7030
rect 12124 6466 12180 6468
rect 12124 6414 12126 6466
rect 12126 6414 12178 6466
rect 12178 6414 12180 6466
rect 12124 6412 12180 6414
rect 13468 6412 13524 6468
rect 12860 6298 12916 6300
rect 12860 6246 12862 6298
rect 12862 6246 12914 6298
rect 12914 6246 12916 6298
rect 12860 6244 12916 6246
rect 12964 6298 13020 6300
rect 12964 6246 12966 6298
rect 12966 6246 13018 6298
rect 13018 6246 13020 6298
rect 12964 6244 13020 6246
rect 13068 6298 13124 6300
rect 13068 6246 13070 6298
rect 13070 6246 13122 6298
rect 13122 6246 13124 6298
rect 13068 6244 13124 6246
rect 14252 5906 14308 5908
rect 14252 5854 14254 5906
rect 14254 5854 14306 5906
rect 14306 5854 14308 5906
rect 14252 5852 14308 5854
rect 18684 9434 18740 9436
rect 18684 9382 18686 9434
rect 18686 9382 18738 9434
rect 18738 9382 18740 9434
rect 18684 9380 18740 9382
rect 18788 9434 18844 9436
rect 18788 9382 18790 9434
rect 18790 9382 18842 9434
rect 18842 9382 18844 9434
rect 18788 9380 18844 9382
rect 18892 9434 18948 9436
rect 18892 9382 18894 9434
rect 18894 9382 18946 9434
rect 18946 9382 18948 9434
rect 18892 9380 18948 9382
rect 20300 10332 20356 10388
rect 21308 12796 21364 12852
rect 21596 13354 21652 13356
rect 21596 13302 21598 13354
rect 21598 13302 21650 13354
rect 21650 13302 21652 13354
rect 21596 13300 21652 13302
rect 21700 13354 21756 13356
rect 21700 13302 21702 13354
rect 21702 13302 21754 13354
rect 21754 13302 21756 13354
rect 21700 13300 21756 13302
rect 21804 13354 21860 13356
rect 21804 13302 21806 13354
rect 21806 13302 21858 13354
rect 21858 13302 21860 13354
rect 21804 13300 21860 13302
rect 21532 12348 21588 12404
rect 22204 12850 22260 12852
rect 22204 12798 22206 12850
rect 22206 12798 22258 12850
rect 22258 12798 22260 12850
rect 22204 12796 22260 12798
rect 20860 11900 20916 11956
rect 20636 11228 20692 11284
rect 21980 12012 22036 12068
rect 21084 11788 21140 11844
rect 20636 10332 20692 10388
rect 20972 10444 21028 10500
rect 20188 9714 20244 9716
rect 20188 9662 20190 9714
rect 20190 9662 20242 9714
rect 20242 9662 20244 9714
rect 20188 9660 20244 9662
rect 18684 7866 18740 7868
rect 18684 7814 18686 7866
rect 18686 7814 18738 7866
rect 18738 7814 18740 7866
rect 18684 7812 18740 7814
rect 18788 7866 18844 7868
rect 18788 7814 18790 7866
rect 18790 7814 18842 7866
rect 18842 7814 18844 7866
rect 18788 7812 18844 7814
rect 18892 7866 18948 7868
rect 18892 7814 18894 7866
rect 18894 7814 18946 7866
rect 18946 7814 18948 7866
rect 18892 7812 18948 7814
rect 19852 8876 19908 8932
rect 20300 8930 20356 8932
rect 20300 8878 20302 8930
rect 20302 8878 20354 8930
rect 20354 8878 20356 8930
rect 20300 8876 20356 8878
rect 20188 8764 20244 8820
rect 20972 9996 21028 10052
rect 20636 9436 20692 9492
rect 20748 9212 20804 9268
rect 20636 8876 20692 8932
rect 21596 11786 21652 11788
rect 21596 11734 21598 11786
rect 21598 11734 21650 11786
rect 21650 11734 21652 11786
rect 21596 11732 21652 11734
rect 21700 11786 21756 11788
rect 21700 11734 21702 11786
rect 21702 11734 21754 11786
rect 21754 11734 21756 11786
rect 21700 11732 21756 11734
rect 21804 11786 21860 11788
rect 21804 11734 21806 11786
rect 21806 11734 21858 11786
rect 21858 11734 21860 11786
rect 21804 11732 21860 11734
rect 22092 11900 22148 11956
rect 21420 11394 21476 11396
rect 21420 11342 21422 11394
rect 21422 11342 21474 11394
rect 21474 11342 21476 11394
rect 21420 11340 21476 11342
rect 21980 11282 22036 11284
rect 21980 11230 21982 11282
rect 21982 11230 22034 11282
rect 22034 11230 22036 11282
rect 21980 11228 22036 11230
rect 21308 10108 21364 10164
rect 21644 10610 21700 10612
rect 21644 10558 21646 10610
rect 21646 10558 21698 10610
rect 21698 10558 21700 10610
rect 21644 10556 21700 10558
rect 21532 10498 21588 10500
rect 21532 10446 21534 10498
rect 21534 10446 21586 10498
rect 21586 10446 21588 10498
rect 21532 10444 21588 10446
rect 21596 10218 21652 10220
rect 21596 10166 21598 10218
rect 21598 10166 21650 10218
rect 21650 10166 21652 10218
rect 21596 10164 21652 10166
rect 21700 10218 21756 10220
rect 21700 10166 21702 10218
rect 21702 10166 21754 10218
rect 21754 10166 21756 10218
rect 21700 10164 21756 10166
rect 21804 10218 21860 10220
rect 21804 10166 21806 10218
rect 21806 10166 21858 10218
rect 21858 10166 21860 10218
rect 21804 10164 21860 10166
rect 23660 16882 23716 16884
rect 23660 16830 23662 16882
rect 23662 16830 23714 16882
rect 23714 16830 23716 16882
rect 23660 16828 23716 16830
rect 23884 16882 23940 16884
rect 23884 16830 23886 16882
rect 23886 16830 23938 16882
rect 23938 16830 23940 16882
rect 23884 16828 23940 16830
rect 24508 18842 24564 18844
rect 24508 18790 24510 18842
rect 24510 18790 24562 18842
rect 24562 18790 24564 18842
rect 24508 18788 24564 18790
rect 24612 18842 24668 18844
rect 24612 18790 24614 18842
rect 24614 18790 24666 18842
rect 24666 18790 24668 18842
rect 24612 18788 24668 18790
rect 24716 18842 24772 18844
rect 24716 18790 24718 18842
rect 24718 18790 24770 18842
rect 24770 18790 24772 18842
rect 24716 18788 24772 18790
rect 24108 18620 24164 18676
rect 24108 18450 24164 18452
rect 24108 18398 24110 18450
rect 24110 18398 24162 18450
rect 24162 18398 24164 18450
rect 24108 18396 24164 18398
rect 24508 17274 24564 17276
rect 24508 17222 24510 17274
rect 24510 17222 24562 17274
rect 24562 17222 24564 17274
rect 24508 17220 24564 17222
rect 24612 17274 24668 17276
rect 24612 17222 24614 17274
rect 24614 17222 24666 17274
rect 24666 17222 24668 17274
rect 24612 17220 24668 17222
rect 24716 17274 24772 17276
rect 24716 17222 24718 17274
rect 24718 17222 24770 17274
rect 24770 17222 24772 17274
rect 24716 17220 24772 17222
rect 24108 16828 24164 16884
rect 22764 12402 22820 12404
rect 22764 12350 22766 12402
rect 22766 12350 22818 12402
rect 22818 12350 22820 12402
rect 22764 12348 22820 12350
rect 23212 12962 23268 12964
rect 23212 12910 23214 12962
rect 23214 12910 23266 12962
rect 23266 12910 23268 12962
rect 23212 12908 23268 12910
rect 23884 15036 23940 15092
rect 23660 14812 23716 14868
rect 23436 14588 23492 14644
rect 23660 14252 23716 14308
rect 22988 12012 23044 12068
rect 23324 11228 23380 11284
rect 23884 13970 23940 13972
rect 23884 13918 23886 13970
rect 23886 13918 23938 13970
rect 23938 13918 23940 13970
rect 23884 13916 23940 13918
rect 24332 15932 24388 15988
rect 24508 15706 24564 15708
rect 24508 15654 24510 15706
rect 24510 15654 24562 15706
rect 24562 15654 24564 15706
rect 24508 15652 24564 15654
rect 24612 15706 24668 15708
rect 24612 15654 24614 15706
rect 24614 15654 24666 15706
rect 24666 15654 24668 15706
rect 24612 15652 24668 15654
rect 24716 15706 24772 15708
rect 24716 15654 24718 15706
rect 24718 15654 24770 15706
rect 24770 15654 24772 15706
rect 24716 15652 24772 15654
rect 24332 14700 24388 14756
rect 24508 14138 24564 14140
rect 24508 14086 24510 14138
rect 24510 14086 24562 14138
rect 24562 14086 24564 14138
rect 24508 14084 24564 14086
rect 24612 14138 24668 14140
rect 24612 14086 24614 14138
rect 24614 14086 24666 14138
rect 24666 14086 24668 14138
rect 24612 14084 24668 14086
rect 24716 14138 24772 14140
rect 24716 14086 24718 14138
rect 24718 14086 24770 14138
rect 24770 14086 24772 14138
rect 24716 14084 24772 14086
rect 24220 13692 24276 13748
rect 24220 12796 24276 12852
rect 24220 12572 24276 12628
rect 23548 11394 23604 11396
rect 23548 11342 23550 11394
rect 23550 11342 23602 11394
rect 23602 11342 23604 11394
rect 23548 11340 23604 11342
rect 22764 9884 22820 9940
rect 21868 9324 21924 9380
rect 21420 9100 21476 9156
rect 21756 9100 21812 9156
rect 21644 9042 21700 9044
rect 21644 8990 21646 9042
rect 21646 8990 21698 9042
rect 21698 8990 21700 9042
rect 21644 8988 21700 8990
rect 21196 8652 21252 8708
rect 18284 6636 18340 6692
rect 17836 6076 17892 6132
rect 18684 6298 18740 6300
rect 18684 6246 18686 6298
rect 18686 6246 18738 6298
rect 18738 6246 18740 6298
rect 18684 6244 18740 6246
rect 18788 6298 18844 6300
rect 18788 6246 18790 6298
rect 18790 6246 18842 6298
rect 18842 6246 18844 6298
rect 18788 6244 18844 6246
rect 18892 6298 18948 6300
rect 18892 6246 18894 6298
rect 18894 6246 18946 6298
rect 18946 6246 18948 6298
rect 18892 6244 18948 6246
rect 18508 6130 18564 6132
rect 18508 6078 18510 6130
rect 18510 6078 18562 6130
rect 18562 6078 18564 6130
rect 18508 6076 18564 6078
rect 18732 6076 18788 6132
rect 17052 5852 17108 5908
rect 19740 6076 19796 6132
rect 20076 7474 20132 7476
rect 20076 7422 20078 7474
rect 20078 7422 20130 7474
rect 20130 7422 20132 7474
rect 20076 7420 20132 7422
rect 20636 6636 20692 6692
rect 19964 5852 20020 5908
rect 20412 5906 20468 5908
rect 20412 5854 20414 5906
rect 20414 5854 20466 5906
rect 20466 5854 20468 5906
rect 20412 5852 20468 5854
rect 21596 8650 21652 8652
rect 21596 8598 21598 8650
rect 21598 8598 21650 8650
rect 21650 8598 21652 8650
rect 21596 8596 21652 8598
rect 21700 8650 21756 8652
rect 21700 8598 21702 8650
rect 21702 8598 21754 8650
rect 21754 8598 21756 8650
rect 21700 8596 21756 8598
rect 21804 8650 21860 8652
rect 21804 8598 21806 8650
rect 21806 8598 21858 8650
rect 21858 8598 21860 8650
rect 21804 8596 21860 8598
rect 21644 8482 21700 8484
rect 21644 8430 21646 8482
rect 21646 8430 21698 8482
rect 21698 8430 21700 8482
rect 21644 8428 21700 8430
rect 22764 9266 22820 9268
rect 22764 9214 22766 9266
rect 22766 9214 22818 9266
rect 22818 9214 22820 9266
rect 22764 9212 22820 9214
rect 21532 7698 21588 7700
rect 21532 7646 21534 7698
rect 21534 7646 21586 7698
rect 21586 7646 21588 7698
rect 21532 7644 21588 7646
rect 21980 8258 22036 8260
rect 21980 8206 21982 8258
rect 21982 8206 22034 8258
rect 22034 8206 22036 8258
rect 21980 8204 22036 8206
rect 21596 7082 21652 7084
rect 21596 7030 21598 7082
rect 21598 7030 21650 7082
rect 21650 7030 21652 7082
rect 21596 7028 21652 7030
rect 21700 7082 21756 7084
rect 21700 7030 21702 7082
rect 21702 7030 21754 7082
rect 21754 7030 21756 7082
rect 21700 7028 21756 7030
rect 21804 7082 21860 7084
rect 21804 7030 21806 7082
rect 21806 7030 21858 7082
rect 21858 7030 21860 7082
rect 21804 7028 21860 7030
rect 20748 6524 20804 6580
rect 22764 8428 22820 8484
rect 23548 9996 23604 10052
rect 23548 9324 23604 9380
rect 23436 8428 23492 8484
rect 23884 9042 23940 9044
rect 23884 8990 23886 9042
rect 23886 8990 23938 9042
rect 23938 8990 23940 9042
rect 23884 8988 23940 8990
rect 22652 7698 22708 7700
rect 22652 7646 22654 7698
rect 22654 7646 22706 7698
rect 22706 7646 22708 7698
rect 22652 7644 22708 7646
rect 22204 7420 22260 7476
rect 23324 7474 23380 7476
rect 23324 7422 23326 7474
rect 23326 7422 23378 7474
rect 23378 7422 23380 7474
rect 23324 7420 23380 7422
rect 23212 6748 23268 6804
rect 22092 6578 22148 6580
rect 22092 6526 22094 6578
rect 22094 6526 22146 6578
rect 22146 6526 22148 6578
rect 22092 6524 22148 6526
rect 21980 5852 22036 5908
rect 22428 5852 22484 5908
rect 9948 5514 10004 5516
rect 9948 5462 9950 5514
rect 9950 5462 10002 5514
rect 10002 5462 10004 5514
rect 9948 5460 10004 5462
rect 10052 5514 10108 5516
rect 10052 5462 10054 5514
rect 10054 5462 10106 5514
rect 10106 5462 10108 5514
rect 10052 5460 10108 5462
rect 10156 5514 10212 5516
rect 10156 5462 10158 5514
rect 10158 5462 10210 5514
rect 10210 5462 10212 5514
rect 10156 5460 10212 5462
rect 15772 5514 15828 5516
rect 15772 5462 15774 5514
rect 15774 5462 15826 5514
rect 15826 5462 15828 5514
rect 15772 5460 15828 5462
rect 15876 5514 15932 5516
rect 15876 5462 15878 5514
rect 15878 5462 15930 5514
rect 15930 5462 15932 5514
rect 15876 5460 15932 5462
rect 15980 5514 16036 5516
rect 15980 5462 15982 5514
rect 15982 5462 16034 5514
rect 16034 5462 16036 5514
rect 15980 5460 16036 5462
rect 21596 5514 21652 5516
rect 21596 5462 21598 5514
rect 21598 5462 21650 5514
rect 21650 5462 21652 5514
rect 21596 5460 21652 5462
rect 21700 5514 21756 5516
rect 21700 5462 21702 5514
rect 21702 5462 21754 5514
rect 21754 5462 21756 5514
rect 21700 5460 21756 5462
rect 21804 5514 21860 5516
rect 21804 5462 21806 5514
rect 21806 5462 21858 5514
rect 21858 5462 21860 5514
rect 21804 5460 21860 5462
rect 7036 4730 7092 4732
rect 7036 4678 7038 4730
rect 7038 4678 7090 4730
rect 7090 4678 7092 4730
rect 7036 4676 7092 4678
rect 7140 4730 7196 4732
rect 7140 4678 7142 4730
rect 7142 4678 7194 4730
rect 7194 4678 7196 4730
rect 7140 4676 7196 4678
rect 7244 4730 7300 4732
rect 7244 4678 7246 4730
rect 7246 4678 7298 4730
rect 7298 4678 7300 4730
rect 7244 4676 7300 4678
rect 12860 4730 12916 4732
rect 12860 4678 12862 4730
rect 12862 4678 12914 4730
rect 12914 4678 12916 4730
rect 12860 4676 12916 4678
rect 12964 4730 13020 4732
rect 12964 4678 12966 4730
rect 12966 4678 13018 4730
rect 13018 4678 13020 4730
rect 12964 4676 13020 4678
rect 13068 4730 13124 4732
rect 13068 4678 13070 4730
rect 13070 4678 13122 4730
rect 13122 4678 13124 4730
rect 13068 4676 13124 4678
rect 18684 4730 18740 4732
rect 18684 4678 18686 4730
rect 18686 4678 18738 4730
rect 18738 4678 18740 4730
rect 18684 4676 18740 4678
rect 18788 4730 18844 4732
rect 18788 4678 18790 4730
rect 18790 4678 18842 4730
rect 18842 4678 18844 4730
rect 18788 4676 18844 4678
rect 18892 4730 18948 4732
rect 18892 4678 18894 4730
rect 18894 4678 18946 4730
rect 18946 4678 18948 4730
rect 18892 4676 18948 4678
rect 4124 3946 4180 3948
rect 4124 3894 4126 3946
rect 4126 3894 4178 3946
rect 4178 3894 4180 3946
rect 4124 3892 4180 3894
rect 4228 3946 4284 3948
rect 4228 3894 4230 3946
rect 4230 3894 4282 3946
rect 4282 3894 4284 3946
rect 4228 3892 4284 3894
rect 4332 3946 4388 3948
rect 4332 3894 4334 3946
rect 4334 3894 4386 3946
rect 4386 3894 4388 3946
rect 4332 3892 4388 3894
rect 9948 3946 10004 3948
rect 9948 3894 9950 3946
rect 9950 3894 10002 3946
rect 10002 3894 10004 3946
rect 9948 3892 10004 3894
rect 10052 3946 10108 3948
rect 10052 3894 10054 3946
rect 10054 3894 10106 3946
rect 10106 3894 10108 3946
rect 10052 3892 10108 3894
rect 10156 3946 10212 3948
rect 10156 3894 10158 3946
rect 10158 3894 10210 3946
rect 10210 3894 10212 3946
rect 10156 3892 10212 3894
rect 15772 3946 15828 3948
rect 15772 3894 15774 3946
rect 15774 3894 15826 3946
rect 15826 3894 15828 3946
rect 15772 3892 15828 3894
rect 15876 3946 15932 3948
rect 15876 3894 15878 3946
rect 15878 3894 15930 3946
rect 15930 3894 15932 3946
rect 15876 3892 15932 3894
rect 15980 3946 16036 3948
rect 15980 3894 15982 3946
rect 15982 3894 16034 3946
rect 16034 3894 16036 3946
rect 15980 3892 16036 3894
rect 21596 3946 21652 3948
rect 21596 3894 21598 3946
rect 21598 3894 21650 3946
rect 21650 3894 21652 3946
rect 21596 3892 21652 3894
rect 21700 3946 21756 3948
rect 21700 3894 21702 3946
rect 21702 3894 21754 3946
rect 21754 3894 21756 3946
rect 21700 3892 21756 3894
rect 21804 3946 21860 3948
rect 21804 3894 21806 3946
rect 21806 3894 21858 3946
rect 21858 3894 21860 3946
rect 21804 3892 21860 3894
rect 23436 3442 23492 3444
rect 23436 3390 23438 3442
rect 23438 3390 23490 3442
rect 23490 3390 23492 3442
rect 23436 3388 23492 3390
rect 23660 5234 23716 5236
rect 23660 5182 23662 5234
rect 23662 5182 23714 5234
rect 23714 5182 23716 5234
rect 23660 5180 23716 5182
rect 24508 12570 24564 12572
rect 24508 12518 24510 12570
rect 24510 12518 24562 12570
rect 24562 12518 24564 12570
rect 24508 12516 24564 12518
rect 24612 12570 24668 12572
rect 24612 12518 24614 12570
rect 24614 12518 24666 12570
rect 24666 12518 24668 12570
rect 24612 12516 24668 12518
rect 24716 12570 24772 12572
rect 24716 12518 24718 12570
rect 24718 12518 24770 12570
rect 24770 12518 24772 12570
rect 24716 12516 24772 12518
rect 24332 11900 24388 11956
rect 24892 11340 24948 11396
rect 24508 11002 24564 11004
rect 24508 10950 24510 11002
rect 24510 10950 24562 11002
rect 24562 10950 24564 11002
rect 24508 10948 24564 10950
rect 24612 11002 24668 11004
rect 24612 10950 24614 11002
rect 24614 10950 24666 11002
rect 24666 10950 24668 11002
rect 24612 10948 24668 10950
rect 24716 11002 24772 11004
rect 24716 10950 24718 11002
rect 24718 10950 24770 11002
rect 24770 10950 24772 11002
rect 24716 10948 24772 10950
rect 24508 9434 24564 9436
rect 24508 9382 24510 9434
rect 24510 9382 24562 9434
rect 24562 9382 24564 9434
rect 24508 9380 24564 9382
rect 24612 9434 24668 9436
rect 24612 9382 24614 9434
rect 24614 9382 24666 9434
rect 24666 9382 24668 9434
rect 24612 9380 24668 9382
rect 24716 9434 24772 9436
rect 24716 9382 24718 9434
rect 24718 9382 24770 9434
rect 24770 9382 24772 9434
rect 24716 9380 24772 9382
rect 24220 8988 24276 9044
rect 24508 7866 24564 7868
rect 24508 7814 24510 7866
rect 24510 7814 24562 7866
rect 24562 7814 24564 7866
rect 24508 7812 24564 7814
rect 24612 7866 24668 7868
rect 24612 7814 24614 7866
rect 24614 7814 24666 7866
rect 24666 7814 24668 7866
rect 24612 7812 24668 7814
rect 24716 7866 24772 7868
rect 24716 7814 24718 7866
rect 24718 7814 24770 7866
rect 24770 7814 24772 7866
rect 24716 7812 24772 7814
rect 24220 6802 24276 6804
rect 24220 6750 24222 6802
rect 24222 6750 24274 6802
rect 24274 6750 24276 6802
rect 24220 6748 24276 6750
rect 24508 6298 24564 6300
rect 24508 6246 24510 6298
rect 24510 6246 24562 6298
rect 24562 6246 24564 6298
rect 24508 6244 24564 6246
rect 24612 6298 24668 6300
rect 24612 6246 24614 6298
rect 24614 6246 24666 6298
rect 24666 6246 24668 6298
rect 24612 6244 24668 6246
rect 24716 6298 24772 6300
rect 24716 6246 24718 6298
rect 24718 6246 24770 6298
rect 24770 6246 24772 6298
rect 24716 6244 24772 6246
rect 24220 5852 24276 5908
rect 24220 5180 24276 5236
rect 24508 4730 24564 4732
rect 24508 4678 24510 4730
rect 24510 4678 24562 4730
rect 24562 4678 24564 4730
rect 24508 4676 24564 4678
rect 24612 4730 24668 4732
rect 24612 4678 24614 4730
rect 24614 4678 24666 4730
rect 24666 4678 24668 4730
rect 24612 4676 24668 4678
rect 24716 4730 24772 4732
rect 24716 4678 24718 4730
rect 24718 4678 24770 4730
rect 24770 4678 24772 4730
rect 24716 4676 24772 4678
rect 24220 3836 24276 3892
rect 23884 3388 23940 3444
rect 7036 3162 7092 3164
rect 7036 3110 7038 3162
rect 7038 3110 7090 3162
rect 7090 3110 7092 3162
rect 7036 3108 7092 3110
rect 7140 3162 7196 3164
rect 7140 3110 7142 3162
rect 7142 3110 7194 3162
rect 7194 3110 7196 3162
rect 7140 3108 7196 3110
rect 7244 3162 7300 3164
rect 7244 3110 7246 3162
rect 7246 3110 7298 3162
rect 7298 3110 7300 3162
rect 7244 3108 7300 3110
rect 12860 3162 12916 3164
rect 12860 3110 12862 3162
rect 12862 3110 12914 3162
rect 12914 3110 12916 3162
rect 12860 3108 12916 3110
rect 12964 3162 13020 3164
rect 12964 3110 12966 3162
rect 12966 3110 13018 3162
rect 13018 3110 13020 3162
rect 12964 3108 13020 3110
rect 13068 3162 13124 3164
rect 13068 3110 13070 3162
rect 13070 3110 13122 3162
rect 13122 3110 13124 3162
rect 13068 3108 13124 3110
rect 18684 3162 18740 3164
rect 18684 3110 18686 3162
rect 18686 3110 18738 3162
rect 18738 3110 18740 3162
rect 18684 3108 18740 3110
rect 18788 3162 18844 3164
rect 18788 3110 18790 3162
rect 18790 3110 18842 3162
rect 18842 3110 18844 3162
rect 18788 3108 18844 3110
rect 18892 3162 18948 3164
rect 18892 3110 18894 3162
rect 18894 3110 18946 3162
rect 18946 3110 18948 3162
rect 18892 3108 18948 3110
rect 24508 3162 24564 3164
rect 24508 3110 24510 3162
rect 24510 3110 24562 3162
rect 24562 3110 24564 3162
rect 24508 3108 24564 3110
rect 24612 3162 24668 3164
rect 24612 3110 24614 3162
rect 24614 3110 24666 3162
rect 24666 3110 24668 3162
rect 24612 3108 24668 3110
rect 24716 3162 24772 3164
rect 24716 3110 24718 3162
rect 24718 3110 24770 3162
rect 24770 3110 24772 3162
rect 24716 3108 24772 3110
rect 23996 1820 24052 1876
<< metal3 >>
rect 25200 24052 26000 24080
rect 20290 23996 20300 24052
rect 20356 23996 26000 24052
rect 25200 23968 26000 23996
rect 4114 22708 4124 22764
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4388 22708 4398 22764
rect 9938 22708 9948 22764
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 10212 22708 10222 22764
rect 15762 22708 15772 22764
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 16036 22708 16046 22764
rect 21586 22708 21596 22764
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21860 22708 21870 22764
rect 21298 22540 21308 22596
rect 21364 22540 22428 22596
rect 22484 22540 22494 22596
rect 19170 22092 19180 22148
rect 19236 22092 20860 22148
rect 20916 22092 24948 22148
rect 24892 22036 24948 22092
rect 25200 22036 26000 22064
rect 24892 21980 26000 22036
rect 7026 21924 7036 21980
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7300 21924 7310 21980
rect 12850 21924 12860 21980
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 13124 21924 13134 21980
rect 18674 21924 18684 21980
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18948 21924 18958 21980
rect 24498 21924 24508 21980
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24772 21924 24782 21980
rect 25200 21952 26000 21980
rect 21074 21868 21084 21924
rect 21140 21868 23660 21924
rect 23716 21868 23726 21924
rect 7634 21756 7644 21812
rect 7700 21756 8204 21812
rect 8260 21756 8270 21812
rect 17490 21644 17500 21700
rect 17556 21644 18508 21700
rect 18564 21644 21420 21700
rect 21476 21644 21486 21700
rect 13010 21532 13020 21588
rect 13076 21532 15708 21588
rect 15764 21532 16268 21588
rect 16324 21532 17948 21588
rect 18004 21532 18396 21588
rect 18452 21532 18462 21588
rect 20178 21532 20188 21588
rect 20244 21532 23548 21588
rect 23604 21532 23614 21588
rect 18722 21420 18732 21476
rect 18788 21420 20412 21476
rect 20468 21420 20478 21476
rect 2258 21308 2268 21364
rect 2324 21308 5068 21364
rect 5124 21308 9660 21364
rect 9716 21308 9726 21364
rect 16482 21308 16492 21364
rect 16548 21308 17500 21364
rect 17556 21308 17566 21364
rect 4114 21140 4124 21196
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4388 21140 4398 21196
rect 9938 21140 9948 21196
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 10212 21140 10222 21196
rect 15762 21140 15772 21196
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 16036 21140 16046 21196
rect 21586 21140 21596 21196
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21860 21140 21870 21196
rect 7858 20748 7868 20804
rect 7924 20748 8652 20804
rect 8708 20748 8718 20804
rect 19506 20748 19516 20804
rect 19572 20748 20860 20804
rect 20916 20748 20926 20804
rect 22418 20748 22428 20804
rect 22484 20748 23212 20804
rect 23268 20748 23996 20804
rect 24052 20748 24062 20804
rect 20626 20636 20636 20692
rect 20692 20636 21756 20692
rect 21812 20636 21822 20692
rect 7746 20524 7756 20580
rect 7812 20524 9996 20580
rect 10052 20524 10062 20580
rect 20402 20524 20412 20580
rect 20468 20524 21868 20580
rect 21924 20524 21934 20580
rect 8418 20412 8428 20468
rect 8484 20412 10444 20468
rect 10500 20412 10510 20468
rect 7026 20356 7036 20412
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7300 20356 7310 20412
rect 12850 20356 12860 20412
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 13124 20356 13134 20412
rect 18674 20356 18684 20412
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18948 20356 18958 20412
rect 24498 20356 24508 20412
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24772 20356 24782 20412
rect 7634 20300 7644 20356
rect 7700 20300 8316 20356
rect 8372 20300 10556 20356
rect 10612 20300 10622 20356
rect 6738 20188 6748 20244
rect 6804 20188 8092 20244
rect 8148 20188 9884 20244
rect 9940 20188 9950 20244
rect 20850 20188 20860 20244
rect 20916 20188 21868 20244
rect 21924 20188 23212 20244
rect 23268 20188 23278 20244
rect 13234 20076 13244 20132
rect 13300 20076 14140 20132
rect 14196 20076 14924 20132
rect 14980 20076 15148 20132
rect 15204 20076 15214 20132
rect 16566 20076 16604 20132
rect 16660 20076 16670 20132
rect 17266 20076 17276 20132
rect 17332 20076 17948 20132
rect 18004 20076 18732 20132
rect 18788 20076 19404 20132
rect 19460 20076 20524 20132
rect 20580 20076 21196 20132
rect 21252 20076 21262 20132
rect 25200 20020 26000 20048
rect 7970 19964 7980 20020
rect 8036 19964 9548 20020
rect 9604 19964 10780 20020
rect 10836 19964 10846 20020
rect 21074 19964 21084 20020
rect 21140 19964 21532 20020
rect 21588 19964 26000 20020
rect 25200 19936 26000 19964
rect 5394 19852 5404 19908
rect 5460 19852 6636 19908
rect 6692 19852 8316 19908
rect 8372 19852 8382 19908
rect 9874 19852 9884 19908
rect 9940 19852 11228 19908
rect 11284 19852 11294 19908
rect 12898 19740 12908 19796
rect 12964 19740 13804 19796
rect 13860 19740 13870 19796
rect 15092 19740 16044 19796
rect 16100 19740 16110 19796
rect 16706 19740 16716 19796
rect 16772 19740 17836 19796
rect 17892 19740 17902 19796
rect 19954 19740 19964 19796
rect 20020 19740 21644 19796
rect 21700 19740 22036 19796
rect 15092 19684 15148 19740
rect 11778 19628 11788 19684
rect 11844 19628 15148 19684
rect 16482 19628 16492 19684
rect 16548 19628 16828 19684
rect 16884 19628 16894 19684
rect 4114 19572 4124 19628
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4388 19572 4398 19628
rect 9938 19572 9948 19628
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 10212 19572 10222 19628
rect 15762 19572 15772 19628
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 16036 19572 16046 19628
rect 21586 19572 21596 19628
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21860 19572 21870 19628
rect 21980 19460 22036 19740
rect 10658 19404 10668 19460
rect 10724 19404 11900 19460
rect 11956 19404 11966 19460
rect 18162 19404 18172 19460
rect 18228 19404 21420 19460
rect 21476 19404 21486 19460
rect 21634 19404 21644 19460
rect 21700 19404 22036 19460
rect 19842 19292 19852 19348
rect 19908 19292 20076 19348
rect 20132 19292 21532 19348
rect 21588 19292 22092 19348
rect 22148 19292 22876 19348
rect 22932 19292 22942 19348
rect 13906 19180 13916 19236
rect 13972 19180 14364 19236
rect 14420 19180 14430 19236
rect 14578 19180 14588 19236
rect 14644 19180 15372 19236
rect 15428 19180 15438 19236
rect 16930 19180 16940 19236
rect 16996 19180 19628 19236
rect 19684 19180 19694 19236
rect 21298 19180 21308 19236
rect 21364 19180 22988 19236
rect 23044 19180 23054 19236
rect 8642 19068 8652 19124
rect 8708 19068 9436 19124
rect 9492 19068 9772 19124
rect 9828 19068 9838 19124
rect 10098 19068 10108 19124
rect 10164 19068 10892 19124
rect 10948 19068 11452 19124
rect 11508 19068 11900 19124
rect 11956 19068 11966 19124
rect 9314 18956 9324 19012
rect 9380 18956 10332 19012
rect 10388 18956 10398 19012
rect 12338 18956 12348 19012
rect 12404 18956 14476 19012
rect 14532 18956 14542 19012
rect 14802 18956 14812 19012
rect 14868 18956 15260 19012
rect 15316 18956 16604 19012
rect 16660 18956 16670 19012
rect 20066 18956 20076 19012
rect 20132 18956 22092 19012
rect 22148 18956 22158 19012
rect 7026 18788 7036 18844
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7300 18788 7310 18844
rect 12850 18788 12860 18844
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 13124 18788 13134 18844
rect 18674 18788 18684 18844
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18948 18788 18958 18844
rect 24498 18788 24508 18844
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24772 18788 24782 18844
rect 5170 18620 5180 18676
rect 5236 18620 6748 18676
rect 6804 18620 6814 18676
rect 11106 18620 11116 18676
rect 11172 18620 12012 18676
rect 12068 18620 12078 18676
rect 14354 18620 14364 18676
rect 14420 18620 15148 18676
rect 15204 18620 15214 18676
rect 22754 18620 22764 18676
rect 22820 18620 24108 18676
rect 24164 18620 25284 18676
rect 1922 18508 1932 18564
rect 1988 18508 2940 18564
rect 2996 18508 3006 18564
rect 4610 18508 4620 18564
rect 4676 18508 7756 18564
rect 7812 18508 7822 18564
rect 3602 18396 3612 18452
rect 3668 18396 4396 18452
rect 4452 18396 4956 18452
rect 5012 18396 5628 18452
rect 5684 18396 5694 18452
rect 7298 18396 7308 18452
rect 7364 18396 8988 18452
rect 9044 18396 9772 18452
rect 9828 18396 9838 18452
rect 12226 18396 12236 18452
rect 12292 18396 12908 18452
rect 12964 18396 12974 18452
rect 14130 18396 14140 18452
rect 14196 18396 15148 18452
rect 15204 18396 15214 18452
rect 15474 18396 15484 18452
rect 15540 18396 16268 18452
rect 16324 18396 17388 18452
rect 17444 18396 17454 18452
rect 20626 18396 20636 18452
rect 20692 18396 23548 18452
rect 23604 18396 24108 18452
rect 24164 18396 24174 18452
rect 3826 18284 3836 18340
rect 3892 18284 4284 18340
rect 4340 18284 5572 18340
rect 6402 18284 6412 18340
rect 6468 18284 12572 18340
rect 12628 18284 14812 18340
rect 14868 18284 15148 18340
rect 15250 18284 15260 18340
rect 15316 18284 16156 18340
rect 16212 18284 16828 18340
rect 16884 18284 16894 18340
rect 20402 18284 20412 18340
rect 20468 18284 22876 18340
rect 22932 18284 22942 18340
rect 5516 18228 5572 18284
rect 15092 18228 15148 18284
rect 25228 18228 25284 18620
rect 3154 18172 3164 18228
rect 3220 18172 4844 18228
rect 4900 18172 4910 18228
rect 5506 18172 5516 18228
rect 5572 18172 8540 18228
rect 8596 18172 9884 18228
rect 9940 18172 9950 18228
rect 15092 18172 16380 18228
rect 16436 18172 17612 18228
rect 17668 18172 17678 18228
rect 20514 18172 20524 18228
rect 20580 18172 21532 18228
rect 21588 18172 21868 18228
rect 21924 18172 21934 18228
rect 25004 18172 25284 18228
rect 4114 18004 4124 18060
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4388 18004 4398 18060
rect 9938 18004 9948 18060
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 10212 18004 10222 18060
rect 15762 18004 15772 18060
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 16036 18004 16046 18060
rect 21586 18004 21596 18060
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21860 18004 21870 18060
rect 25004 18004 25060 18172
rect 25200 18004 26000 18032
rect 25004 17948 26000 18004
rect 25200 17920 26000 17948
rect 2482 17836 2492 17892
rect 2548 17836 4284 17892
rect 4340 17836 4350 17892
rect 9314 17836 9324 17892
rect 9380 17836 10780 17892
rect 10836 17836 11340 17892
rect 11396 17836 23100 17892
rect 23156 17836 23166 17892
rect 20738 17724 20748 17780
rect 20804 17724 21980 17780
rect 22036 17724 22046 17780
rect 17154 17612 17164 17668
rect 17220 17612 18060 17668
rect 18116 17612 19180 17668
rect 19236 17612 20300 17668
rect 20356 17612 20366 17668
rect 3938 17500 3948 17556
rect 4004 17500 12908 17556
rect 12964 17500 16940 17556
rect 16996 17500 17006 17556
rect 19506 17388 19516 17444
rect 19572 17388 20748 17444
rect 20804 17388 20814 17444
rect 21970 17388 21980 17444
rect 22036 17388 23884 17444
rect 23940 17388 23950 17444
rect 13906 17276 13916 17332
rect 13972 17276 16268 17332
rect 16324 17276 16334 17332
rect 7026 17220 7036 17276
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7300 17220 7310 17276
rect 12850 17220 12860 17276
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 13124 17220 13134 17276
rect 18674 17220 18684 17276
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18948 17220 18958 17276
rect 24498 17220 24508 17276
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24772 17220 24782 17276
rect 4386 17052 4396 17108
rect 4452 17052 4956 17108
rect 5012 17052 11004 17108
rect 11060 17052 11070 17108
rect 3154 16940 3164 16996
rect 3220 16940 3724 16996
rect 3780 16940 3790 16996
rect 7858 16940 7868 16996
rect 7924 16940 8428 16996
rect 8484 16940 9660 16996
rect 9716 16940 9726 16996
rect 16146 16940 16156 16996
rect 16212 16940 16492 16996
rect 16548 16940 23436 16996
rect 23492 16940 23502 16996
rect 5730 16828 5740 16884
rect 5796 16828 6748 16884
rect 6804 16828 6814 16884
rect 22306 16828 22316 16884
rect 22372 16828 23324 16884
rect 23380 16828 23660 16884
rect 23716 16828 23726 16884
rect 23874 16828 23884 16884
rect 23940 16828 24108 16884
rect 24164 16828 24174 16884
rect 9538 16716 9548 16772
rect 9604 16716 11004 16772
rect 11060 16716 11070 16772
rect 11778 16716 11788 16772
rect 11844 16716 13580 16772
rect 13636 16716 13646 16772
rect 5730 16604 5740 16660
rect 5796 16604 6300 16660
rect 6356 16604 6366 16660
rect 10434 16604 10444 16660
rect 10500 16604 11900 16660
rect 11956 16604 11966 16660
rect 13458 16604 13468 16660
rect 13524 16604 15484 16660
rect 15540 16604 15550 16660
rect 19282 16492 19292 16548
rect 19348 16492 20188 16548
rect 20244 16492 21308 16548
rect 21364 16492 21374 16548
rect 4114 16436 4124 16492
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4388 16436 4398 16492
rect 9938 16436 9948 16492
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 10212 16436 10222 16492
rect 15762 16436 15772 16492
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 16036 16436 16046 16492
rect 21586 16436 21596 16492
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21860 16436 21870 16492
rect 2034 16268 2044 16324
rect 2100 16268 2492 16324
rect 2548 16268 3388 16324
rect 3444 16268 3454 16324
rect 5170 16268 5180 16324
rect 5236 16268 6076 16324
rect 6132 16268 6142 16324
rect 14466 16268 14476 16324
rect 14532 16268 14812 16324
rect 14868 16268 14878 16324
rect 17266 16156 17276 16212
rect 17332 16156 20636 16212
rect 20692 16156 20702 16212
rect 2370 16044 2380 16100
rect 2436 16044 5852 16100
rect 5908 16044 5918 16100
rect 6514 16044 6524 16100
rect 6580 16044 7644 16100
rect 7700 16044 7710 16100
rect 8754 16044 8764 16100
rect 8820 16044 14924 16100
rect 14980 16044 14990 16100
rect 19618 16044 19628 16100
rect 19684 16044 21532 16100
rect 21588 16044 21598 16100
rect 25200 15988 26000 16016
rect 14690 15932 14700 15988
rect 14756 15932 15036 15988
rect 15092 15932 15596 15988
rect 15652 15932 15662 15988
rect 18050 15932 18060 15988
rect 18116 15932 20076 15988
rect 20132 15932 20142 15988
rect 24322 15932 24332 15988
rect 24388 15932 26000 15988
rect 25200 15904 26000 15932
rect 2482 15820 2492 15876
rect 2548 15820 3612 15876
rect 3668 15820 4732 15876
rect 4788 15820 4798 15876
rect 5506 15820 5516 15876
rect 5572 15820 7308 15876
rect 7364 15820 7374 15876
rect 7026 15652 7036 15708
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7300 15652 7310 15708
rect 12850 15652 12860 15708
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 13124 15652 13134 15708
rect 18674 15652 18684 15708
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18948 15652 18958 15708
rect 24498 15652 24508 15708
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24772 15652 24782 15708
rect 14914 15596 14924 15652
rect 14980 15596 17388 15652
rect 17444 15596 17454 15652
rect 15138 15484 15148 15540
rect 15204 15484 16660 15540
rect 16604 15428 16660 15484
rect 2706 15372 2716 15428
rect 2772 15372 4620 15428
rect 4676 15372 5404 15428
rect 5460 15372 5470 15428
rect 14466 15372 14476 15428
rect 14532 15372 15484 15428
rect 15540 15372 15550 15428
rect 16594 15372 16604 15428
rect 16660 15372 17388 15428
rect 17444 15372 17454 15428
rect 2034 15260 2044 15316
rect 2100 15260 2380 15316
rect 2436 15260 2446 15316
rect 3154 15260 3164 15316
rect 3220 15260 4060 15316
rect 4116 15260 4396 15316
rect 4452 15260 6636 15316
rect 6692 15260 6702 15316
rect 15586 15260 15596 15316
rect 15652 15260 16492 15316
rect 16548 15260 17612 15316
rect 17668 15260 17780 15316
rect 19394 15260 19404 15316
rect 19460 15260 20524 15316
rect 20580 15260 20590 15316
rect 21298 15260 21308 15316
rect 21364 15260 21980 15316
rect 22036 15260 22046 15316
rect 11890 15148 11900 15204
rect 11956 15148 14364 15204
rect 14420 15148 15260 15204
rect 15316 15148 15326 15204
rect 17724 15092 17780 15260
rect 1810 15036 1820 15092
rect 1876 15036 3052 15092
rect 3108 15036 5628 15092
rect 5684 15036 5694 15092
rect 7746 15036 7756 15092
rect 7812 15036 9660 15092
rect 9716 15036 9726 15092
rect 12338 15036 12348 15092
rect 12404 15036 15708 15092
rect 15764 15036 16380 15092
rect 16436 15036 16446 15092
rect 16706 15036 16716 15092
rect 16772 15036 16782 15092
rect 17724 15036 21644 15092
rect 21700 15036 21710 15092
rect 21858 15036 21868 15092
rect 21924 15036 23884 15092
rect 23940 15036 23950 15092
rect 16716 14980 16772 15036
rect 2594 14924 2604 14980
rect 2660 14924 3164 14980
rect 3220 14924 3230 14980
rect 16482 14924 16492 14980
rect 16548 14924 16772 14980
rect 4114 14868 4124 14924
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4388 14868 4398 14924
rect 9938 14868 9948 14924
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 10212 14868 10222 14924
rect 15762 14868 15772 14924
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 16036 14868 16046 14924
rect 21586 14868 21596 14924
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21860 14868 21870 14924
rect 23650 14812 23660 14868
rect 23716 14812 24220 14868
rect 24276 14812 24286 14868
rect 23492 14700 24332 14756
rect 24388 14700 24398 14756
rect 12898 14588 12908 14644
rect 12964 14588 16492 14644
rect 16548 14588 16558 14644
rect 23426 14588 23436 14644
rect 23492 14588 23548 14700
rect 1922 14476 1932 14532
rect 1988 14476 2940 14532
rect 2996 14476 3006 14532
rect 6402 14476 6412 14532
rect 6468 14476 7084 14532
rect 7140 14476 8428 14532
rect 8484 14476 8494 14532
rect 4386 14252 4396 14308
rect 4452 14252 8652 14308
rect 8708 14252 8718 14308
rect 23650 14252 23660 14308
rect 23716 14252 23884 14308
rect 23940 14252 23950 14308
rect 7026 14084 7036 14140
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7300 14084 7310 14140
rect 12850 14084 12860 14140
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 13124 14084 13134 14140
rect 18674 14084 18684 14140
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18948 14084 18958 14140
rect 24498 14084 24508 14140
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24772 14084 24782 14140
rect 25200 13972 26000 14000
rect 4946 13916 4956 13972
rect 5012 13916 8428 13972
rect 16594 13916 16604 13972
rect 16660 13916 17388 13972
rect 17444 13916 17454 13972
rect 22306 13916 22316 13972
rect 22372 13916 23884 13972
rect 23940 13916 23950 13972
rect 24444 13916 26000 13972
rect 6178 13804 6188 13860
rect 6244 13804 6860 13860
rect 6916 13804 6926 13860
rect 8372 13748 8428 13916
rect 6402 13692 6412 13748
rect 6468 13692 7084 13748
rect 7140 13692 7150 13748
rect 8372 13692 11228 13748
rect 11284 13692 11294 13748
rect 12450 13692 12460 13748
rect 12516 13692 14140 13748
rect 14196 13692 14206 13748
rect 19954 13692 19964 13748
rect 20020 13692 20300 13748
rect 20356 13692 24220 13748
rect 24276 13692 24286 13748
rect 2706 13580 2716 13636
rect 2772 13580 6972 13636
rect 7028 13580 7980 13636
rect 8036 13580 8046 13636
rect 8306 13580 8316 13636
rect 8372 13580 9548 13636
rect 9604 13580 9614 13636
rect 24444 13524 24500 13916
rect 25200 13888 26000 13916
rect 5282 13468 5292 13524
rect 5348 13468 6076 13524
rect 6132 13468 6142 13524
rect 20514 13468 20524 13524
rect 20580 13468 24500 13524
rect 20402 13356 20412 13412
rect 20468 13356 21420 13412
rect 21476 13356 21486 13412
rect 4114 13300 4124 13356
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4388 13300 4398 13356
rect 9938 13300 9948 13356
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 10212 13300 10222 13356
rect 15762 13300 15772 13356
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 16036 13300 16046 13356
rect 21586 13300 21596 13356
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21860 13300 21870 13356
rect 16706 13020 16716 13076
rect 16772 13020 18284 13076
rect 18340 13020 18350 13076
rect 5954 12908 5964 12964
rect 6020 12908 7868 12964
rect 7924 12908 7934 12964
rect 20738 12908 20748 12964
rect 20804 12908 23212 12964
rect 23268 12908 23278 12964
rect 18386 12796 18396 12852
rect 18452 12796 21308 12852
rect 21364 12796 21374 12852
rect 22194 12796 22204 12852
rect 22260 12796 24220 12852
rect 24276 12796 24286 12852
rect 24182 12572 24220 12628
rect 24276 12572 24286 12628
rect 7026 12516 7036 12572
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7300 12516 7310 12572
rect 12850 12516 12860 12572
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 13124 12516 13134 12572
rect 18674 12516 18684 12572
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18948 12516 18958 12572
rect 24498 12516 24508 12572
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24772 12516 24782 12572
rect 14242 12348 14252 12404
rect 14308 12348 15484 12404
rect 15540 12348 17500 12404
rect 17556 12348 17566 12404
rect 19282 12348 19292 12404
rect 19348 12348 19628 12404
rect 19684 12348 20860 12404
rect 20916 12348 20926 12404
rect 21522 12348 21532 12404
rect 21588 12348 22764 12404
rect 22820 12348 22830 12404
rect 10658 12236 10668 12292
rect 10724 12236 12684 12292
rect 12740 12236 12750 12292
rect 15586 12236 15596 12292
rect 15652 12236 16380 12292
rect 16436 12236 16446 12292
rect 11666 12124 11676 12180
rect 11732 12124 14812 12180
rect 14868 12124 16940 12180
rect 16996 12124 17006 12180
rect 14242 12012 14252 12068
rect 14308 12012 15036 12068
rect 15092 12012 15102 12068
rect 15362 12012 15372 12068
rect 15428 12012 16828 12068
rect 16884 12012 16894 12068
rect 21970 12012 21980 12068
rect 22036 12012 22988 12068
rect 23044 12012 23054 12068
rect 25200 11956 26000 11984
rect 20850 11900 20860 11956
rect 20916 11900 22092 11956
rect 22148 11900 22158 11956
rect 24322 11900 24332 11956
rect 24388 11900 26000 11956
rect 25200 11872 26000 11900
rect 14690 11788 14700 11844
rect 14756 11788 15596 11844
rect 15652 11788 15662 11844
rect 19730 11788 19740 11844
rect 19796 11788 20300 11844
rect 20356 11788 21084 11844
rect 21140 11788 21150 11844
rect 4114 11732 4124 11788
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4388 11732 4398 11788
rect 9938 11732 9948 11788
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 10212 11732 10222 11788
rect 15762 11732 15772 11788
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 16036 11732 16046 11788
rect 21586 11732 21596 11788
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21860 11732 21870 11788
rect 4834 11676 4844 11732
rect 4900 11676 5964 11732
rect 6020 11676 6030 11732
rect 11218 11564 11228 11620
rect 11284 11564 14476 11620
rect 14532 11564 14542 11620
rect 3378 11452 3388 11508
rect 3444 11452 5516 11508
rect 5572 11452 6860 11508
rect 6916 11452 6926 11508
rect 11442 11340 11452 11396
rect 11508 11340 14924 11396
rect 14980 11340 15484 11396
rect 15540 11340 15550 11396
rect 20066 11340 20076 11396
rect 20132 11340 21420 11396
rect 21476 11340 21486 11396
rect 23538 11340 23548 11396
rect 23604 11340 24892 11396
rect 24948 11340 24958 11396
rect 6850 11228 6860 11284
rect 6916 11228 7868 11284
rect 7924 11228 9324 11284
rect 9380 11228 11340 11284
rect 11396 11228 11406 11284
rect 12674 11228 12684 11284
rect 12740 11228 13580 11284
rect 13636 11228 13646 11284
rect 20626 11228 20636 11284
rect 20692 11228 21980 11284
rect 22036 11228 23324 11284
rect 23380 11228 23390 11284
rect 7026 10948 7036 11004
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7300 10948 7310 11004
rect 12850 10948 12860 11004
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 13124 10948 13134 11004
rect 18674 10948 18684 11004
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18948 10948 18958 11004
rect 24498 10948 24508 11004
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24772 10948 24782 11004
rect 3490 10668 3500 10724
rect 3556 10668 4620 10724
rect 4676 10668 9772 10724
rect 9828 10668 9838 10724
rect 10210 10668 10220 10724
rect 10276 10668 10668 10724
rect 10724 10668 10734 10724
rect 2034 10556 2044 10612
rect 2100 10556 3276 10612
rect 3332 10556 4844 10612
rect 4900 10556 4910 10612
rect 8754 10556 8764 10612
rect 8820 10556 10444 10612
rect 10500 10556 10510 10612
rect 19618 10556 19628 10612
rect 19684 10556 21644 10612
rect 21700 10556 21710 10612
rect 20962 10444 20972 10500
rect 21028 10444 21532 10500
rect 21588 10444 21598 10500
rect 19506 10332 19516 10388
rect 19572 10332 20300 10388
rect 20356 10332 20636 10388
rect 20692 10332 20702 10388
rect 4114 10164 4124 10220
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4388 10164 4398 10220
rect 9938 10164 9948 10220
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 10212 10164 10222 10220
rect 15762 10164 15772 10220
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 16036 10164 16046 10220
rect 21586 10164 21596 10220
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21860 10164 21870 10220
rect 17378 10108 17388 10164
rect 17444 10108 21308 10164
rect 21364 10108 21374 10164
rect 10322 9996 10332 10052
rect 10388 9996 12012 10052
rect 12068 9996 12078 10052
rect 20962 9996 20972 10052
rect 21028 9996 23548 10052
rect 23604 9996 23614 10052
rect 25200 9940 26000 9968
rect 22754 9884 22764 9940
rect 22820 9884 26000 9940
rect 25200 9856 26000 9884
rect 18162 9660 18172 9716
rect 18228 9660 20188 9716
rect 20244 9660 20254 9716
rect 20626 9436 20636 9492
rect 20692 9436 21924 9492
rect 7026 9380 7036 9436
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7300 9380 7310 9436
rect 12850 9380 12860 9436
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 13124 9380 13134 9436
rect 18674 9380 18684 9436
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18948 9380 18958 9436
rect 21868 9380 21924 9436
rect 24498 9380 24508 9436
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24772 9380 24782 9436
rect 7410 9324 7420 9380
rect 7476 9324 7486 9380
rect 14802 9324 14812 9380
rect 14868 9324 15148 9380
rect 21858 9324 21868 9380
rect 21924 9324 23548 9380
rect 23604 9324 23614 9380
rect 7420 9268 7476 9324
rect 7186 9212 7196 9268
rect 7252 9212 7476 9268
rect 15092 9268 15148 9324
rect 15092 9212 16380 9268
rect 16436 9212 16446 9268
rect 20738 9212 20748 9268
rect 20804 9212 22764 9268
rect 22820 9212 22830 9268
rect 21410 9100 21420 9156
rect 21476 9100 21756 9156
rect 21812 9100 21822 9156
rect 12562 8988 12572 9044
rect 12628 8988 15372 9044
rect 15428 8988 15820 9044
rect 15876 8988 15886 9044
rect 21410 8988 21420 9044
rect 21476 8988 21644 9044
rect 21700 8988 23884 9044
rect 23940 8988 24220 9044
rect 24276 8988 24286 9044
rect 15474 8876 15484 8932
rect 15540 8876 16828 8932
rect 16884 8876 17388 8932
rect 17444 8876 17454 8932
rect 19842 8876 19852 8932
rect 19908 8876 20300 8932
rect 20356 8876 20636 8932
rect 20692 8876 20702 8932
rect 3154 8764 3164 8820
rect 3220 8764 4844 8820
rect 4900 8764 4910 8820
rect 20178 8764 20188 8820
rect 20244 8764 22036 8820
rect 21186 8652 21196 8708
rect 21252 8652 21476 8708
rect 4114 8596 4124 8652
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4388 8596 4398 8652
rect 9938 8596 9948 8652
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 10212 8596 10222 8652
rect 15762 8596 15772 8652
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 16036 8596 16046 8652
rect 21420 8484 21476 8652
rect 21586 8596 21596 8652
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21860 8596 21870 8652
rect 21420 8428 21644 8484
rect 21700 8428 21710 8484
rect 3714 8316 3724 8372
rect 3780 8316 6412 8372
rect 6468 8316 10332 8372
rect 10388 8316 10398 8372
rect 21980 8260 22036 8764
rect 22754 8428 22764 8484
rect 22820 8428 23436 8484
rect 23492 8428 23502 8484
rect 21970 8204 21980 8260
rect 22036 8204 22046 8260
rect 25200 7924 26000 7952
rect 24892 7868 26000 7924
rect 7026 7812 7036 7868
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7300 7812 7310 7868
rect 12850 7812 12860 7868
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 13124 7812 13134 7868
rect 18674 7812 18684 7868
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18948 7812 18958 7868
rect 24498 7812 24508 7868
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24772 7812 24782 7868
rect 10434 7756 10444 7812
rect 10500 7756 10836 7812
rect 10780 7700 10836 7756
rect 24892 7700 24948 7868
rect 25200 7840 26000 7868
rect 7756 7644 10556 7700
rect 10612 7644 10622 7700
rect 10780 7644 12852 7700
rect 21410 7644 21420 7700
rect 21476 7644 21532 7700
rect 21588 7644 21598 7700
rect 22642 7644 22652 7700
rect 22708 7644 24948 7700
rect 4946 7532 4956 7588
rect 5012 7532 5852 7588
rect 5908 7532 5918 7588
rect 6626 7532 6636 7588
rect 6692 7532 7196 7588
rect 7252 7532 7262 7588
rect 7756 7476 7812 7644
rect 12796 7588 12852 7644
rect 8306 7532 8316 7588
rect 8372 7532 9212 7588
rect 9268 7532 9278 7588
rect 11106 7532 11116 7588
rect 11172 7532 12012 7588
rect 12068 7532 12078 7588
rect 12786 7532 12796 7588
rect 12852 7532 15596 7588
rect 15652 7532 15662 7588
rect 4834 7420 4844 7476
rect 4900 7420 5628 7476
rect 5684 7420 7756 7476
rect 7812 7420 7822 7476
rect 9650 7420 9660 7476
rect 9716 7420 10332 7476
rect 10388 7420 10398 7476
rect 20066 7420 20076 7476
rect 20132 7420 22204 7476
rect 22260 7420 23324 7476
rect 23380 7420 23390 7476
rect 10994 7308 11004 7364
rect 11060 7308 13916 7364
rect 13972 7308 16268 7364
rect 16324 7308 16334 7364
rect 4722 7196 4732 7252
rect 4788 7196 5516 7252
rect 5572 7196 5582 7252
rect 4114 7028 4124 7084
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4388 7028 4398 7084
rect 9938 7028 9948 7084
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 10212 7028 10222 7084
rect 15762 7028 15772 7084
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 16036 7028 16046 7084
rect 21586 7028 21596 7084
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21860 7028 21870 7084
rect 23202 6748 23212 6804
rect 23268 6748 24220 6804
rect 24276 6748 24286 6804
rect 8306 6636 8316 6692
rect 8372 6636 8876 6692
rect 8932 6636 8942 6692
rect 18274 6636 18284 6692
rect 18340 6636 20636 6692
rect 20692 6636 20702 6692
rect 20738 6524 20748 6580
rect 20804 6524 22092 6580
rect 22148 6524 22158 6580
rect 12114 6412 12124 6468
rect 12180 6412 13468 6468
rect 13524 6412 13534 6468
rect 7026 6244 7036 6300
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7300 6244 7310 6300
rect 12850 6244 12860 6300
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 13124 6244 13134 6300
rect 18674 6244 18684 6300
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18948 6244 18958 6300
rect 24498 6244 24508 6300
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24772 6244 24782 6300
rect 17826 6076 17836 6132
rect 17892 6076 18508 6132
rect 18564 6076 18574 6132
rect 18722 6076 18732 6132
rect 18788 6076 19740 6132
rect 19796 6076 19806 6132
rect 25200 5908 26000 5936
rect 14242 5852 14252 5908
rect 14308 5852 17052 5908
rect 17108 5852 17118 5908
rect 19954 5852 19964 5908
rect 20020 5852 20412 5908
rect 20468 5852 21980 5908
rect 22036 5852 22428 5908
rect 22484 5852 22494 5908
rect 24210 5852 24220 5908
rect 24276 5852 26000 5908
rect 25200 5824 26000 5852
rect 4114 5460 4124 5516
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4388 5460 4398 5516
rect 9938 5460 9948 5516
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 10212 5460 10222 5516
rect 15762 5460 15772 5516
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 16036 5460 16046 5516
rect 21586 5460 21596 5516
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21860 5460 21870 5516
rect 23650 5180 23660 5236
rect 23716 5180 24220 5236
rect 24276 5180 24286 5236
rect 7026 4676 7036 4732
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7300 4676 7310 4732
rect 12850 4676 12860 4732
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 13124 4676 13134 4732
rect 18674 4676 18684 4732
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18948 4676 18958 4732
rect 24498 4676 24508 4732
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24772 4676 24782 4732
rect 4114 3892 4124 3948
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4388 3892 4398 3948
rect 9938 3892 9948 3948
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 10212 3892 10222 3948
rect 15762 3892 15772 3948
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 16036 3892 16046 3948
rect 21586 3892 21596 3948
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21860 3892 21870 3948
rect 25200 3892 26000 3920
rect 24210 3836 24220 3892
rect 24276 3836 26000 3892
rect 25200 3808 26000 3836
rect 23426 3388 23436 3444
rect 23492 3388 23884 3444
rect 23940 3388 23950 3444
rect 7026 3108 7036 3164
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7300 3108 7310 3164
rect 12850 3108 12860 3164
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 13124 3108 13134 3164
rect 18674 3108 18684 3164
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18948 3108 18958 3164
rect 24498 3108 24508 3164
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24772 3108 24782 3164
rect 25200 1876 26000 1904
rect 23986 1820 23996 1876
rect 24052 1820 26000 1876
rect 25200 1792 26000 1820
<< via3 >>
rect 4124 22708 4180 22764
rect 4228 22708 4284 22764
rect 4332 22708 4388 22764
rect 9948 22708 10004 22764
rect 10052 22708 10108 22764
rect 10156 22708 10212 22764
rect 15772 22708 15828 22764
rect 15876 22708 15932 22764
rect 15980 22708 16036 22764
rect 21596 22708 21652 22764
rect 21700 22708 21756 22764
rect 21804 22708 21860 22764
rect 7036 21924 7092 21980
rect 7140 21924 7196 21980
rect 7244 21924 7300 21980
rect 12860 21924 12916 21980
rect 12964 21924 13020 21980
rect 13068 21924 13124 21980
rect 18684 21924 18740 21980
rect 18788 21924 18844 21980
rect 18892 21924 18948 21980
rect 24508 21924 24564 21980
rect 24612 21924 24668 21980
rect 24716 21924 24772 21980
rect 4124 21140 4180 21196
rect 4228 21140 4284 21196
rect 4332 21140 4388 21196
rect 9948 21140 10004 21196
rect 10052 21140 10108 21196
rect 10156 21140 10212 21196
rect 15772 21140 15828 21196
rect 15876 21140 15932 21196
rect 15980 21140 16036 21196
rect 21596 21140 21652 21196
rect 21700 21140 21756 21196
rect 21804 21140 21860 21196
rect 7036 20356 7092 20412
rect 7140 20356 7196 20412
rect 7244 20356 7300 20412
rect 12860 20356 12916 20412
rect 12964 20356 13020 20412
rect 13068 20356 13124 20412
rect 18684 20356 18740 20412
rect 18788 20356 18844 20412
rect 18892 20356 18948 20412
rect 24508 20356 24564 20412
rect 24612 20356 24668 20412
rect 24716 20356 24772 20412
rect 16604 20076 16660 20132
rect 4124 19572 4180 19628
rect 4228 19572 4284 19628
rect 4332 19572 4388 19628
rect 9948 19572 10004 19628
rect 10052 19572 10108 19628
rect 10156 19572 10212 19628
rect 15772 19572 15828 19628
rect 15876 19572 15932 19628
rect 15980 19572 16036 19628
rect 21596 19572 21652 19628
rect 21700 19572 21756 19628
rect 21804 19572 21860 19628
rect 7036 18788 7092 18844
rect 7140 18788 7196 18844
rect 7244 18788 7300 18844
rect 12860 18788 12916 18844
rect 12964 18788 13020 18844
rect 13068 18788 13124 18844
rect 18684 18788 18740 18844
rect 18788 18788 18844 18844
rect 18892 18788 18948 18844
rect 24508 18788 24564 18844
rect 24612 18788 24668 18844
rect 24716 18788 24772 18844
rect 4124 18004 4180 18060
rect 4228 18004 4284 18060
rect 4332 18004 4388 18060
rect 9948 18004 10004 18060
rect 10052 18004 10108 18060
rect 10156 18004 10212 18060
rect 15772 18004 15828 18060
rect 15876 18004 15932 18060
rect 15980 18004 16036 18060
rect 21596 18004 21652 18060
rect 21700 18004 21756 18060
rect 21804 18004 21860 18060
rect 7036 17220 7092 17276
rect 7140 17220 7196 17276
rect 7244 17220 7300 17276
rect 12860 17220 12916 17276
rect 12964 17220 13020 17276
rect 13068 17220 13124 17276
rect 18684 17220 18740 17276
rect 18788 17220 18844 17276
rect 18892 17220 18948 17276
rect 24508 17220 24564 17276
rect 24612 17220 24668 17276
rect 24716 17220 24772 17276
rect 23884 16828 23940 16884
rect 4124 16436 4180 16492
rect 4228 16436 4284 16492
rect 4332 16436 4388 16492
rect 9948 16436 10004 16492
rect 10052 16436 10108 16492
rect 10156 16436 10212 16492
rect 15772 16436 15828 16492
rect 15876 16436 15932 16492
rect 15980 16436 16036 16492
rect 21596 16436 21652 16492
rect 21700 16436 21756 16492
rect 21804 16436 21860 16492
rect 7036 15652 7092 15708
rect 7140 15652 7196 15708
rect 7244 15652 7300 15708
rect 12860 15652 12916 15708
rect 12964 15652 13020 15708
rect 13068 15652 13124 15708
rect 18684 15652 18740 15708
rect 18788 15652 18844 15708
rect 18892 15652 18948 15708
rect 24508 15652 24564 15708
rect 24612 15652 24668 15708
rect 24716 15652 24772 15708
rect 4124 14868 4180 14924
rect 4228 14868 4284 14924
rect 4332 14868 4388 14924
rect 9948 14868 10004 14924
rect 10052 14868 10108 14924
rect 10156 14868 10212 14924
rect 15772 14868 15828 14924
rect 15876 14868 15932 14924
rect 15980 14868 16036 14924
rect 21596 14868 21652 14924
rect 21700 14868 21756 14924
rect 21804 14868 21860 14924
rect 24220 14812 24276 14868
rect 23884 14252 23940 14308
rect 7036 14084 7092 14140
rect 7140 14084 7196 14140
rect 7244 14084 7300 14140
rect 12860 14084 12916 14140
rect 12964 14084 13020 14140
rect 13068 14084 13124 14140
rect 18684 14084 18740 14140
rect 18788 14084 18844 14140
rect 18892 14084 18948 14140
rect 24508 14084 24564 14140
rect 24612 14084 24668 14140
rect 24716 14084 24772 14140
rect 16604 13916 16660 13972
rect 4124 13300 4180 13356
rect 4228 13300 4284 13356
rect 4332 13300 4388 13356
rect 9948 13300 10004 13356
rect 10052 13300 10108 13356
rect 10156 13300 10212 13356
rect 15772 13300 15828 13356
rect 15876 13300 15932 13356
rect 15980 13300 16036 13356
rect 21596 13300 21652 13356
rect 21700 13300 21756 13356
rect 21804 13300 21860 13356
rect 24220 12572 24276 12628
rect 7036 12516 7092 12572
rect 7140 12516 7196 12572
rect 7244 12516 7300 12572
rect 12860 12516 12916 12572
rect 12964 12516 13020 12572
rect 13068 12516 13124 12572
rect 18684 12516 18740 12572
rect 18788 12516 18844 12572
rect 18892 12516 18948 12572
rect 24508 12516 24564 12572
rect 24612 12516 24668 12572
rect 24716 12516 24772 12572
rect 4124 11732 4180 11788
rect 4228 11732 4284 11788
rect 4332 11732 4388 11788
rect 9948 11732 10004 11788
rect 10052 11732 10108 11788
rect 10156 11732 10212 11788
rect 15772 11732 15828 11788
rect 15876 11732 15932 11788
rect 15980 11732 16036 11788
rect 21596 11732 21652 11788
rect 21700 11732 21756 11788
rect 21804 11732 21860 11788
rect 7036 10948 7092 11004
rect 7140 10948 7196 11004
rect 7244 10948 7300 11004
rect 12860 10948 12916 11004
rect 12964 10948 13020 11004
rect 13068 10948 13124 11004
rect 18684 10948 18740 11004
rect 18788 10948 18844 11004
rect 18892 10948 18948 11004
rect 24508 10948 24564 11004
rect 24612 10948 24668 11004
rect 24716 10948 24772 11004
rect 4124 10164 4180 10220
rect 4228 10164 4284 10220
rect 4332 10164 4388 10220
rect 9948 10164 10004 10220
rect 10052 10164 10108 10220
rect 10156 10164 10212 10220
rect 15772 10164 15828 10220
rect 15876 10164 15932 10220
rect 15980 10164 16036 10220
rect 21596 10164 21652 10220
rect 21700 10164 21756 10220
rect 21804 10164 21860 10220
rect 7036 9380 7092 9436
rect 7140 9380 7196 9436
rect 7244 9380 7300 9436
rect 12860 9380 12916 9436
rect 12964 9380 13020 9436
rect 13068 9380 13124 9436
rect 18684 9380 18740 9436
rect 18788 9380 18844 9436
rect 18892 9380 18948 9436
rect 24508 9380 24564 9436
rect 24612 9380 24668 9436
rect 24716 9380 24772 9436
rect 21420 8988 21476 9044
rect 4124 8596 4180 8652
rect 4228 8596 4284 8652
rect 4332 8596 4388 8652
rect 9948 8596 10004 8652
rect 10052 8596 10108 8652
rect 10156 8596 10212 8652
rect 15772 8596 15828 8652
rect 15876 8596 15932 8652
rect 15980 8596 16036 8652
rect 21596 8596 21652 8652
rect 21700 8596 21756 8652
rect 21804 8596 21860 8652
rect 7036 7812 7092 7868
rect 7140 7812 7196 7868
rect 7244 7812 7300 7868
rect 12860 7812 12916 7868
rect 12964 7812 13020 7868
rect 13068 7812 13124 7868
rect 18684 7812 18740 7868
rect 18788 7812 18844 7868
rect 18892 7812 18948 7868
rect 24508 7812 24564 7868
rect 24612 7812 24668 7868
rect 24716 7812 24772 7868
rect 21420 7644 21476 7700
rect 4124 7028 4180 7084
rect 4228 7028 4284 7084
rect 4332 7028 4388 7084
rect 9948 7028 10004 7084
rect 10052 7028 10108 7084
rect 10156 7028 10212 7084
rect 15772 7028 15828 7084
rect 15876 7028 15932 7084
rect 15980 7028 16036 7084
rect 21596 7028 21652 7084
rect 21700 7028 21756 7084
rect 21804 7028 21860 7084
rect 7036 6244 7092 6300
rect 7140 6244 7196 6300
rect 7244 6244 7300 6300
rect 12860 6244 12916 6300
rect 12964 6244 13020 6300
rect 13068 6244 13124 6300
rect 18684 6244 18740 6300
rect 18788 6244 18844 6300
rect 18892 6244 18948 6300
rect 24508 6244 24564 6300
rect 24612 6244 24668 6300
rect 24716 6244 24772 6300
rect 4124 5460 4180 5516
rect 4228 5460 4284 5516
rect 4332 5460 4388 5516
rect 9948 5460 10004 5516
rect 10052 5460 10108 5516
rect 10156 5460 10212 5516
rect 15772 5460 15828 5516
rect 15876 5460 15932 5516
rect 15980 5460 16036 5516
rect 21596 5460 21652 5516
rect 21700 5460 21756 5516
rect 21804 5460 21860 5516
rect 7036 4676 7092 4732
rect 7140 4676 7196 4732
rect 7244 4676 7300 4732
rect 12860 4676 12916 4732
rect 12964 4676 13020 4732
rect 13068 4676 13124 4732
rect 18684 4676 18740 4732
rect 18788 4676 18844 4732
rect 18892 4676 18948 4732
rect 24508 4676 24564 4732
rect 24612 4676 24668 4732
rect 24716 4676 24772 4732
rect 4124 3892 4180 3948
rect 4228 3892 4284 3948
rect 4332 3892 4388 3948
rect 9948 3892 10004 3948
rect 10052 3892 10108 3948
rect 10156 3892 10212 3948
rect 15772 3892 15828 3948
rect 15876 3892 15932 3948
rect 15980 3892 16036 3948
rect 21596 3892 21652 3948
rect 21700 3892 21756 3948
rect 21804 3892 21860 3948
rect 7036 3108 7092 3164
rect 7140 3108 7196 3164
rect 7244 3108 7300 3164
rect 12860 3108 12916 3164
rect 12964 3108 13020 3164
rect 13068 3108 13124 3164
rect 18684 3108 18740 3164
rect 18788 3108 18844 3164
rect 18892 3108 18948 3164
rect 24508 3108 24564 3164
rect 24612 3108 24668 3164
rect 24716 3108 24772 3164
<< metal4 >>
rect 4096 22764 4416 22796
rect 4096 22708 4124 22764
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4388 22708 4416 22764
rect 4096 21196 4416 22708
rect 4096 21140 4124 21196
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4388 21140 4416 21196
rect 4096 19628 4416 21140
rect 4096 19572 4124 19628
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4388 19572 4416 19628
rect 4096 18060 4416 19572
rect 4096 18004 4124 18060
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4388 18004 4416 18060
rect 4096 16492 4416 18004
rect 4096 16436 4124 16492
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4388 16436 4416 16492
rect 4096 14924 4416 16436
rect 4096 14868 4124 14924
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4388 14868 4416 14924
rect 4096 13356 4416 14868
rect 4096 13300 4124 13356
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4388 13300 4416 13356
rect 4096 11788 4416 13300
rect 4096 11732 4124 11788
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4388 11732 4416 11788
rect 4096 10220 4416 11732
rect 4096 10164 4124 10220
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4388 10164 4416 10220
rect 4096 8652 4416 10164
rect 4096 8596 4124 8652
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4388 8596 4416 8652
rect 4096 7084 4416 8596
rect 4096 7028 4124 7084
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4388 7028 4416 7084
rect 4096 5516 4416 7028
rect 4096 5460 4124 5516
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4388 5460 4416 5516
rect 4096 3948 4416 5460
rect 4096 3892 4124 3948
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4388 3892 4416 3948
rect 4096 3076 4416 3892
rect 7008 21980 7328 22796
rect 7008 21924 7036 21980
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7300 21924 7328 21980
rect 7008 20412 7328 21924
rect 7008 20356 7036 20412
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7300 20356 7328 20412
rect 7008 18844 7328 20356
rect 7008 18788 7036 18844
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7300 18788 7328 18844
rect 7008 17276 7328 18788
rect 7008 17220 7036 17276
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7300 17220 7328 17276
rect 7008 15708 7328 17220
rect 7008 15652 7036 15708
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7300 15652 7328 15708
rect 7008 14140 7328 15652
rect 7008 14084 7036 14140
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7300 14084 7328 14140
rect 7008 12572 7328 14084
rect 7008 12516 7036 12572
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7300 12516 7328 12572
rect 7008 11004 7328 12516
rect 7008 10948 7036 11004
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7300 10948 7328 11004
rect 7008 9436 7328 10948
rect 7008 9380 7036 9436
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7300 9380 7328 9436
rect 7008 7868 7328 9380
rect 7008 7812 7036 7868
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7300 7812 7328 7868
rect 7008 6300 7328 7812
rect 7008 6244 7036 6300
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7300 6244 7328 6300
rect 7008 4732 7328 6244
rect 7008 4676 7036 4732
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7300 4676 7328 4732
rect 7008 3164 7328 4676
rect 7008 3108 7036 3164
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7300 3108 7328 3164
rect 7008 3076 7328 3108
rect 9920 22764 10240 22796
rect 9920 22708 9948 22764
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 10212 22708 10240 22764
rect 9920 21196 10240 22708
rect 9920 21140 9948 21196
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 10212 21140 10240 21196
rect 9920 19628 10240 21140
rect 9920 19572 9948 19628
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 10212 19572 10240 19628
rect 9920 18060 10240 19572
rect 9920 18004 9948 18060
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 10212 18004 10240 18060
rect 9920 16492 10240 18004
rect 9920 16436 9948 16492
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 10212 16436 10240 16492
rect 9920 14924 10240 16436
rect 9920 14868 9948 14924
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 10212 14868 10240 14924
rect 9920 13356 10240 14868
rect 9920 13300 9948 13356
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 10212 13300 10240 13356
rect 9920 11788 10240 13300
rect 9920 11732 9948 11788
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 10212 11732 10240 11788
rect 9920 10220 10240 11732
rect 9920 10164 9948 10220
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 10212 10164 10240 10220
rect 9920 8652 10240 10164
rect 9920 8596 9948 8652
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 10212 8596 10240 8652
rect 9920 7084 10240 8596
rect 9920 7028 9948 7084
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 10212 7028 10240 7084
rect 9920 5516 10240 7028
rect 9920 5460 9948 5516
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 10212 5460 10240 5516
rect 9920 3948 10240 5460
rect 9920 3892 9948 3948
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 10212 3892 10240 3948
rect 9920 3076 10240 3892
rect 12832 21980 13152 22796
rect 12832 21924 12860 21980
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 13124 21924 13152 21980
rect 12832 20412 13152 21924
rect 12832 20356 12860 20412
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 13124 20356 13152 20412
rect 12832 18844 13152 20356
rect 12832 18788 12860 18844
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 13124 18788 13152 18844
rect 12832 17276 13152 18788
rect 12832 17220 12860 17276
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 13124 17220 13152 17276
rect 12832 15708 13152 17220
rect 12832 15652 12860 15708
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 13124 15652 13152 15708
rect 12832 14140 13152 15652
rect 12832 14084 12860 14140
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 13124 14084 13152 14140
rect 12832 12572 13152 14084
rect 12832 12516 12860 12572
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 13124 12516 13152 12572
rect 12832 11004 13152 12516
rect 12832 10948 12860 11004
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 13124 10948 13152 11004
rect 12832 9436 13152 10948
rect 12832 9380 12860 9436
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 13124 9380 13152 9436
rect 12832 7868 13152 9380
rect 12832 7812 12860 7868
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 13124 7812 13152 7868
rect 12832 6300 13152 7812
rect 12832 6244 12860 6300
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 13124 6244 13152 6300
rect 12832 4732 13152 6244
rect 12832 4676 12860 4732
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 13124 4676 13152 4732
rect 12832 3164 13152 4676
rect 12832 3108 12860 3164
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 13124 3108 13152 3164
rect 12832 3076 13152 3108
rect 15744 22764 16064 22796
rect 15744 22708 15772 22764
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 16036 22708 16064 22764
rect 15744 21196 16064 22708
rect 15744 21140 15772 21196
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 16036 21140 16064 21196
rect 15744 19628 16064 21140
rect 18656 21980 18976 22796
rect 18656 21924 18684 21980
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18948 21924 18976 21980
rect 18656 20412 18976 21924
rect 18656 20356 18684 20412
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18948 20356 18976 20412
rect 15744 19572 15772 19628
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 16036 19572 16064 19628
rect 15744 18060 16064 19572
rect 15744 18004 15772 18060
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 16036 18004 16064 18060
rect 15744 16492 16064 18004
rect 15744 16436 15772 16492
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 16036 16436 16064 16492
rect 15744 14924 16064 16436
rect 15744 14868 15772 14924
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 16036 14868 16064 14924
rect 15744 13356 16064 14868
rect 16604 20132 16660 20142
rect 16604 13972 16660 20076
rect 16604 13906 16660 13916
rect 18656 18844 18976 20356
rect 18656 18788 18684 18844
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18948 18788 18976 18844
rect 18656 17276 18976 18788
rect 18656 17220 18684 17276
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18948 17220 18976 17276
rect 18656 15708 18976 17220
rect 18656 15652 18684 15708
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18948 15652 18976 15708
rect 18656 14140 18976 15652
rect 18656 14084 18684 14140
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18948 14084 18976 14140
rect 15744 13300 15772 13356
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 16036 13300 16064 13356
rect 15744 11788 16064 13300
rect 15744 11732 15772 11788
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 16036 11732 16064 11788
rect 15744 10220 16064 11732
rect 15744 10164 15772 10220
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 16036 10164 16064 10220
rect 15744 8652 16064 10164
rect 15744 8596 15772 8652
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 16036 8596 16064 8652
rect 15744 7084 16064 8596
rect 15744 7028 15772 7084
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 16036 7028 16064 7084
rect 15744 5516 16064 7028
rect 15744 5460 15772 5516
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 16036 5460 16064 5516
rect 15744 3948 16064 5460
rect 15744 3892 15772 3948
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 16036 3892 16064 3948
rect 15744 3076 16064 3892
rect 18656 12572 18976 14084
rect 18656 12516 18684 12572
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18948 12516 18976 12572
rect 18656 11004 18976 12516
rect 18656 10948 18684 11004
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18948 10948 18976 11004
rect 18656 9436 18976 10948
rect 18656 9380 18684 9436
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18948 9380 18976 9436
rect 18656 7868 18976 9380
rect 21568 22764 21888 22796
rect 21568 22708 21596 22764
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21860 22708 21888 22764
rect 21568 21196 21888 22708
rect 21568 21140 21596 21196
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21860 21140 21888 21196
rect 21568 19628 21888 21140
rect 21568 19572 21596 19628
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21860 19572 21888 19628
rect 21568 18060 21888 19572
rect 21568 18004 21596 18060
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21860 18004 21888 18060
rect 21568 16492 21888 18004
rect 24480 21980 24800 22796
rect 24480 21924 24508 21980
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24772 21924 24800 21980
rect 24480 20412 24800 21924
rect 24480 20356 24508 20412
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24772 20356 24800 20412
rect 24480 18844 24800 20356
rect 24480 18788 24508 18844
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24772 18788 24800 18844
rect 24480 17276 24800 18788
rect 24480 17220 24508 17276
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24772 17220 24800 17276
rect 21568 16436 21596 16492
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21860 16436 21888 16492
rect 21568 14924 21888 16436
rect 21568 14868 21596 14924
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21860 14868 21888 14924
rect 21568 13356 21888 14868
rect 23884 16884 23940 16894
rect 23884 14308 23940 16828
rect 24480 15708 24800 17220
rect 24480 15652 24508 15708
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24772 15652 24800 15708
rect 23884 14242 23940 14252
rect 24220 14868 24276 14878
rect 21568 13300 21596 13356
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21860 13300 21888 13356
rect 21568 11788 21888 13300
rect 24220 12628 24276 14812
rect 24220 12562 24276 12572
rect 24480 14140 24800 15652
rect 24480 14084 24508 14140
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24772 14084 24800 14140
rect 24480 12572 24800 14084
rect 21568 11732 21596 11788
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21860 11732 21888 11788
rect 21568 10220 21888 11732
rect 21568 10164 21596 10220
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21860 10164 21888 10220
rect 18656 7812 18684 7868
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18948 7812 18976 7868
rect 18656 6300 18976 7812
rect 21420 9044 21476 9054
rect 21420 7700 21476 8988
rect 21420 7634 21476 7644
rect 21568 8652 21888 10164
rect 21568 8596 21596 8652
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21860 8596 21888 8652
rect 18656 6244 18684 6300
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18948 6244 18976 6300
rect 18656 4732 18976 6244
rect 18656 4676 18684 4732
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18948 4676 18976 4732
rect 18656 3164 18976 4676
rect 18656 3108 18684 3164
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18948 3108 18976 3164
rect 18656 3076 18976 3108
rect 21568 7084 21888 8596
rect 21568 7028 21596 7084
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21860 7028 21888 7084
rect 21568 5516 21888 7028
rect 21568 5460 21596 5516
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21860 5460 21888 5516
rect 21568 3948 21888 5460
rect 21568 3892 21596 3948
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21860 3892 21888 3948
rect 21568 3076 21888 3892
rect 24480 12516 24508 12572
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24772 12516 24800 12572
rect 24480 11004 24800 12516
rect 24480 10948 24508 11004
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24772 10948 24800 11004
rect 24480 9436 24800 10948
rect 24480 9380 24508 9436
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24772 9380 24800 9436
rect 24480 7868 24800 9380
rect 24480 7812 24508 7868
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24772 7812 24800 7868
rect 24480 6300 24800 7812
rect 24480 6244 24508 6300
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24772 6244 24800 6300
rect 24480 4732 24800 6244
rect 24480 4676 24508 4732
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24772 4676 24800 4732
rect 24480 3164 24800 4676
rect 24480 3108 24508 3164
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24772 3108 24800 3164
rect 24480 3076 24800 3108
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _177_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12432 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _178_
timestamp 1698431365
transform 1 0 11424 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11648 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _181_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _182_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14672 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _183_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20272 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1698431365
transform -1 0 16800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16688 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _186_
timestamp 1698431365
transform 1 0 17808 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _188_
timestamp 1698431365
transform -1 0 22960 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _189_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698431365
transform 1 0 20272 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _191_
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _192_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _193_
timestamp 1698431365
transform 1 0 21280 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _194_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698431365
transform 1 0 21168 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _196_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22400 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _197_
timestamp 1698431365
transform -1 0 20272 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _198_
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1698431365
transform -1 0 17920 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _200_
timestamp 1698431365
transform -1 0 17920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _201_
timestamp 1698431365
transform -1 0 20160 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _202_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19488 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _203_
timestamp 1698431365
transform 1 0 16240 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _204_
timestamp 1698431365
transform 1 0 17808 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _206_
timestamp 1698431365
transform -1 0 20048 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _207_
timestamp 1698431365
transform -1 0 18704 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _208_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _209_
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _210_
timestamp 1698431365
transform -1 0 21840 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _211_
timestamp 1698431365
transform -1 0 22400 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _212_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _213_
timestamp 1698431365
transform -1 0 19712 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _214_
timestamp 1698431365
transform -1 0 20832 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _215_
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _216_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _217_
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _218_
timestamp 1698431365
transform -1 0 21840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _219_
timestamp 1698431365
transform -1 0 20160 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _220_
timestamp 1698431365
transform -1 0 17024 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _221_
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _222_
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _223_
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _224_
timestamp 1698431365
transform 1 0 21504 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _225_
timestamp 1698431365
transform -1 0 22960 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _226_
timestamp 1698431365
transform -1 0 20832 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _227_
timestamp 1698431365
transform -1 0 17696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _228_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _229_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _230_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _231_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14896 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _232_
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _233_
timestamp 1698431365
transform 1 0 15680 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _234_
timestamp 1698431365
transform 1 0 15568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _235_
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _236_
timestamp 1698431365
transform -1 0 15904 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _237_
timestamp 1698431365
transform 1 0 15344 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _238_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15232 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _239_
timestamp 1698431365
transform -1 0 15344 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _240_
timestamp 1698431365
transform -1 0 13888 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _241_
timestamp 1698431365
transform -1 0 15456 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _242_
timestamp 1698431365
transform -1 0 14672 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _243_
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _244_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14000 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _245_
timestamp 1698431365
transform 1 0 13664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _246_
timestamp 1698431365
transform -1 0 15680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _247_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15232 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _248_
timestamp 1698431365
transform -1 0 13664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _249_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _250_
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _251_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _252_
timestamp 1698431365
transform -1 0 12208 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _253_
timestamp 1698431365
transform -1 0 24304 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _254_
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _255_
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _256_
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _257_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24416 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _258_
timestamp 1698431365
transform 1 0 22960 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _259_
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _260_
timestamp 1698431365
transform -1 0 24080 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _261_
timestamp 1698431365
transform -1 0 23856 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _262_
timestamp 1698431365
transform 1 0 22400 0 1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _263_
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _264_
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _265_
timestamp 1698431365
transform -1 0 24304 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _266_
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _267_
timestamp 1698431365
transform 1 0 22400 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _268_
timestamp 1698431365
transform 1 0 13664 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _269_
timestamp 1698431365
transform 1 0 14112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _270_
timestamp 1698431365
transform 1 0 14560 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _271_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24304 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _272_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11536 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _273_
timestamp 1698431365
transform -1 0 8736 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _274_
timestamp 1698431365
transform 1 0 7728 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _275_
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _276_
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _277_
timestamp 1698431365
transform 1 0 6496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _278_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9744 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _279_
timestamp 1698431365
transform -1 0 9632 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _280_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _281_
timestamp 1698431365
transform 1 0 9184 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _282_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10752 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _283_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _284_
timestamp 1698431365
transform 1 0 11760 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _285_
timestamp 1698431365
transform 1 0 10304 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _286_
timestamp 1698431365
transform -1 0 8288 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _287_
timestamp 1698431365
transform 1 0 6608 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _288_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5152 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _289_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4592 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _290_
timestamp 1698431365
transform -1 0 9072 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _291_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7504 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _292_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _293_
timestamp 1698431365
transform 1 0 1792 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _294_
timestamp 1698431365
transform -1 0 13104 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _295_
timestamp 1698431365
transform -1 0 6608 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _296_
timestamp 1698431365
transform 1 0 10528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _297_
timestamp 1698431365
transform 1 0 7504 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _298_
timestamp 1698431365
transform 1 0 9744 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _299_
timestamp 1698431365
transform -1 0 10192 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _300_
timestamp 1698431365
transform 1 0 11088 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _301_
timestamp 1698431365
transform -1 0 11760 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _302_
timestamp 1698431365
transform -1 0 4592 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _303_
timestamp 1698431365
transform 1 0 3248 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _304_
timestamp 1698431365
transform -1 0 4032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _305_
timestamp 1698431365
transform 1 0 3584 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _306_
timestamp 1698431365
transform 1 0 4144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _307_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8624 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _308_
timestamp 1698431365
transform -1 0 7952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _309_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4592 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _310_
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _311_
timestamp 1698431365
transform 1 0 6160 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _312_
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _313_
timestamp 1698431365
transform 1 0 4928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _314_
timestamp 1698431365
transform 1 0 6048 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _315_
timestamp 1698431365
transform -1 0 3136 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _316_
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _317_
timestamp 1698431365
transform -1 0 7392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _318_
timestamp 1698431365
transform -1 0 3248 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _319_
timestamp 1698431365
transform 1 0 2912 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _320_
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _321_
timestamp 1698431365
transform 1 0 1904 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _322_
timestamp 1698431365
transform -1 0 3360 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _323_
timestamp 1698431365
transform -1 0 2240 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _324_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3360 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _325_
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _326_
timestamp 1698431365
transform 1 0 6048 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _327_
timestamp 1698431365
transform 1 0 6832 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _328_
timestamp 1698431365
transform -1 0 16688 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _329_
timestamp 1698431365
transform 1 0 12208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _330_
timestamp 1698431365
transform -1 0 11536 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _331_
timestamp 1698431365
transform -1 0 22400 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _332_
timestamp 1698431365
transform 1 0 15232 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _333_
timestamp 1698431365
transform 1 0 15904 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _334_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _335_
timestamp 1698431365
transform -1 0 12880 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _336_
timestamp 1698431365
transform -1 0 11088 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _337_
timestamp 1698431365
transform -1 0 16128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _338_
timestamp 1698431365
transform -1 0 10752 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _339_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _340_
timestamp 1698431365
transform 1 0 8288 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _341_
timestamp 1698431365
transform -1 0 12096 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _342_
timestamp 1698431365
transform 1 0 4256 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _343_
timestamp 1698431365
transform 1 0 2912 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _344_
timestamp 1698431365
transform 1 0 2016 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _345_
timestamp 1698431365
transform 1 0 3584 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _346_
timestamp 1698431365
transform 1 0 2576 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _347_
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _348_
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _349_
timestamp 1698431365
transform 1 0 5264 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _350_
timestamp 1698431365
transform -1 0 4928 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _351_
timestamp 1698431365
transform 1 0 9744 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _352_
timestamp 1698431365
transform 1 0 8624 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _353_
timestamp 1698431365
transform -1 0 8512 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _354_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _355_
timestamp 1698431365
transform 1 0 8960 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _356_
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _357_
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _358_
timestamp 1698431365
transform 1 0 3136 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _359_
timestamp 1698431365
transform 1 0 6832 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _360_
timestamp 1698431365
transform -1 0 14448 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _361_
timestamp 1698431365
transform -1 0 15680 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _362_
timestamp 1698431365
transform 1 0 16912 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _363_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _364_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _365_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _366_
timestamp 1698431365
transform 1 0 17360 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _367_
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _368_
timestamp 1698431365
transform 1 0 20160 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _369_
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _370_
timestamp 1698431365
transform -1 0 23856 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _371_
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _372_
timestamp 1698431365
transform 1 0 17808 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _373_
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _374_
timestamp 1698431365
transform 1 0 15456 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _375_
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _376_
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _377_
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _378_
timestamp 1698431365
transform 1 0 7504 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _379_
timestamp 1698431365
transform -1 0 17360 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _380_
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _381_
timestamp 1698431365
transform 1 0 11536 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _382_
timestamp 1698431365
transform 1 0 10864 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _383_
timestamp 1698431365
transform 1 0 12768 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _384_
timestamp 1698431365
transform 1 0 9520 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _385_
timestamp 1698431365
transform 1 0 7728 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _386_
timestamp 1698431365
transform 1 0 5712 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _387_
timestamp 1698431365
transform 1 0 1792 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _388_
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _389_
timestamp 1698431365
transform 1 0 6608 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _390_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _391_
timestamp 1698431365
transform 1 0 4592 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__CLK $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__CLK
timestamp 1698431365
transform 1 0 22736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__CLK
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__CLK
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__CLK
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__CLK
timestamp 1698431365
transform 1 0 19376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__CLK
timestamp 1698431365
transform -1 0 18816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__CLK
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__CLK
timestamp 1698431365
transform -1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__CLK
timestamp 1698431365
transform 1 0 16240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 11200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 23520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 19264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 23744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 22736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 22848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 24304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 20272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 23744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11424 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 11648 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1698431365
transform 1 0 7168 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 15344 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_188 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_174
timestamp 1698431365
transform 1 0 20832 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_190
timestamp 1698431365
transform 1 0 22624 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_45
timestamp 1698431365
transform 1 0 6384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_78
timestamp 1698431365
transform 1 0 10080 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_94
timestamp 1698431365
transform 1 0 11872 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_197
timestamp 1698431365
transform 1 0 23408 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_10
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_14
timestamp 1698431365
transform 1 0 2912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_45
timestamp 1698431365
transform 1 0 6384 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_61
timestamp 1698431365
transform 1 0 8176 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_117
timestamp 1698431365
transform 1 0 14448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_133
timestamp 1698431365
transform 1 0 16240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_157
timestamp 1698431365
transform 1 0 18928 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_174
timestamp 1698431365
transform 1 0 20832 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_182
timestamp 1698431365
transform 1 0 21728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_186
timestamp 1698431365
transform 1 0 22176 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_205
timestamp 1698431365
transform 1 0 24304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_18
timestamp 1698431365
transform 1 0 3360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_57
timestamp 1698431365
transform 1 0 7728 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_64
timestamp 1698431365
transform 1 0 8512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_80
timestamp 1698431365
transform 1 0 10304 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_88
timestamp 1698431365
transform 1 0 11200 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_98
timestamp 1698431365
transform 1 0 12320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_102
timestamp 1698431365
transform 1 0 12768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_65
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_105
timestamp 1698431365
transform 1 0 13104 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_109
timestamp 1698431365
transform 1 0 13552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_158
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_162
timestamp 1698431365
transform 1 0 19488 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_169
timestamp 1698431365
transform 1 0 20272 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_183
timestamp 1698431365
transform 1 0 21840 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_187
timestamp 1698431365
transform 1 0 22288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_203
timestamp 1698431365
transform 1 0 24080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_205
timestamp 1698431365
transform 1 0 24304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_31
timestamp 1698431365
transform 1 0 4816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_45
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_99
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_131
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_147
timestamp 1698431365
transform 1 0 17808 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_155
timestamp 1698431365
transform 1 0 18704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_159
timestamp 1698431365
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_205
timestamp 1698431365
transform 1 0 24304 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_10
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_41
timestamp 1698431365
transform 1 0 5936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_55
timestamp 1698431365
transform 1 0 7504 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_63
timestamp 1698431365
transform 1 0 8400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_87
timestamp 1698431365
transform 1 0 11088 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_96
timestamp 1698431365
transform 1 0 12096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_98
timestamp 1698431365
transform 1 0 12320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_188
timestamp 1698431365
transform 1 0 22400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_192
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_205
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_97
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_127
timestamp 1698431365
transform 1 0 15568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_143
timestamp 1698431365
transform 1 0 17360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_147
timestamp 1698431365
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_12
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_87
timestamp 1698431365
transform 1 0 11088 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_117
timestamp 1698431365
transform 1 0 14448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_119
timestamp 1698431365
transform 1 0 14672 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_122
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_171
timestamp 1698431365
transform 1 0 20496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_175
timestamp 1698431365
transform 1 0 20944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_177
timestamp 1698431365
transform 1 0 21168 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_186
timestamp 1698431365
transform 1 0 22176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_188
timestamp 1698431365
transform 1 0 22400 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_205
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_10
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_20
timestamp 1698431365
transform 1 0 3584 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_92
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_96
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_122
timestamp 1698431365
transform 1 0 15008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_124
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_33
timestamp 1698431365
transform 1 0 5040 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_37
timestamp 1698431365
transform 1 0 5488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_120
timestamp 1698431365
transform 1 0 14784 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_188
timestamp 1698431365
transform 1 0 22400 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_190
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_205
timestamp 1698431365
transform 1 0 24304 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_31
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_54
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_56
timestamp 1698431365
transform 1 0 7616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_86
timestamp 1698431365
transform 1 0 10976 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_111
timestamp 1698431365
transform 1 0 13776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_113
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_143
timestamp 1698431365
transform 1 0 17360 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_147
timestamp 1698431365
transform 1 0 17808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_149
timestamp 1698431365
transform 1 0 18032 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_162
timestamp 1698431365
transform 1 0 19488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_166
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_183
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_203
timestamp 1698431365
transform 1 0 24080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_205
timestamp 1698431365
transform 1 0 24304 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_30
timestamp 1698431365
transform 1 0 4704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_53
timestamp 1698431365
transform 1 0 7280 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_55
timestamp 1698431365
transform 1 0 7504 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_64
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_86
timestamp 1698431365
transform 1 0 10976 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_161
timestamp 1698431365
transform 1 0 19376 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_197
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_199
timestamp 1698431365
transform 1 0 23632 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_22
timestamp 1698431365
transform 1 0 3808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_24
timestamp 1698431365
transform 1 0 4032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_33
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_41
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_54
timestamp 1698431365
transform 1 0 7392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_84
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_92
timestamp 1698431365
transform 1 0 11648 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_96
timestamp 1698431365
transform 1 0 12096 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_120
timestamp 1698431365
transform 1 0 14784 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_132
timestamp 1698431365
transform 1 0 16128 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_197
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_4
timestamp 1698431365
transform 1 0 1792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_38
timestamp 1698431365
transform 1 0 5600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_42
timestamp 1698431365
transform 1 0 6048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_65
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_101
timestamp 1698431365
transform 1 0 12656 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_109
timestamp 1698431365
transform 1 0 13552 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_113
timestamp 1698431365
transform 1 0 14000 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_130
timestamp 1698431365
transform 1 0 15904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_148
timestamp 1698431365
transform 1 0 17920 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_164
timestamp 1698431365
transform 1 0 19712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_178
timestamp 1698431365
transform 1 0 21280 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_180
timestamp 1698431365
transform 1 0 21504 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_27
timestamp 1698431365
transform 1 0 4368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_49
timestamp 1698431365
transform 1 0 6832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_51
timestamp 1698431365
transform 1 0 7056 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_102
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_112
timestamp 1698431365
transform 1 0 13888 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_137
timestamp 1698431365
transform 1 0 16688 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_170
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_8
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_12
timestamp 1698431365
transform 1 0 2688 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_20
timestamp 1698431365
transform 1 0 3584 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_51
timestamp 1698431365
transform 1 0 7056 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698431365
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_84
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_205
timestamp 1698431365
transform 1 0 24304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_24
timestamp 1698431365
transform 1 0 4032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_29
timestamp 1698431365
transform 1 0 4592 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_33
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_55
timestamp 1698431365
transform 1 0 7504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_69
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_78
timestamp 1698431365
transform 1 0 10080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_82
timestamp 1698431365
transform 1 0 10528 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_91
timestamp 1698431365
transform 1 0 11536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_113
timestamp 1698431365
transform 1 0 14000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_119
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_142
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_146
timestamp 1698431365
transform 1 0 17696 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_153
timestamp 1698431365
transform 1 0 18480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_157
timestamp 1698431365
transform 1 0 18928 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_164
timestamp 1698431365
transform 1 0 19712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_166
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_193
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_197
timestamp 1698431365
transform 1 0 23408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_199
timestamp 1698431365
transform 1 0 23632 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_105
timestamp 1698431365
transform 1 0 13104 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_127
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_148
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_156
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_10
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_14
timestamp 1698431365
transform 1 0 2912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_16
timestamp 1698431365
transform 1 0 3136 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_67
timestamp 1698431365
transform 1 0 8848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_90
timestamp 1698431365
transform 1 0 11424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_128
timestamp 1698431365
transform 1 0 15680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_132
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_169
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_201
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_205
timestamp 1698431365
transform 1 0 24304 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_22
timestamp 1698431365
transform 1 0 3808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_24
timestamp 1698431365
transform 1 0 4032 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_34
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_42
timestamp 1698431365
transform 1 0 6048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_62
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_64
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_79
timestamp 1698431365
transform 1 0 10192 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_92
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_100
timestamp 1698431365
transform 1 0 12544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_118
timestamp 1698431365
transform 1 0 14560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_126
timestamp 1698431365
transform 1 0 15456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_152
timestamp 1698431365
transform 1 0 18368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_154
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_157
timestamp 1698431365
transform 1 0 18928 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_205
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_85
timestamp 1698431365
transform 1 0 10864 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_125
timestamp 1698431365
transform 1 0 15344 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_155
timestamp 1698431365
transform 1 0 18704 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_205
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_18
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_26
timestamp 1698431365
transform 1 0 4256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_30
timestamp 1698431365
transform 1 0 4704 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_131
timestamp 1698431365
transform 1 0 16016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_135
timestamp 1698431365
transform 1 0 16464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_205
timestamp 1698431365
transform 1 0 24304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_36
timestamp 1698431365
transform 1 0 5376 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_86
timestamp 1698431365
transform 1 0 10976 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_94
timestamp 1698431365
transform 1 0 11872 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_98
timestamp 1698431365
transform 1 0 12320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_110
timestamp 1698431365
transform 1 0 13664 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_126
timestamp 1698431365
transform 1 0 15456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_134
timestamp 1698431365
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_138
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_156
timestamp 1698431365
transform 1 0 18816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_160
timestamp 1698431365
transform 1 0 19264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 24416 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 24416 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 22288 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 20272 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 24416 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 22960 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 20832 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 13664 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_25 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 24640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_26
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_27
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 24640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_28
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_29
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_30
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_31
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 24640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_32
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_33
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 24640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_34
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_35
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 24640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_36
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_37
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 24640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_38
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_39
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_40
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_41
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 24640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_42
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_43
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 24640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 24640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer1
timestamp 1698431365
transform -1 0 10976 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer2
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer3
timestamp 1698431365
transform -1 0 24416 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer4
timestamp 1698431365
transform -1 0 24416 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_50 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_51
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_52
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_53
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_54
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_55
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_56
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_57
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_60
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_63
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_64
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_65
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_66
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_67
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_68
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_69
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_70
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_71
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_72
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_73
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_74
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_75
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_76
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_77
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_78
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_79
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_80
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_81
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_82
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_83
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_84
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_85
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_86
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_87
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_88
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_89
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_90
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_91
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_92
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_93
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_94
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_95
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_96
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_97
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_98
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_99
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_100
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_101
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_102
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_103
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_104
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_105
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_106
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_107
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_108
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_109
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_110
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_111
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_112
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_113
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_114
timestamp 1698431365
transform 1 0 8960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_115
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_116
timestamp 1698431365
transform 1 0 16576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_117
timestamp 1698431365
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_118
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 310 870
<< labels >>
flabel metal3 s 25200 1792 26000 1904 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 25200 21952 26000 22064 0 FreeSans 448 0 0 0 custom_settings[10]
port 1 nsew signal input
flabel metal3 s 25200 23968 26000 24080 0 FreeSans 448 0 0 0 custom_settings[11]
port 2 nsew signal input
flabel metal3 s 25200 3808 26000 3920 0 FreeSans 448 0 0 0 custom_settings[1]
port 3 nsew signal input
flabel metal3 s 25200 5824 26000 5936 0 FreeSans 448 0 0 0 custom_settings[2]
port 4 nsew signal input
flabel metal3 s 25200 7840 26000 7952 0 FreeSans 448 0 0 0 custom_settings[3]
port 5 nsew signal input
flabel metal3 s 25200 9856 26000 9968 0 FreeSans 448 0 0 0 custom_settings[4]
port 6 nsew signal input
flabel metal3 s 25200 11872 26000 11984 0 FreeSans 448 0 0 0 custom_settings[5]
port 7 nsew signal input
flabel metal3 s 25200 13888 26000 14000 0 FreeSans 448 0 0 0 custom_settings[6]
port 8 nsew signal input
flabel metal3 s 25200 15904 26000 16016 0 FreeSans 448 0 0 0 custom_settings[7]
port 9 nsew signal input
flabel metal3 s 25200 17920 26000 18032 0 FreeSans 448 0 0 0 custom_settings[8]
port 10 nsew signal input
flabel metal3 s 25200 19936 26000 20048 0 FreeSans 448 0 0 0 custom_settings[9]
port 11 nsew signal input
flabel metal2 s 21280 25200 21392 26000 0 FreeSans 448 90 0 0 io_out
port 12 nsew signal tristate
flabel metal2 s 12768 25200 12880 26000 0 FreeSans 448 90 0 0 rst_n
port 13 nsew signal input
flabel metal4 s 4096 3076 4416 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 9920 3076 10240 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 15744 3076 16064 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 21568 3076 21888 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 7008 3076 7328 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 12832 3076 13152 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 18656 3076 18976 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 24480 3076 24800 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal2 s 4256 25200 4368 26000 0 FreeSans 448 90 0 0 wb_clk_i
port 16 nsew signal input
rlabel metal1 12992 22736 12992 22736 0 vdd
rlabel via1 13072 21952 13072 21952 0 vss
rlabel metal2 8680 13664 8680 13664 0 _000_
rlabel metal2 6664 12488 6664 12488 0 _001_
rlabel metal2 3192 11760 3192 11760 0 _002_
rlabel metal2 2576 13048 2576 13048 0 _003_
rlabel metal2 7448 9128 7448 9128 0 _004_
rlabel metal2 12152 10920 12152 10920 0 _005_
rlabel metal2 9352 9576 9352 9576 0 _006_
rlabel metal2 2520 10304 2520 10304 0 _007_
rlabel metal2 2520 7896 2520 7896 0 _008_
rlabel metal2 4088 6216 4088 6216 0 _009_
rlabel metal2 7784 5824 7784 5824 0 _010_
rlabel metal2 13496 6216 13496 6216 0 _011_
rlabel metal2 14840 9128 14840 9128 0 _012_
rlabel metal3 18200 6104 18200 6104 0 _013_
rlabel metal2 20776 6664 20776 6664 0 _014_
rlabel metal2 18200 9408 18200 9408 0 _015_
rlabel metal2 22120 9072 22120 9072 0 _016_
rlabel metal2 18312 14168 18312 14168 0 _017_
rlabel metal2 18200 10248 18200 10248 0 _018_
rlabel metal2 21336 13216 21336 13216 0 _019_
rlabel metal2 20104 15680 20104 15680 0 _020_
rlabel metal3 21672 18312 21672 18312 0 _021_
rlabel metal2 17976 19600 17976 19600 0 _022_
rlabel metal2 20440 21168 20440 21168 0 _023_
rlabel metal2 20328 20160 20328 20160 0 _024_
rlabel metal2 16408 20272 16408 20272 0 _025_
rlabel metal2 2968 20412 2968 20412 0 _026_
rlabel metal2 5992 13888 5992 13888 0 _027_
rlabel metal2 2520 15960 2520 15960 0 _028_
rlabel metal2 6440 14112 6440 14112 0 _029_
rlabel metal2 16744 12600 16744 12600 0 _030_
rlabel metal2 16072 7784 16072 7784 0 _031_
rlabel metal2 12488 12992 12488 12992 0 _032_
rlabel metal2 13608 16520 13608 16520 0 _033_
rlabel metal2 13944 20832 13944 20832 0 _034_
rlabel metal3 11312 19432 11312 19432 0 _035_
rlabel metal2 9912 14336 9912 14336 0 _036_
rlabel metal2 5544 11088 5544 11088 0 _037_
rlabel metal2 23744 11480 23744 11480 0 _038_
rlabel metal2 24080 15960 24080 15960 0 _039_
rlabel metal2 24136 10080 24136 10080 0 _040_
rlabel metal2 23128 15596 23128 15596 0 _041_
rlabel metal2 22568 16352 22568 16352 0 _042_
rlabel metal2 23240 16352 23240 16352 0 _043_
rlabel metal2 16296 17136 16296 17136 0 _044_
rlabel metal2 14728 16912 14728 16912 0 _045_
rlabel metal2 16184 17024 16184 17024 0 _046_
rlabel metal2 23128 17472 23128 17472 0 _047_
rlabel metal2 10920 18480 10920 18480 0 _048_
rlabel metal2 10584 19880 10584 19880 0 _049_
rlabel metal3 9072 19096 9072 19096 0 _050_
rlabel metal2 10360 17472 10360 17472 0 _051_
rlabel metal2 7840 19992 7840 19992 0 _052_
rlabel metal2 8120 20496 8120 20496 0 _053_
rlabel metal2 8904 20608 8904 20608 0 _054_
rlabel metal2 9128 19600 9128 19600 0 _055_
rlabel metal2 9576 18256 9576 18256 0 _056_
rlabel metal2 10080 16744 10080 16744 0 _057_
rlabel metal3 8792 16968 8792 16968 0 _058_
rlabel metal2 2744 15736 2744 15736 0 _059_
rlabel metal2 12936 17976 12936 17976 0 _060_
rlabel metal2 9576 20048 9576 20048 0 _061_
rlabel metal2 7672 13832 7672 13832 0 _062_
rlabel metal2 5208 19320 5208 19320 0 _063_
rlabel metal2 4480 17640 4480 17640 0 _064_
rlabel metal2 8568 17864 8568 17864 0 _065_
rlabel metal3 4704 18424 4704 18424 0 _066_
rlabel metal2 2968 18368 2968 18368 0 _067_
rlabel metal2 16408 18592 16408 18592 0 _068_
rlabel metal2 3192 17584 3192 17584 0 _069_
rlabel metal2 11368 18816 11368 18816 0 _070_
rlabel metal3 8904 20552 8904 20552 0 _071_
rlabel metal2 10024 20160 10024 20160 0 _072_
rlabel metal2 11256 19936 11256 19936 0 _073_
rlabel metal2 11592 19264 11592 19264 0 _074_
rlabel metal3 7728 17080 7728 17080 0 _075_
rlabel metal3 5544 15288 5544 15288 0 _076_
rlabel metal2 4088 14504 4088 14504 0 _077_
rlabel metal2 3304 16408 3304 16408 0 _078_
rlabel metal2 4984 13720 4984 13720 0 _079_
rlabel metal2 7672 15680 7672 15680 0 _080_
rlabel metal2 6216 13776 6216 13776 0 _081_
rlabel metal2 6104 16576 6104 16576 0 _082_
rlabel metal3 5712 13496 5712 13496 0 _083_
rlabel metal2 6216 13048 6216 13048 0 _084_
rlabel metal2 2464 15288 2464 15288 0 _085_
rlabel metal2 6664 14280 6664 14280 0 _086_
rlabel metal2 3192 11256 3192 11256 0 _087_
rlabel metal2 7000 13552 7000 13552 0 _088_
rlabel metal2 2352 14280 2352 14280 0 _089_
rlabel metal2 2856 15008 2856 15008 0 _090_
rlabel metal2 3080 14504 3080 14504 0 _091_
rlabel metal2 6776 14840 6776 14840 0 _092_
rlabel metal2 7112 9128 7112 9128 0 _093_
rlabel metal2 11760 8120 11760 8120 0 _094_
rlabel metal3 11704 12264 11704 12264 0 _095_
rlabel metal2 14504 11424 14504 11424 0 _096_
rlabel metal3 16072 15288 16072 15288 0 _097_
rlabel metal2 16184 13216 16184 13216 0 _098_
rlabel metal2 14840 9520 14840 9520 0 _099_
rlabel metal3 13160 11256 13160 11256 0 _100_
rlabel metal2 10808 9744 10808 9744 0 _101_
rlabel metal2 12824 7504 12824 7504 0 _102_
rlabel metal2 6440 7896 6440 7896 0 _103_
rlabel metal2 9688 9296 9688 9296 0 _104_
rlabel metal3 5264 7448 5264 7448 0 _105_
rlabel metal2 4536 9968 4536 9968 0 _106_
rlabel metal2 2296 10752 2296 10752 0 _107_
rlabel metal2 3864 8400 3864 8400 0 _108_
rlabel metal2 2296 7924 2296 7924 0 _109_
rlabel metal3 6944 7560 6944 7560 0 _110_
rlabel metal2 4760 6944 4760 6944 0 _111_
rlabel metal2 9800 6888 9800 6888 0 _112_
rlabel metal3 8624 6664 8624 6664 0 _113_
rlabel metal2 12600 7784 12600 7784 0 _114_
rlabel metal2 11760 6664 11760 6664 0 _115_
rlabel metal2 15064 9100 15064 9100 0 _116_
rlabel metal2 15288 10976 15288 10976 0 _117_
rlabel metal2 19656 9408 19656 9408 0 _118_
rlabel metal2 15960 17808 15960 17808 0 _119_
rlabel metal2 20328 16744 20328 16744 0 _120_
rlabel metal2 18312 16268 18312 16268 0 _121_
rlabel metal2 22456 5936 22456 5936 0 _122_
rlabel metal2 20552 6160 20552 6160 0 _123_
rlabel metal3 20160 17416 20160 17416 0 _124_
rlabel metal2 20384 8456 20384 8456 0 _125_
rlabel metal2 20776 10136 20776 10136 0 _126_
rlabel metal2 21728 7336 21728 7336 0 _127_
rlabel metal3 20776 11368 20776 11368 0 _128_
rlabel metal2 20328 11984 20328 11984 0 _129_
rlabel metal2 16072 19880 16072 19880 0 _130_
rlabel metal3 17024 15400 17024 15400 0 _131_
rlabel metal2 20888 12096 20888 12096 0 _132_
rlabel metal3 17528 13048 17528 13048 0 _133_
rlabel metal2 17976 14000 17976 14000 0 _134_
rlabel metal2 19208 10920 19208 10920 0 _135_
rlabel metal2 18704 9688 18704 9688 0 _136_
rlabel metal2 21168 12040 21168 12040 0 _137_
rlabel metal2 22176 12264 22176 12264 0 _138_
rlabel metal3 20608 16072 20608 16072 0 _139_
rlabel metal2 20552 18032 20552 18032 0 _140_
rlabel metal3 19992 15288 19992 15288 0 _141_
rlabel metal2 20104 18704 20104 18704 0 _142_
rlabel metal3 21840 19432 21840 19432 0 _143_
rlabel metal2 21448 19376 21448 19376 0 _144_
rlabel metal2 19656 19600 19656 19600 0 _145_
rlabel metal2 16744 19600 16744 19600 0 _146_
rlabel metal2 20160 20664 20160 20664 0 _147_
rlabel metal2 22008 20328 22008 20328 0 _148_
rlabel metal2 20664 20384 20664 20384 0 _149_
rlabel metal3 17024 13944 17024 13944 0 _150_
rlabel metal2 16856 19824 16856 19824 0 _151_
rlabel metal2 16520 20720 16520 20720 0 _152_
rlabel metal3 16128 12040 16128 12040 0 _153_
rlabel metal2 15736 8400 15736 8400 0 _154_
rlabel metal2 14672 14728 14672 14728 0 _155_
rlabel metal2 15624 15568 15624 15568 0 _156_
rlabel metal2 15064 16016 15064 16016 0 _157_
rlabel metal2 13944 15960 13944 15960 0 _158_
rlabel metal2 15176 19376 15176 19376 0 _159_
rlabel metal2 15008 18200 15008 18200 0 _160_
rlabel metal2 14168 18480 14168 18480 0 _161_
rlabel metal2 14280 19320 14280 19320 0 _162_
rlabel metal3 15008 19208 15008 19208 0 _163_
rlabel metal2 12376 19096 12376 19096 0 _164_
rlabel metal2 12600 19488 12600 19488 0 _165_
rlabel metal2 9576 13664 9576 13664 0 _166_
rlabel metal2 15288 15148 15288 15148 0 _167_
rlabel metal2 22568 15512 22568 15512 0 _168_
rlabel metal2 22568 15204 22568 15204 0 _169_
rlabel metal2 23688 18144 23688 18144 0 _170_
rlabel metal2 24136 15260 24136 15260 0 _171_
rlabel metal2 24136 15624 24136 15624 0 _172_
rlabel metal2 24080 5992 24080 5992 0 _173_
rlabel metal2 24528 20664 24528 20664 0 _174_
rlabel metal2 22904 7840 22904 7840 0 _175_
rlabel metal2 22624 10696 22624 10696 0 _176_
rlabel metal2 22232 8176 22232 8176 0 baud_delay\[0\]
rlabel metal2 21896 20160 21896 20160 0 baud_delay\[10\]
rlabel metal3 22848 20776 22848 20776 0 baud_delay\[11\]
rlabel metal2 23240 6328 23240 6328 0 baud_delay\[1\]
rlabel metal2 21896 9240 21896 9240 0 baud_delay\[2\]
rlabel metal3 24080 9016 24080 9016 0 baud_delay\[3\]
rlabel metal3 22120 13720 22120 13720 0 baud_delay\[4\]
rlabel metal2 20328 10416 20328 10416 0 baud_delay\[5\]
rlabel metal2 21784 12096 21784 12096 0 baud_delay\[6\]
rlabel metal2 20216 16352 20216 16352 0 baud_delay\[7\]
rlabel metal2 22008 17920 22008 17920 0 baud_delay\[8\]
rlabel metal2 22120 19712 22120 19712 0 baud_delay\[9\]
rlabel metal2 10864 12152 10864 12152 0 char_at\[0\]
rlabel metal3 9632 10584 9632 10584 0 char_at\[1\]
rlabel metal2 4928 9016 4928 9016 0 char_at\[2\]
rlabel metal2 4200 7924 4200 7924 0 char_at\[3\]
rlabel metal2 7616 7448 7616 7448 0 char_at\[4\]
rlabel metal3 10024 7448 10024 7448 0 char_at\[5\]
rlabel metal2 11984 12040 11984 12040 0 char_at\[6\]
rlabel metal2 8288 19208 8288 19208 0 char_pointer\[0\]
rlabel metal2 8456 21112 8456 21112 0 char_pointer\[1\]
rlabel metal3 6216 18536 6216 18536 0 char_pointer\[2\]
rlabel metal2 10472 19096 10472 19096 0 char_pointer\[3\]
rlabel metal2 14952 12600 14952 12600 0 clknet_0_wb_clk_i
rlabel metal2 6944 5096 6944 5096 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 2296 21056 2296 21056 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 17080 6272 17080 6272 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 14896 10808 14896 10808 0 clknet_2_3__leaf_wb_clk_i
rlabel metal3 24626 1848 24626 1848 0 custom_settings[0]
rlabel metal2 20888 22232 20888 22232 0 custom_settings[10]
rlabel metal2 20160 22344 20160 22344 0 custom_settings[11]
rlabel metal2 24248 4088 24248 4088 0 custom_settings[1]
rlabel metal2 24248 5488 24248 5488 0 custom_settings[2]
rlabel metal3 23800 7672 23800 7672 0 custom_settings[3]
rlabel metal2 22792 9576 22792 9576 0 custom_settings[4]
rlabel metal2 24304 10808 24304 10808 0 custom_settings[5]
rlabel metal2 20552 13216 20552 13216 0 custom_settings[6]
rlabel metal2 23492 14616 23492 14616 0 custom_settings[7]
rlabel metal2 24136 18816 24136 18816 0 custom_settings[8]
rlabel metal3 23170 19992 23170 19992 0 custom_settings[9]
rlabel metal2 14560 14392 14560 14392 0 frame_counter\[0\]
rlabel metal2 14280 17192 14280 17192 0 frame_counter\[1\]
rlabel metal2 15288 19768 15288 19768 0 frame_counter\[2\]
rlabel metal2 12824 20104 12824 20104 0 frame_counter\[3\]
rlabel metal2 21336 23898 21336 23898 0 io_out
rlabel metal2 23632 3416 23632 3416 0 net1
rlabel metal2 22344 14224 22344 14224 0 net10
rlabel metal2 22400 17640 22400 17640 0 net11
rlabel metal2 21336 19656 21336 19656 0 net12
rlabel metal2 12040 20272 12040 20272 0 net13
rlabel metal2 18536 21280 18536 21280 0 net14
rlabel metal3 8176 18424 8176 18424 0 net15
rlabel metal2 8232 18424 8232 18424 0 net16
rlabel metal2 22008 16464 22008 16464 0 net17
rlabel metal2 23912 14728 23912 14728 0 net18
rlabel metal2 21112 22008 21112 22008 0 net2
rlabel metal2 20216 21840 20216 21840 0 net3
rlabel metal2 23744 5880 23744 5880 0 net4
rlabel metal2 23856 8232 23856 8232 0 net5
rlabel metal2 22792 8288 22792 8288 0 net6
rlabel metal2 21000 9632 21000 9632 0 net7
rlabel metal2 22568 12208 22568 12208 0 net8
rlabel metal2 20776 12880 20776 12880 0 net9
rlabel metal2 12768 22456 12768 22456 0 rst_n
rlabel metal2 14280 12712 14280 12712 0 uart_frame\[0\]
rlabel metal2 13944 11816 13944 11816 0 uart_frame\[1\]
rlabel metal2 10024 9520 10024 9520 0 uart_frame\[2\]
rlabel metal2 4648 10304 4648 10304 0 uart_frame\[3\]
rlabel metal2 4648 8372 4648 8372 0 uart_frame\[4\]
rlabel metal2 5880 6496 5880 6496 0 uart_frame\[5\]
rlabel metal2 9240 7224 9240 7224 0 uart_frame\[6\]
rlabel metal2 12040 7504 12040 7504 0 uart_frame\[7\]
rlabel metal2 11032 7728 11032 7728 0 uart_frame\[8\]
rlabel metal2 12600 8960 12600 8960 0 uart_frame\[9\]
rlabel metal3 6692 13944 6692 13944 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 26000 26000
<< end >>
