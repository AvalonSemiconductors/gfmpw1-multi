VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avali_logo
  CLASS BLOCK ;
  FOREIGN avali_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 293.500 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 94.000 201.500 107.500 202.000 ;
        RECT 89.000 201.000 114.000 201.500 ;
        RECT 85.000 200.500 119.000 201.000 ;
        RECT 82.500 200.000 122.500 200.500 ;
        RECT 80.000 199.500 122.500 200.000 ;
        RECT 77.500 199.000 122.000 199.500 ;
        RECT 75.500 198.500 122.000 199.000 ;
        RECT 74.000 198.000 121.500 198.500 ;
        RECT 72.000 197.500 121.500 198.000 ;
        RECT 70.500 197.000 121.000 197.500 ;
        RECT 69.000 196.500 121.000 197.000 ;
        RECT 67.500 196.000 120.500 196.500 ;
        RECT 66.000 195.500 120.000 196.000 ;
        RECT 65.000 195.000 120.000 195.500 ;
        RECT 63.500 194.500 119.500 195.000 ;
        RECT 62.500 194.000 119.500 194.500 ;
        RECT 61.000 193.500 119.000 194.000 ;
        RECT 60.000 193.000 119.000 193.500 ;
        RECT 59.000 192.500 118.500 193.000 ;
        RECT 58.000 192.000 118.500 192.500 ;
        RECT 57.000 191.500 118.000 192.000 ;
        RECT 56.000 191.000 118.000 191.500 ;
        RECT 55.000 190.500 117.500 191.000 ;
        RECT 54.000 190.000 117.500 190.500 ;
        RECT 53.000 189.500 117.000 190.000 ;
        RECT 52.000 189.000 116.500 189.500 ;
        RECT 51.000 188.500 116.500 189.000 ;
        RECT 50.000 188.000 116.000 188.500 ;
        RECT 49.500 187.500 116.000 188.000 ;
        RECT 48.500 187.000 115.500 187.500 ;
        RECT 48.000 186.500 115.500 187.000 ;
        RECT 47.000 186.000 115.000 186.500 ;
        RECT 46.000 185.500 115.000 186.000 ;
        RECT 45.500 185.000 114.500 185.500 ;
        RECT 44.500 184.500 114.500 185.000 ;
        RECT 44.000 184.000 93.000 184.500 ;
        RECT 110.500 184.000 114.000 184.500 ;
        RECT 43.000 183.500 89.000 184.000 ;
        RECT 42.500 183.000 86.000 183.500 ;
        RECT 42.000 182.500 83.500 183.000 ;
        RECT 41.000 182.000 81.500 182.500 ;
        RECT 40.500 181.500 79.500 182.000 ;
        RECT 40.000 181.000 77.500 181.500 ;
        RECT 39.000 180.500 76.000 181.000 ;
        RECT 38.500 180.000 74.500 180.500 ;
        RECT 38.000 179.500 73.000 180.000 ;
        RECT 37.000 179.000 71.500 179.500 ;
        RECT 36.500 178.500 70.500 179.000 ;
        RECT 36.000 178.000 69.000 178.500 ;
        RECT 35.500 177.500 68.000 178.000 ;
        RECT 35.000 177.000 67.000 177.500 ;
        RECT 34.500 176.500 65.500 177.000 ;
        RECT 33.500 176.000 64.500 176.500 ;
        RECT 33.000 175.500 63.500 176.000 ;
        RECT 32.500 175.000 62.500 175.500 ;
        RECT 32.000 174.500 61.500 175.000 ;
        RECT 31.500 174.000 61.000 174.500 ;
        RECT 31.000 173.500 60.000 174.000 ;
        RECT 30.500 173.000 59.000 173.500 ;
        RECT 30.000 172.500 58.000 173.000 ;
        RECT 29.500 172.000 57.500 172.500 ;
        RECT 29.000 171.500 56.500 172.000 ;
        RECT 28.500 171.000 56.000 171.500 ;
        RECT 28.000 170.500 55.000 171.000 ;
        RECT 27.500 170.000 54.000 170.500 ;
        RECT 27.000 169.500 53.500 170.000 ;
        RECT 26.500 169.000 53.000 169.500 ;
        RECT 26.000 168.500 52.000 169.000 ;
        RECT 26.000 168.000 51.500 168.500 ;
        RECT 25.500 167.500 50.500 168.000 ;
        RECT 25.000 167.000 50.000 167.500 ;
        RECT 24.500 166.500 49.500 167.000 ;
        RECT 24.000 166.000 49.000 166.500 ;
        RECT 23.500 165.500 48.000 166.000 ;
        RECT 23.000 165.000 47.500 165.500 ;
        RECT 23.000 164.500 47.000 165.000 ;
        RECT 22.500 164.000 46.500 164.500 ;
        RECT 22.000 163.500 46.000 164.000 ;
        RECT 21.500 163.000 45.500 163.500 ;
        RECT 21.000 162.500 44.500 163.000 ;
        RECT 21.000 162.000 44.000 162.500 ;
        RECT 20.500 161.500 43.500 162.000 ;
        RECT 20.000 161.000 43.000 161.500 ;
        RECT 19.500 160.500 42.500 161.000 ;
        RECT 19.500 160.000 42.000 160.500 ;
        RECT 19.000 159.500 41.500 160.000 ;
        RECT 18.500 159.000 41.000 159.500 ;
        RECT 18.500 158.500 40.500 159.000 ;
        RECT 18.000 158.000 40.000 158.500 ;
        RECT 17.500 157.500 39.500 158.000 ;
        RECT 17.000 156.500 39.000 157.500 ;
        RECT 16.500 156.000 38.500 156.500 ;
        RECT 16.500 155.500 38.000 156.000 ;
        RECT 16.000 155.000 37.500 155.500 ;
        RECT 15.500 154.500 37.000 155.000 ;
        RECT 15.500 154.000 36.500 154.500 ;
        RECT 15.000 153.500 36.000 154.000 ;
        RECT 14.500 153.000 36.000 153.500 ;
        RECT 14.500 152.500 35.500 153.000 ;
        RECT 14.000 152.000 35.000 152.500 ;
        RECT 14.000 151.500 34.500 152.000 ;
        RECT 13.500 151.000 34.500 151.500 ;
        RECT 13.000 150.500 34.000 151.000 ;
        RECT 13.000 150.000 33.500 150.500 ;
        RECT 12.500 149.000 33.000 150.000 ;
        RECT 12.000 148.500 32.500 149.000 ;
        RECT 12.000 148.000 32.000 148.500 ;
        RECT 11.500 147.500 32.000 148.000 ;
        RECT 11.500 147.000 31.500 147.500 ;
        RECT 11.000 146.000 31.000 147.000 ;
        RECT 10.500 145.500 30.500 146.000 ;
        RECT 10.500 145.000 30.000 145.500 ;
        RECT 10.000 144.500 30.000 145.000 ;
        RECT 10.000 144.000 29.500 144.500 ;
        RECT 9.500 143.000 29.000 144.000 ;
        RECT 9.000 142.000 28.500 143.000 ;
        RECT 8.500 141.000 28.000 142.000 ;
        RECT 8.500 140.500 27.500 141.000 ;
        RECT 8.000 140.000 27.500 140.500 ;
        RECT 8.000 139.500 27.000 140.000 ;
        RECT 7.500 139.000 27.000 139.500 ;
        RECT 7.500 138.500 26.500 139.000 ;
        RECT 7.000 138.000 26.500 138.500 ;
        RECT 7.000 137.000 26.000 138.000 ;
        RECT 6.500 136.000 25.500 137.000 ;
        RECT 6.500 135.500 25.000 136.000 ;
        RECT 6.000 135.000 25.000 135.500 ;
        RECT 6.000 134.500 24.500 135.000 ;
        RECT 5.500 134.000 24.500 134.500 ;
        RECT 5.500 133.000 24.000 134.000 ;
        RECT 5.000 131.500 23.500 133.000 ;
        RECT 4.500 130.000 23.000 131.500 ;
        RECT 4.500 129.500 22.500 130.000 ;
        RECT 4.000 129.000 22.500 129.500 ;
        RECT 4.000 128.000 22.000 129.000 ;
        RECT 3.500 127.500 22.000 128.000 ;
        RECT 3.500 126.000 21.500 127.500 ;
        RECT 3.000 124.000 21.000 126.000 ;
        RECT 2.500 122.500 20.500 124.000 ;
        RECT 2.500 121.500 20.000 122.500 ;
        RECT 2.000 120.500 20.000 121.500 ;
        RECT 2.000 119.000 19.500 120.500 ;
        RECT 1.500 118.000 19.500 119.000 ;
        RECT 1.500 116.000 19.000 118.000 ;
        RECT 1.000 115.500 19.000 116.000 ;
        RECT 1.000 112.500 18.500 115.500 ;
        RECT 0.500 112.000 18.500 112.500 ;
        RECT 0.500 107.500 18.000 112.000 ;
        RECT 0.500 106.500 17.500 107.500 ;
        RECT 0.000 95.500 17.500 106.500 ;
        RECT 0.500 94.500 17.500 95.500 ;
        RECT 0.500 89.500 18.000 94.500 ;
        RECT 1.000 86.500 18.500 89.500 ;
        RECT 1.000 86.000 19.000 86.500 ;
        RECT 1.500 84.000 19.000 86.000 ;
        RECT 1.500 83.000 19.500 84.000 ;
        RECT 2.000 81.500 19.500 83.000 ;
        RECT 2.000 80.000 20.000 81.500 ;
        RECT 2.500 79.500 20.000 80.000 ;
        RECT 2.500 78.000 20.500 79.500 ;
        RECT 3.000 76.000 21.000 78.000 ;
        RECT 3.500 74.500 21.500 76.000 ;
        RECT 3.500 74.000 22.000 74.500 ;
        RECT 4.000 73.000 22.000 74.000 ;
        RECT 4.000 72.500 22.500 73.000 ;
        RECT 4.500 72.000 22.500 72.500 ;
        RECT 4.500 70.500 23.000 72.000 ;
        RECT 5.000 69.000 23.500 70.500 ;
        RECT 5.500 68.000 24.000 69.000 ;
        RECT 5.500 67.500 24.500 68.000 ;
        RECT 6.000 67.000 24.500 67.500 ;
        RECT 6.000 66.500 25.000 67.000 ;
        RECT 6.500 66.000 25.000 66.500 ;
        RECT 6.500 65.000 25.500 66.000 ;
        RECT 7.000 64.500 25.500 65.000 ;
        RECT 7.000 63.500 26.000 64.500 ;
        RECT 7.500 62.500 26.500 63.500 ;
        RECT 8.000 61.500 27.000 62.500 ;
        RECT 8.000 61.000 27.500 61.500 ;
        RECT 8.500 60.000 28.000 61.000 ;
        RECT 9.000 59.000 28.500 60.000 ;
        RECT 9.500 58.000 29.000 59.000 ;
        RECT 10.000 57.500 29.500 58.000 ;
        RECT 10.000 57.000 30.000 57.500 ;
        RECT 10.500 56.500 30.000 57.000 ;
        RECT 10.500 56.000 30.500 56.500 ;
        RECT 11.000 55.000 31.000 56.000 ;
        RECT 11.500 54.000 31.500 55.000 ;
        RECT 12.000 53.500 32.000 54.000 ;
        RECT 12.000 53.000 32.500 53.500 ;
        RECT 12.500 52.000 33.000 53.000 ;
        RECT 13.000 51.500 33.500 52.000 ;
        RECT 13.000 51.000 34.000 51.500 ;
        RECT 13.500 50.500 34.000 51.000 ;
        RECT 14.000 50.000 34.500 50.500 ;
        RECT 14.000 49.500 35.000 50.000 ;
        RECT 14.500 49.000 35.500 49.500 ;
        RECT 14.500 48.500 36.000 49.000 ;
        RECT 15.000 48.000 36.000 48.500 ;
        RECT 15.500 47.500 36.500 48.000 ;
        RECT 15.500 47.000 37.000 47.500 ;
        RECT 16.000 46.500 37.500 47.000 ;
        RECT 16.000 46.000 38.000 46.500 ;
        RECT 16.500 45.500 38.500 46.000 ;
        RECT 17.000 45.000 38.500 45.500 ;
        RECT 17.000 44.500 39.000 45.000 ;
        RECT 17.500 44.000 39.500 44.500 ;
        RECT 18.000 43.500 40.000 44.000 ;
        RECT 18.000 43.000 40.500 43.500 ;
        RECT 18.500 42.500 41.000 43.000 ;
        RECT 19.000 42.000 41.500 42.500 ;
        RECT 19.500 41.500 42.000 42.000 ;
        RECT 19.500 41.000 42.500 41.500 ;
        RECT 20.000 40.500 43.000 41.000 ;
        RECT 20.500 40.000 43.500 40.500 ;
        RECT 21.000 39.500 44.000 40.000 ;
        RECT 21.000 39.000 44.500 39.500 ;
        RECT 21.500 38.500 45.000 39.000 ;
        RECT 22.000 38.000 46.000 38.500 ;
        RECT 22.500 37.500 46.500 38.000 ;
        RECT 22.500 37.000 47.000 37.500 ;
        RECT 23.000 36.500 47.500 37.000 ;
        RECT 23.500 36.000 48.000 36.500 ;
        RECT 24.000 35.500 48.500 36.000 ;
        RECT 24.500 35.000 49.500 35.500 ;
        RECT 25.000 34.500 50.000 35.000 ;
        RECT 25.500 34.000 50.500 34.500 ;
        RECT 25.500 33.500 51.000 34.000 ;
        RECT 26.000 33.000 52.000 33.500 ;
        RECT 26.500 32.500 52.500 33.000 ;
        RECT 27.000 32.000 53.000 32.500 ;
        RECT 27.500 31.500 54.000 32.000 ;
        RECT 28.000 31.000 54.500 31.500 ;
        RECT 28.500 30.500 55.500 31.000 ;
        RECT 29.000 30.000 56.000 30.500 ;
        RECT 29.500 29.500 57.000 30.000 ;
        RECT 30.000 29.000 57.500 29.500 ;
        RECT 30.500 28.500 58.500 29.000 ;
        RECT 31.000 28.000 59.500 28.500 ;
        RECT 31.500 27.500 60.500 28.000 ;
        RECT 32.000 27.000 61.500 27.500 ;
        RECT 32.500 26.500 61.500 27.000 ;
        RECT 33.000 26.000 61.500 26.500 ;
        RECT 33.500 25.500 61.500 26.000 ;
        RECT 34.000 25.000 61.500 25.500 ;
        RECT 35.000 24.500 61.500 25.000 ;
        RECT 35.500 24.000 61.500 24.500 ;
        RECT 36.000 23.500 61.500 24.000 ;
        RECT 36.500 23.000 61.500 23.500 ;
        RECT 37.000 22.500 61.000 23.000 ;
        RECT 38.000 22.000 61.000 22.500 ;
        RECT 38.500 21.500 61.000 22.000 ;
        RECT 39.000 21.000 61.000 21.500 ;
        RECT 39.500 20.500 61.000 21.000 ;
        RECT 40.500 20.000 61.000 20.500 ;
        RECT 41.000 19.500 61.000 20.000 ;
        RECT 41.500 19.000 61.000 19.500 ;
        RECT 42.500 18.500 61.000 19.000 ;
        RECT 43.000 18.000 60.500 18.500 ;
        RECT 44.000 17.500 60.500 18.000 ;
        RECT 44.500 17.000 60.500 17.500 ;
        RECT 45.000 16.500 60.500 17.000 ;
        RECT 46.000 16.000 60.500 16.500 ;
        RECT 47.000 15.500 60.500 16.000 ;
        RECT 47.500 15.000 60.500 15.500 ;
        RECT 48.500 14.500 60.500 15.000 ;
        RECT 49.000 14.000 60.000 14.500 ;
        RECT 50.000 13.500 60.000 14.000 ;
        RECT 51.000 13.000 60.000 13.500 ;
        RECT 51.500 12.500 60.000 13.000 ;
        RECT 52.500 12.000 60.000 12.500 ;
        RECT 53.500 11.500 60.000 12.000 ;
        RECT 54.500 11.000 60.000 11.500 ;
        RECT 55.500 10.500 60.000 11.000 ;
        RECT 56.000 10.000 59.500 10.500 ;
        RECT 57.000 9.500 59.500 10.000 ;
        RECT 58.000 9.000 59.500 9.500 ;
        RECT 59.000 8.500 59.500 9.000 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 196.000 292.500 197.000 293.000 ;
        RECT 195.500 292.000 197.000 292.500 ;
        RECT 195.000 291.000 197.000 292.000 ;
        RECT 194.500 290.500 197.500 291.000 ;
        RECT 194.000 290.000 197.500 290.500 ;
        RECT 193.500 289.500 197.500 290.000 ;
        RECT 193.000 289.000 197.500 289.500 ;
        RECT 192.500 288.000 198.000 289.000 ;
        RECT 192.000 287.500 198.000 288.000 ;
        RECT 191.500 287.000 198.500 287.500 ;
        RECT 191.000 286.500 198.500 287.000 ;
        RECT 190.500 285.500 198.500 286.500 ;
        RECT 190.000 285.000 199.000 285.500 ;
        RECT 189.500 284.500 199.000 285.000 ;
        RECT 189.000 284.000 199.000 284.500 ;
        RECT 188.500 283.500 199.000 284.000 ;
        RECT 188.000 282.500 199.500 283.500 ;
        RECT 187.500 282.000 199.500 282.500 ;
        RECT 187.000 281.500 199.500 282.000 ;
        RECT 186.500 281.000 200.000 281.500 ;
        RECT 186.000 280.000 200.000 281.000 ;
        RECT 185.500 279.500 200.000 280.000 ;
        RECT 185.000 279.000 200.500 279.500 ;
        RECT 184.500 278.500 200.500 279.000 ;
        RECT 184.000 277.500 200.500 278.500 ;
        RECT 183.500 277.000 201.000 277.500 ;
        RECT 183.000 276.500 201.000 277.000 ;
        RECT 182.500 276.000 201.000 276.500 ;
        RECT 182.000 275.500 201.000 276.000 ;
        RECT 182.000 275.000 201.500 275.500 ;
        RECT 181.500 274.500 201.500 275.000 ;
        RECT 181.000 274.000 201.500 274.500 ;
        RECT 180.500 273.500 201.500 274.000 ;
        RECT 180.000 273.000 201.500 273.500 ;
        RECT 180.000 272.500 202.000 273.000 ;
        RECT 179.500 272.000 202.000 272.500 ;
        RECT 179.000 271.500 202.000 272.000 ;
        RECT 178.500 271.000 202.000 271.500 ;
        RECT 178.000 270.500 202.000 271.000 ;
        RECT 178.000 270.000 202.500 270.500 ;
        RECT 177.500 269.500 202.500 270.000 ;
        RECT 177.000 269.000 202.500 269.500 ;
        RECT 176.500 268.500 202.500 269.000 ;
        RECT 176.000 268.000 202.500 268.500 ;
        RECT 176.000 267.500 203.000 268.000 ;
        RECT 175.500 267.000 203.000 267.500 ;
        RECT 175.000 266.500 203.000 267.000 ;
        RECT 174.500 266.000 203.000 266.500 ;
        RECT 174.000 265.000 203.000 266.000 ;
        RECT 173.500 264.500 203.000 265.000 ;
        RECT 173.000 264.000 203.500 264.500 ;
        RECT 172.500 263.500 203.500 264.000 ;
        RECT 172.000 262.500 203.500 263.500 ;
        RECT 171.500 262.000 203.500 262.500 ;
        RECT 171.000 261.500 203.500 262.000 ;
        RECT 170.500 260.500 203.500 261.500 ;
        RECT 170.000 260.000 203.500 260.500 ;
        RECT 169.500 259.500 203.500 260.000 ;
        RECT 169.000 259.000 203.500 259.500 ;
        RECT 168.500 258.000 203.500 259.000 ;
        RECT 168.000 257.500 204.000 258.000 ;
        RECT 167.500 257.000 204.000 257.500 ;
        RECT 167.000 256.000 204.000 257.000 ;
        RECT 166.500 255.500 204.000 256.000 ;
        RECT 166.000 255.000 203.500 255.500 ;
        RECT 165.500 254.000 203.500 255.000 ;
        RECT 165.000 253.500 203.500 254.000 ;
        RECT 164.500 253.000 203.500 253.500 ;
        RECT 164.000 252.500 203.500 253.000 ;
        RECT 163.500 251.500 203.500 252.500 ;
        RECT 163.000 251.000 203.500 251.500 ;
        RECT 162.500 250.500 203.500 251.000 ;
        RECT 162.000 249.500 203.500 250.500 ;
        RECT 161.500 249.000 203.000 249.500 ;
        RECT 161.000 248.500 203.000 249.000 ;
        RECT 160.500 247.500 203.000 248.500 ;
        RECT 160.000 247.000 203.000 247.500 ;
        RECT 159.500 246.500 203.000 247.000 ;
        RECT 159.000 245.500 202.500 246.500 ;
        RECT 158.500 245.000 202.500 245.500 ;
        RECT 158.000 244.500 202.500 245.000 ;
        RECT 157.500 243.500 202.500 244.500 ;
        RECT 157.000 243.000 202.000 243.500 ;
        RECT 156.500 242.500 202.000 243.000 ;
        RECT 156.000 241.500 202.000 242.500 ;
        RECT 155.500 241.000 201.500 241.500 ;
        RECT 155.000 240.000 201.500 241.000 ;
        RECT 154.500 239.500 201.500 240.000 ;
        RECT 154.000 239.000 201.000 239.500 ;
        RECT 153.500 238.000 201.000 239.000 ;
        RECT 153.000 237.500 201.000 238.000 ;
        RECT 152.500 237.000 200.500 237.500 ;
        RECT 152.000 236.000 200.500 237.000 ;
        RECT 151.500 235.500 200.500 236.000 ;
        RECT 151.000 234.500 200.000 235.500 ;
        RECT 150.500 234.000 200.000 234.500 ;
        RECT 150.000 233.500 199.500 234.000 ;
        RECT 149.500 232.500 199.500 233.500 ;
        RECT 149.000 232.000 199.000 232.500 ;
        RECT 148.500 231.000 199.000 232.000 ;
        RECT 148.000 230.500 199.000 231.000 ;
        RECT 147.500 230.000 198.500 230.500 ;
        RECT 147.000 229.000 198.500 230.000 ;
        RECT 146.500 228.500 198.000 229.000 ;
        RECT 146.000 227.500 198.000 228.500 ;
        RECT 145.500 227.000 197.500 227.500 ;
        RECT 145.000 226.000 197.500 227.000 ;
        RECT 144.500 225.500 197.000 226.000 ;
        RECT 144.000 224.500 197.000 225.500 ;
        RECT 143.500 224.000 196.500 224.500 ;
        RECT 143.000 223.500 196.500 224.000 ;
        RECT 142.500 223.000 196.500 223.500 ;
        RECT 142.500 222.500 196.000 223.000 ;
        RECT 142.000 222.000 196.000 222.500 ;
        RECT 141.500 221.500 196.000 222.000 ;
        RECT 141.500 221.000 195.500 221.500 ;
        RECT 141.000 220.500 195.500 221.000 ;
        RECT 140.500 220.000 195.500 220.500 ;
        RECT 140.500 219.500 195.000 220.000 ;
        RECT 140.000 219.000 195.000 219.500 ;
        RECT 139.500 218.500 195.000 219.000 ;
        RECT 139.500 218.000 194.500 218.500 ;
        RECT 139.000 217.500 194.500 218.000 ;
        RECT 138.500 217.000 194.500 217.500 ;
        RECT 138.500 216.500 194.000 217.000 ;
        RECT 138.000 216.000 194.000 216.500 ;
        RECT 137.500 215.000 193.500 216.000 ;
        RECT 137.000 214.500 193.500 215.000 ;
        RECT 136.500 213.500 193.000 214.500 ;
        RECT 136.000 213.000 193.000 213.500 ;
        RECT 136.000 212.500 192.500 213.000 ;
        RECT 135.500 212.000 192.500 212.500 ;
        RECT 135.000 211.000 192.000 212.000 ;
        RECT 134.500 210.500 192.000 211.000 ;
        RECT 134.000 209.500 191.500 210.500 ;
        RECT 133.500 209.000 191.500 209.500 ;
        RECT 133.000 208.000 191.000 209.000 ;
        RECT 132.500 207.000 190.500 208.000 ;
        RECT 132.000 206.500 190.500 207.000 ;
        RECT 131.500 205.500 190.000 206.500 ;
        RECT 131.000 205.000 190.000 205.500 ;
        RECT 130.500 204.000 189.500 205.000 ;
        RECT 130.000 203.000 189.000 204.000 ;
        RECT 129.500 202.500 189.000 203.000 ;
        RECT 129.000 201.500 188.500 202.500 ;
        RECT 128.500 200.500 188.000 201.500 ;
        RECT 128.000 200.000 188.000 200.500 ;
        RECT 127.500 199.000 187.500 200.000 ;
        RECT 127.000 198.000 187.000 199.000 ;
        RECT 126.500 197.500 187.000 198.000 ;
        RECT 126.000 196.500 186.500 197.500 ;
        RECT 125.500 195.500 186.000 196.500 ;
        RECT 125.000 195.000 186.000 195.500 ;
        RECT 124.500 194.000 185.500 195.000 ;
        RECT 124.000 193.000 185.000 194.000 ;
        RECT 123.500 192.500 185.000 193.000 ;
        RECT 123.500 192.000 184.500 192.500 ;
        RECT 123.000 191.500 184.500 192.000 ;
        RECT 123.000 191.000 184.000 191.500 ;
        RECT 122.500 190.500 184.000 191.000 ;
        RECT 122.000 190.000 184.000 190.500 ;
        RECT 122.000 189.500 183.500 190.000 ;
        RECT 121.500 189.000 183.500 189.500 ;
        RECT 121.500 188.500 183.000 189.000 ;
        RECT 121.000 188.000 183.000 188.500 ;
        RECT 121.000 187.500 182.500 188.000 ;
        RECT 120.500 186.500 182.500 187.500 ;
        RECT 120.000 186.000 182.000 186.500 ;
        RECT 119.500 185.500 182.000 186.000 ;
        RECT 119.500 185.000 181.500 185.500 ;
        RECT 119.000 184.000 181.500 185.000 ;
        RECT 118.500 183.000 181.000 184.000 ;
        RECT 118.000 182.000 180.500 183.000 ;
        RECT 117.500 181.000 180.000 182.000 ;
        RECT 117.000 180.500 180.000 181.000 ;
        RECT 117.000 180.000 179.500 180.500 ;
        RECT 116.500 179.500 179.500 180.000 ;
        RECT 116.500 179.000 179.000 179.500 ;
        RECT 116.000 178.000 179.000 179.000 ;
        RECT 115.500 177.000 178.500 178.000 ;
        RECT 115.000 176.000 178.000 177.000 ;
        RECT 114.500 175.000 177.500 176.000 ;
        RECT 114.000 174.500 177.500 175.000 ;
        RECT 114.000 174.000 177.000 174.500 ;
        RECT 113.500 173.500 177.000 174.000 ;
        RECT 113.500 173.000 176.500 173.500 ;
        RECT 113.000 172.500 176.500 173.000 ;
        RECT 113.000 172.000 176.000 172.500 ;
        RECT 112.500 171.000 176.000 172.000 ;
        RECT 112.000 170.000 175.500 171.000 ;
        RECT 111.500 169.000 175.000 170.000 ;
        RECT 111.000 168.000 174.500 169.000 ;
        RECT 110.500 167.500 174.500 168.000 ;
        RECT 110.500 167.000 174.000 167.500 ;
        RECT 110.000 166.500 174.000 167.000 ;
        RECT 110.000 165.500 173.500 166.500 ;
        RECT 109.500 164.500 173.000 165.500 ;
        RECT 109.000 164.000 173.000 164.500 ;
        RECT 109.000 163.500 172.500 164.000 ;
        RECT 108.500 163.000 172.500 163.500 ;
        RECT 108.500 162.500 172.000 163.000 ;
        RECT 108.000 162.000 172.000 162.500 ;
        RECT 108.000 161.000 171.500 162.000 ;
        RECT 107.500 160.500 171.000 161.000 ;
        RECT 107.500 160.000 170.500 160.500 ;
        RECT 107.000 159.500 170.000 160.000 ;
        RECT 107.000 159.000 169.500 159.500 ;
        RECT 106.500 158.500 169.000 159.000 ;
        RECT 106.500 158.000 168.500 158.500 ;
        RECT 106.000 157.500 168.000 158.000 ;
        RECT 106.000 157.000 167.500 157.500 ;
        RECT 106.000 156.500 167.000 157.000 ;
        RECT 105.500 156.000 166.500 156.500 ;
        RECT 105.500 155.500 166.000 156.000 ;
        RECT 105.000 155.000 165.500 155.500 ;
        RECT 105.000 154.500 165.000 155.000 ;
        RECT 105.000 154.000 164.500 154.500 ;
        RECT 104.500 153.500 164.000 154.000 ;
        RECT 104.500 153.000 163.500 153.500 ;
        RECT 104.000 152.500 163.000 153.000 ;
        RECT 104.000 152.000 162.500 152.500 ;
        RECT 103.500 151.500 162.000 152.000 ;
        RECT 103.500 151.000 161.500 151.500 ;
        RECT 103.500 150.500 161.000 151.000 ;
        RECT 103.000 149.500 160.500 150.500 ;
        RECT 102.500 149.000 160.000 149.500 ;
        RECT 102.500 148.500 159.500 149.000 ;
        RECT 102.500 148.000 159.000 148.500 ;
        RECT 102.000 147.500 158.500 148.000 ;
        RECT 102.000 147.000 158.000 147.500 ;
        RECT 101.500 146.500 157.500 147.000 ;
        RECT 101.500 146.000 157.000 146.500 ;
        RECT 101.500 145.500 156.500 146.000 ;
        RECT 101.000 145.000 156.000 145.500 ;
        RECT 101.000 144.500 155.500 145.000 ;
        RECT 100.500 144.000 155.000 144.500 ;
        RECT 100.500 143.500 154.500 144.000 ;
        RECT 100.500 143.000 154.000 143.500 ;
        RECT 100.000 142.500 153.500 143.000 ;
        RECT 100.000 142.000 153.000 142.500 ;
        RECT 99.500 141.500 152.500 142.000 ;
        RECT 99.500 141.000 152.000 141.500 ;
        RECT 99.500 140.500 151.500 141.000 ;
        RECT 99.000 140.000 151.000 140.500 ;
        RECT 99.000 139.500 150.500 140.000 ;
        RECT 99.000 139.000 150.000 139.500 ;
        RECT 98.500 138.500 149.500 139.000 ;
        RECT 98.500 138.000 149.000 138.500 ;
        RECT 98.000 137.500 148.500 138.000 ;
        RECT 98.000 137.000 148.000 137.500 ;
        RECT 98.000 136.500 147.500 137.000 ;
        RECT 97.500 136.000 147.000 136.500 ;
        RECT 97.500 135.500 146.500 136.000 ;
        RECT 97.500 135.000 146.000 135.500 ;
        RECT 97.000 134.500 146.000 135.000 ;
        RECT 97.000 134.000 145.500 134.500 ;
        RECT 96.500 133.500 145.000 134.000 ;
        RECT 96.500 133.000 144.500 133.500 ;
        RECT 96.500 132.500 144.000 133.000 ;
        RECT 96.000 132.000 143.500 132.500 ;
        RECT 96.000 131.500 143.000 132.000 ;
        RECT 96.000 131.000 142.500 131.500 ;
        RECT 95.500 130.500 142.000 131.000 ;
        RECT 95.500 130.000 141.500 130.500 ;
        RECT 95.500 129.500 141.000 130.000 ;
        RECT 95.000 129.000 140.500 129.500 ;
        RECT 95.000 128.500 140.000 129.000 ;
        RECT 94.500 127.500 139.500 128.500 ;
        RECT 94.500 127.000 139.000 127.500 ;
        RECT 94.000 126.500 138.500 127.000 ;
        RECT 94.000 126.000 138.000 126.500 ;
        RECT 94.000 125.500 137.500 126.000 ;
        RECT 93.500 125.000 137.000 125.500 ;
        RECT 93.500 124.500 136.500 125.000 ;
        RECT 93.500 124.000 136.000 124.500 ;
        RECT 93.000 123.500 136.000 124.000 ;
        RECT 93.000 123.000 135.500 123.500 ;
        RECT 93.000 122.500 135.000 123.000 ;
        RECT 92.500 122.000 134.500 122.500 ;
        RECT 92.500 121.500 134.000 122.000 ;
        RECT 92.500 121.000 133.500 121.500 ;
        RECT 92.000 120.000 133.000 121.000 ;
        RECT 92.000 119.500 132.500 120.000 ;
        RECT 91.500 119.000 132.000 119.500 ;
        RECT 91.500 118.500 131.500 119.000 ;
        RECT 91.500 118.000 131.000 118.500 ;
        RECT 91.000 117.000 130.500 118.000 ;
        RECT 91.000 116.500 130.000 117.000 ;
        RECT 90.500 116.000 129.500 116.500 ;
        RECT 90.500 115.500 129.000 116.000 ;
        RECT 90.500 115.000 128.500 115.500 ;
        RECT 90.000 114.000 128.000 115.000 ;
        RECT 90.000 113.500 127.500 114.000 ;
        RECT 89.500 113.000 127.000 113.500 ;
        RECT 89.500 112.500 126.500 113.000 ;
        RECT 89.500 111.500 126.000 112.500 ;
        RECT 89.000 111.000 125.500 111.500 ;
        RECT 89.000 110.500 125.000 111.000 ;
        RECT 89.000 110.000 124.500 110.500 ;
        RECT 88.500 109.500 124.500 110.000 ;
        RECT 88.500 109.000 124.000 109.500 ;
        RECT 88.500 108.500 123.500 109.000 ;
        RECT 88.000 108.000 123.000 108.500 ;
        RECT 88.000 107.000 122.500 108.000 ;
        RECT 87.500 106.500 122.000 107.000 ;
        RECT 87.500 106.000 121.500 106.500 ;
        RECT 87.500 105.500 121.000 106.000 ;
        RECT 87.000 105.000 121.000 105.500 ;
        RECT 87.000 104.500 120.500 105.000 ;
        RECT 87.000 104.000 120.000 104.500 ;
        RECT 87.000 103.500 119.500 104.000 ;
        RECT 86.500 103.000 119.500 103.500 ;
        RECT 86.500 102.500 119.000 103.000 ;
        RECT 86.500 102.000 118.500 102.500 ;
        RECT 86.000 101.000 118.000 102.000 ;
        RECT 86.000 100.500 117.500 101.000 ;
        RECT 85.500 100.000 117.000 100.500 ;
        RECT 85.500 99.000 116.500 100.000 ;
        RECT 85.500 98.500 116.000 99.000 ;
        RECT 85.000 97.500 115.500 98.500 ;
        RECT 85.000 97.000 115.000 97.500 ;
        RECT 84.500 96.500 114.500 97.000 ;
        RECT 84.500 95.500 114.000 96.500 ;
        RECT 84.500 95.000 113.500 95.500 ;
        RECT 84.000 94.500 113.000 95.000 ;
        RECT 84.000 93.500 112.500 94.500 ;
        RECT 83.500 93.000 112.000 93.500 ;
        RECT 83.500 92.000 111.500 93.000 ;
        RECT 83.000 91.500 111.000 92.000 ;
        RECT 83.000 91.000 110.500 91.500 ;
        RECT 83.000 90.000 110.000 91.000 ;
        RECT 82.500 89.500 109.500 90.000 ;
        RECT 82.500 89.000 109.000 89.500 ;
        RECT 82.500 88.500 108.500 89.000 ;
        RECT 82.000 88.000 108.500 88.500 ;
        RECT 82.000 87.500 108.000 88.000 ;
        RECT 82.000 86.500 107.500 87.500 ;
        RECT 81.500 86.000 107.000 86.500 ;
        RECT 81.500 85.000 106.500 86.000 ;
        RECT 81.000 84.500 106.000 85.000 ;
        RECT 81.000 84.000 105.500 84.500 ;
        RECT 81.000 83.000 105.000 84.000 ;
        RECT 80.500 82.500 104.500 83.000 ;
        RECT 80.500 81.500 104.000 82.500 ;
        RECT 80.000 81.000 103.500 81.500 ;
        RECT 80.000 80.000 103.000 81.000 ;
        RECT 80.000 79.500 102.500 80.000 ;
        RECT 79.500 78.500 102.000 79.500 ;
        RECT 79.500 78.000 101.500 78.500 ;
        RECT 79.000 77.000 101.000 78.000 ;
        RECT 79.000 76.500 100.500 77.000 ;
        RECT 79.000 76.000 100.000 76.500 ;
        RECT 78.500 75.500 100.000 76.000 ;
        RECT 78.500 75.000 99.500 75.500 ;
        RECT 78.500 74.500 99.000 75.000 ;
        RECT 78.000 74.000 99.000 74.500 ;
        RECT 78.000 73.500 98.500 74.000 ;
        RECT 78.000 72.500 98.000 73.500 ;
        RECT 77.500 72.000 97.500 72.500 ;
        RECT 77.500 71.000 97.000 72.000 ;
        RECT 77.000 70.500 96.500 71.000 ;
        RECT 77.000 69.500 96.000 70.500 ;
        RECT 77.000 69.000 95.500 69.500 ;
        RECT 76.500 68.000 95.000 69.000 ;
        RECT 76.500 67.500 94.500 68.000 ;
        RECT 76.500 67.000 94.000 67.500 ;
        RECT 76.000 66.500 94.000 67.000 ;
        RECT 76.000 65.500 93.500 66.500 ;
        RECT 76.000 65.000 93.000 65.500 ;
        RECT 75.500 64.000 92.500 65.000 ;
        RECT 75.500 63.500 92.000 64.000 ;
        RECT 75.000 63.000 92.000 63.500 ;
        RECT 75.000 62.500 91.500 63.000 ;
        RECT 75.000 61.500 91.000 62.500 ;
        RECT 74.500 61.000 90.500 61.500 ;
        RECT 74.500 60.000 90.000 61.000 ;
        RECT 74.500 59.500 89.500 60.000 ;
        RECT 74.000 59.000 89.500 59.500 ;
        RECT 74.000 58.000 89.000 59.000 ;
        RECT 74.000 57.500 88.500 58.000 ;
        RECT 73.500 56.500 88.000 57.500 ;
        RECT 73.500 55.500 87.500 56.500 ;
        RECT 73.000 54.500 87.000 55.500 ;
        RECT 73.000 54.000 86.500 54.500 ;
        RECT 73.000 53.500 86.000 54.000 ;
        RECT 72.500 53.000 86.000 53.500 ;
        RECT 72.500 52.000 85.500 53.000 ;
        RECT 72.500 51.500 85.000 52.000 ;
        RECT 72.000 51.000 85.000 51.500 ;
        RECT 72.000 50.000 84.500 51.000 ;
        RECT 72.000 49.000 84.000 50.000 ;
        RECT 71.500 48.500 83.500 49.000 ;
        RECT 71.500 47.500 83.000 48.500 ;
        RECT 71.500 47.000 82.500 47.500 ;
        RECT 71.000 46.500 82.500 47.000 ;
        RECT 71.000 45.500 82.000 46.500 ;
        RECT 71.000 44.500 81.500 45.500 ;
        RECT 70.500 43.500 81.000 44.500 ;
        RECT 70.500 42.500 80.500 43.500 ;
        RECT 70.000 41.500 80.000 42.500 ;
        RECT 70.000 40.500 79.500 41.500 ;
        RECT 70.000 40.000 79.000 40.500 ;
        RECT 69.500 39.500 79.000 40.000 ;
        RECT 69.500 38.500 78.500 39.500 ;
        RECT 69.500 37.500 78.000 38.500 ;
        RECT 69.000 36.500 77.500 37.500 ;
        RECT 69.000 35.500 77.000 36.500 ;
        RECT 69.000 35.000 76.500 35.500 ;
        RECT 68.500 34.500 76.500 35.000 ;
        RECT 68.500 33.500 76.000 34.500 ;
        RECT 68.500 33.000 75.500 33.500 ;
        RECT 68.000 32.500 75.500 33.000 ;
        RECT 68.000 31.500 75.000 32.500 ;
        RECT 68.000 30.500 74.500 31.500 ;
        RECT 67.500 29.500 74.000 30.500 ;
        RECT 67.500 28.500 73.500 29.500 ;
        RECT 67.500 27.500 73.000 28.500 ;
        RECT 67.000 26.500 72.500 27.500 ;
        RECT 67.000 25.500 72.000 26.500 ;
        RECT 67.000 25.000 71.500 25.500 ;
        RECT 66.500 24.500 71.500 25.000 ;
        RECT 66.500 23.500 71.000 24.500 ;
        RECT 66.500 22.500 70.500 23.500 ;
        RECT 66.000 21.500 70.000 22.500 ;
        RECT 66.000 20.500 69.500 21.500 ;
        RECT 66.000 20.000 69.000 20.500 ;
        RECT 65.500 19.500 69.000 20.000 ;
        RECT 65.500 18.500 68.500 19.500 ;
        RECT 65.500 17.500 68.000 18.500 ;
        RECT 65.000 17.000 68.000 17.500 ;
        RECT 65.000 16.000 67.500 17.000 ;
        RECT 65.000 15.000 67.000 16.000 ;
        RECT 65.000 14.500 66.500 15.000 ;
        RECT 64.500 14.000 66.500 14.500 ;
        RECT 64.500 13.000 66.000 14.000 ;
        RECT 64.500 12.000 65.500 13.000 ;
        RECT 64.000 11.000 65.000 12.000 ;
        RECT 64.000 10.000 64.500 11.000 ;
    END
  END vdd
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 250.000 293.500 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 250.000 293.500 ;
      LAYER Metal4 ;
        RECT 243.500 209.000 244.000 209.500 ;
        RECT 243.000 208.500 244.000 209.000 ;
        RECT 242.000 208.000 244.000 208.500 ;
        RECT 241.500 207.500 244.000 208.000 ;
        RECT 240.500 207.000 244.000 207.500 ;
        RECT 240.000 206.500 244.000 207.000 ;
        RECT 239.000 206.000 244.000 206.500 ;
        RECT 238.500 205.500 244.000 206.000 ;
        RECT 237.500 205.000 244.000 205.500 ;
        RECT 236.500 204.500 244.000 205.000 ;
        RECT 236.000 204.000 244.000 204.500 ;
        RECT 235.000 203.500 244.000 204.000 ;
        RECT 234.500 203.000 244.000 203.500 ;
        RECT 233.500 202.500 244.000 203.000 ;
        RECT 233.000 202.000 244.000 202.500 ;
        RECT 232.000 201.500 244.000 202.000 ;
        RECT 231.500 201.000 244.000 201.500 ;
        RECT 230.500 200.500 244.000 201.000 ;
        RECT 230.000 200.000 244.000 200.500 ;
        RECT 229.000 199.500 244.000 200.000 ;
        RECT 228.500 199.000 244.000 199.500 ;
        RECT 227.500 198.500 244.000 199.000 ;
        RECT 227.000 198.000 244.000 198.500 ;
        RECT 226.000 197.500 244.000 198.000 ;
        RECT 225.500 197.000 244.000 197.500 ;
        RECT 225.000 196.500 244.000 197.000 ;
        RECT 224.000 196.000 244.000 196.500 ;
        RECT 223.500 195.500 244.000 196.000 ;
        RECT 222.500 195.000 244.000 195.500 ;
        RECT 222.000 194.500 244.000 195.000 ;
        RECT 221.000 194.000 244.000 194.500 ;
        RECT 220.500 193.500 244.000 194.000 ;
        RECT 220.000 193.000 244.000 193.500 ;
        RECT 219.000 192.500 244.000 193.000 ;
        RECT 218.500 192.000 244.000 192.500 ;
        RECT 217.500 191.500 244.000 192.000 ;
        RECT 217.000 191.000 244.000 191.500 ;
        RECT 216.500 190.500 244.000 191.000 ;
        RECT 215.500 190.000 244.000 190.500 ;
        RECT 215.000 189.500 244.000 190.000 ;
        RECT 214.500 189.000 244.000 189.500 ;
        RECT 213.500 188.500 243.500 189.000 ;
        RECT 213.000 188.000 243.500 188.500 ;
        RECT 212.500 187.500 243.500 188.000 ;
        RECT 211.500 187.000 243.500 187.500 ;
        RECT 211.000 186.500 243.500 187.000 ;
        RECT 210.500 186.000 243.500 186.500 ;
        RECT 209.500 185.500 243.500 186.000 ;
        RECT 209.000 185.000 243.500 185.500 ;
        RECT 208.500 184.500 243.000 185.000 ;
        RECT 207.500 184.000 243.000 184.500 ;
        RECT 207.000 183.500 243.000 184.000 ;
        RECT 206.500 183.000 243.000 183.500 ;
        RECT 205.500 182.500 243.000 183.000 ;
        RECT 205.000 182.000 242.500 182.500 ;
        RECT 204.500 181.500 242.500 182.000 ;
        RECT 204.000 181.000 242.500 181.500 ;
        RECT 203.000 180.500 242.500 181.000 ;
        RECT 202.500 180.000 242.000 180.500 ;
        RECT 202.000 179.500 242.000 180.000 ;
        RECT 201.000 179.000 242.000 179.500 ;
        RECT 200.500 178.500 242.000 179.000 ;
        RECT 200.000 178.000 241.500 178.500 ;
        RECT 199.500 177.500 241.500 178.000 ;
        RECT 199.000 177.000 241.500 177.500 ;
        RECT 198.000 176.500 241.500 177.000 ;
        RECT 197.500 176.000 241.000 176.500 ;
        RECT 197.000 175.500 241.000 176.000 ;
        RECT 196.500 175.000 240.500 175.500 ;
        RECT 195.500 174.500 240.500 175.000 ;
        RECT 195.000 174.000 240.000 174.500 ;
        RECT 194.500 173.500 240.000 174.000 ;
        RECT 194.000 173.000 240.000 173.500 ;
        RECT 193.000 172.500 239.500 173.000 ;
        RECT 192.500 172.000 239.500 172.500 ;
        RECT 192.000 171.500 239.000 172.000 ;
        RECT 191.500 171.000 239.000 171.500 ;
        RECT 191.000 170.500 238.500 171.000 ;
        RECT 190.000 170.000 238.500 170.500 ;
        RECT 189.500 169.500 238.500 170.000 ;
        RECT 189.000 169.000 238.000 169.500 ;
        RECT 188.500 168.500 238.000 169.000 ;
        RECT 188.000 168.000 237.500 168.500 ;
        RECT 187.500 167.500 237.000 168.000 ;
        RECT 186.500 167.000 237.000 167.500 ;
        RECT 186.000 166.500 236.500 167.000 ;
        RECT 185.500 166.000 236.500 166.500 ;
        RECT 185.000 165.500 236.000 166.000 ;
        RECT 184.500 165.000 235.500 165.500 ;
        RECT 183.500 164.500 235.500 165.000 ;
        RECT 183.000 164.000 235.000 164.500 ;
        RECT 182.500 163.500 235.000 164.000 ;
        RECT 182.000 163.000 234.500 163.500 ;
        RECT 181.500 162.500 234.000 163.000 ;
        RECT 181.000 162.000 234.000 162.500 ;
        RECT 180.500 161.500 233.500 162.000 ;
        RECT 180.000 161.000 233.500 161.500 ;
        RECT 179.000 160.500 233.000 161.000 ;
        RECT 178.500 160.000 232.500 160.500 ;
        RECT 178.000 159.500 232.500 160.000 ;
        RECT 177.500 159.000 232.000 159.500 ;
        RECT 177.000 158.500 231.500 159.000 ;
        RECT 176.500 158.000 231.500 158.500 ;
        RECT 176.000 157.500 231.000 158.000 ;
        RECT 175.500 157.000 230.500 157.500 ;
        RECT 174.500 156.500 230.000 157.000 ;
        RECT 174.000 156.000 230.000 156.500 ;
        RECT 173.500 155.500 229.500 156.000 ;
        RECT 173.000 155.000 229.000 155.500 ;
        RECT 172.500 154.500 229.000 155.000 ;
        RECT 172.000 154.000 228.500 154.500 ;
        RECT 171.500 153.500 228.000 154.000 ;
        RECT 171.000 153.000 227.500 153.500 ;
        RECT 170.500 152.500 227.500 153.000 ;
        RECT 170.000 152.000 227.000 152.500 ;
        RECT 169.500 151.500 226.500 152.000 ;
        RECT 168.500 151.000 226.500 151.500 ;
        RECT 168.000 150.500 226.000 151.000 ;
        RECT 167.500 150.000 225.500 150.500 ;
        RECT 167.000 149.500 225.000 150.000 ;
        RECT 166.500 149.000 224.500 149.500 ;
        RECT 166.000 148.500 224.500 149.000 ;
        RECT 165.500 148.000 224.000 148.500 ;
        RECT 165.000 147.500 223.500 148.000 ;
        RECT 164.500 147.000 223.000 147.500 ;
        RECT 164.000 146.500 223.000 147.000 ;
        RECT 163.500 146.000 222.500 146.500 ;
        RECT 163.000 145.500 222.000 146.000 ;
        RECT 162.500 145.000 221.500 145.500 ;
        RECT 162.000 144.500 221.000 145.000 ;
        RECT 161.500 144.000 221.000 144.500 ;
        RECT 161.000 143.500 220.500 144.000 ;
        RECT 160.500 143.000 220.000 143.500 ;
        RECT 160.000 142.500 219.500 143.000 ;
        RECT 159.000 142.000 219.500 142.500 ;
        RECT 158.500 141.500 219.000 142.000 ;
        RECT 158.000 141.000 218.500 141.500 ;
        RECT 157.500 140.500 218.000 141.000 ;
        RECT 157.000 140.000 217.500 140.500 ;
        RECT 156.500 139.500 217.500 140.000 ;
        RECT 156.000 139.000 217.000 139.500 ;
        RECT 155.500 138.500 216.500 139.000 ;
        RECT 155.000 138.000 216.000 138.500 ;
        RECT 154.500 137.500 215.500 138.000 ;
        RECT 154.000 137.000 215.500 137.500 ;
        RECT 153.500 136.500 215.000 137.000 ;
        RECT 153.000 136.000 214.500 136.500 ;
        RECT 152.500 135.500 214.000 136.000 ;
        RECT 152.000 135.000 213.500 135.500 ;
        RECT 151.500 134.500 213.500 135.000 ;
        RECT 151.000 134.000 213.000 134.500 ;
        RECT 150.500 133.500 212.500 134.000 ;
        RECT 150.000 133.000 212.000 133.500 ;
        RECT 149.500 132.500 211.500 133.000 ;
        RECT 149.000 132.000 211.000 132.500 ;
        RECT 148.500 131.500 211.000 132.000 ;
        RECT 148.000 131.000 210.500 131.500 ;
        RECT 147.500 130.500 210.000 131.000 ;
        RECT 147.000 130.000 209.500 130.500 ;
        RECT 146.500 129.500 209.000 130.000 ;
        RECT 146.000 129.000 209.000 129.500 ;
        RECT 145.500 128.500 208.500 129.000 ;
        RECT 145.000 128.000 208.000 128.500 ;
        RECT 144.500 127.500 207.500 128.000 ;
        RECT 144.500 127.000 207.000 127.500 ;
        RECT 144.000 126.500 207.000 127.000 ;
        RECT 143.500 126.000 206.500 126.500 ;
        RECT 143.000 125.500 206.000 126.000 ;
        RECT 142.500 125.000 205.500 125.500 ;
        RECT 142.000 124.500 205.000 125.000 ;
        RECT 141.500 124.000 205.000 124.500 ;
        RECT 141.000 123.500 204.500 124.000 ;
        RECT 140.500 123.000 204.000 123.500 ;
        RECT 140.000 122.500 203.500 123.000 ;
        RECT 139.500 122.000 203.000 122.500 ;
        RECT 139.000 121.500 202.500 122.000 ;
        RECT 138.500 121.000 202.500 121.500 ;
        RECT 138.000 120.500 202.000 121.000 ;
        RECT 137.500 120.000 201.500 120.500 ;
        RECT 137.500 119.500 201.000 120.000 ;
        RECT 137.000 119.000 200.500 119.500 ;
        RECT 136.500 118.500 200.500 119.000 ;
        RECT 136.000 118.000 200.000 118.500 ;
        RECT 135.500 117.500 199.500 118.000 ;
        RECT 135.000 117.000 199.000 117.500 ;
        RECT 134.500 116.500 198.500 117.000 ;
        RECT 134.000 116.000 198.500 116.500 ;
        RECT 133.500 115.500 198.000 116.000 ;
        RECT 133.500 115.000 197.500 115.500 ;
        RECT 133.000 114.500 197.000 115.000 ;
        RECT 132.500 114.000 196.500 114.500 ;
        RECT 132.000 113.500 196.000 114.000 ;
        RECT 131.500 113.000 196.000 113.500 ;
        RECT 201.000 113.000 201.500 113.500 ;
        RECT 131.000 112.500 195.500 113.000 ;
        RECT 200.500 112.500 201.500 113.000 ;
        RECT 131.000 112.000 195.000 112.500 ;
        RECT 200.000 112.000 202.000 112.500 ;
        RECT 130.500 111.500 194.500 112.000 ;
        RECT 199.500 111.500 202.000 112.000 ;
        RECT 130.000 111.000 194.000 111.500 ;
        RECT 199.000 111.000 202.000 111.500 ;
        RECT 129.500 110.500 194.000 111.000 ;
        RECT 129.000 110.000 193.500 110.500 ;
        RECT 198.500 110.000 202.000 111.000 ;
        RECT 128.500 109.500 193.000 110.000 ;
        RECT 198.000 109.500 202.000 110.000 ;
        RECT 128.500 109.000 192.500 109.500 ;
        RECT 197.500 109.000 202.500 109.500 ;
        RECT 128.000 108.500 192.000 109.000 ;
        RECT 197.000 108.500 202.500 109.000 ;
        RECT 127.500 108.000 191.500 108.500 ;
        RECT 196.500 108.000 202.500 108.500 ;
        RECT 127.000 107.500 191.500 108.000 ;
        RECT 196.000 107.500 202.500 108.000 ;
        RECT 126.500 107.000 191.000 107.500 ;
        RECT 126.500 106.500 190.500 107.000 ;
        RECT 195.500 106.500 202.500 107.500 ;
        RECT 126.000 106.000 190.000 106.500 ;
        RECT 195.000 106.000 202.500 106.500 ;
        RECT 125.500 105.500 189.500 106.000 ;
        RECT 194.500 105.500 202.500 106.000 ;
        RECT 125.000 105.000 189.500 105.500 ;
        RECT 194.000 105.000 202.500 105.500 ;
        RECT 125.000 104.500 189.000 105.000 ;
        RECT 193.500 104.500 202.500 105.000 ;
        RECT 124.500 104.000 188.500 104.500 ;
        RECT 193.000 104.000 202.500 104.500 ;
        RECT 124.000 103.500 188.000 104.000 ;
        RECT 192.500 103.500 202.500 104.000 ;
        RECT 123.500 103.000 187.500 103.500 ;
        RECT 123.000 102.500 187.500 103.000 ;
        RECT 192.000 102.500 202.500 103.500 ;
        RECT 123.000 102.000 187.000 102.500 ;
        RECT 191.500 102.000 202.500 102.500 ;
        RECT 122.500 101.500 186.500 102.000 ;
        RECT 191.000 101.500 202.500 102.000 ;
        RECT 122.000 101.000 186.000 101.500 ;
        RECT 190.500 101.000 202.500 101.500 ;
        RECT 121.500 100.500 185.500 101.000 ;
        RECT 190.000 100.500 202.500 101.000 ;
        RECT 121.500 100.000 185.000 100.500 ;
        RECT 189.500 100.000 202.500 100.500 ;
        RECT 121.000 99.500 185.000 100.000 ;
        RECT 189.000 99.500 202.500 100.000 ;
        RECT 248.000 99.500 250.000 100.000 ;
        RECT 120.500 99.000 184.500 99.500 ;
        RECT 120.500 98.500 184.000 99.000 ;
        RECT 188.500 98.500 202.500 99.500 ;
        RECT 246.000 99.000 249.500 99.500 ;
        RECT 244.000 98.500 249.500 99.000 ;
        RECT 120.000 98.000 183.500 98.500 ;
        RECT 188.000 98.000 202.500 98.500 ;
        RECT 242.000 98.000 249.000 98.500 ;
        RECT 119.500 97.500 183.000 98.000 ;
        RECT 187.500 97.500 202.500 98.000 ;
        RECT 239.500 97.500 249.000 98.000 ;
        RECT 119.000 97.000 183.000 97.500 ;
        RECT 187.000 97.000 202.500 97.500 ;
        RECT 237.500 97.000 249.000 97.500 ;
        RECT 119.000 96.500 182.500 97.000 ;
        RECT 186.500 96.500 202.500 97.000 ;
        RECT 235.500 96.500 248.500 97.000 ;
        RECT 118.500 96.000 182.000 96.500 ;
        RECT 186.000 96.000 202.500 96.500 ;
        RECT 233.500 96.000 248.500 96.500 ;
        RECT 118.000 95.500 181.500 96.000 ;
        RECT 185.500 95.500 202.500 96.000 ;
        RECT 231.500 95.500 248.000 96.000 ;
        RECT 117.500 95.000 181.000 95.500 ;
        RECT 185.500 95.000 202.000 95.500 ;
        RECT 229.500 95.000 248.000 95.500 ;
        RECT 117.500 94.500 180.500 95.000 ;
        RECT 185.000 94.500 202.000 95.000 ;
        RECT 227.500 94.500 248.000 95.000 ;
        RECT 117.000 94.000 180.500 94.500 ;
        RECT 184.500 94.000 202.000 94.500 ;
        RECT 225.500 94.000 247.500 94.500 ;
        RECT 116.500 93.500 180.000 94.000 ;
        RECT 184.000 93.500 202.000 94.000 ;
        RECT 223.500 93.500 247.500 94.000 ;
        RECT 116.500 93.000 179.500 93.500 ;
        RECT 184.000 93.000 201.000 93.500 ;
        RECT 221.500 93.000 247.000 93.500 ;
        RECT 116.000 92.500 179.000 93.000 ;
        RECT 184.000 92.500 199.500 93.000 ;
        RECT 219.500 92.500 247.000 93.000 ;
        RECT 115.500 91.500 178.500 92.500 ;
        RECT 184.000 92.000 198.500 92.500 ;
        RECT 217.500 92.000 246.500 92.500 ;
        RECT 184.000 91.500 197.000 92.000 ;
        RECT 216.000 91.500 246.500 92.000 ;
        RECT 115.000 91.000 178.000 91.500 ;
        RECT 184.000 91.000 195.500 91.500 ;
        RECT 214.000 91.000 246.000 91.500 ;
        RECT 114.500 90.500 177.500 91.000 ;
        RECT 184.000 90.500 194.500 91.000 ;
        RECT 212.000 90.500 246.000 91.000 ;
        RECT 114.000 90.000 177.000 90.500 ;
        RECT 184.000 90.000 193.000 90.500 ;
        RECT 210.000 90.000 245.500 90.500 ;
        RECT 114.000 89.500 176.500 90.000 ;
        RECT 184.000 89.500 191.500 90.000 ;
        RECT 208.500 89.500 245.500 90.000 ;
        RECT 113.500 89.000 176.000 89.500 ;
        RECT 113.000 88.500 176.000 89.000 ;
        RECT 184.000 89.000 190.000 89.500 ;
        RECT 206.500 89.000 245.000 89.500 ;
        RECT 184.000 88.500 189.000 89.000 ;
        RECT 204.500 88.500 245.000 89.000 ;
        RECT 113.000 88.000 175.500 88.500 ;
        RECT 184.000 88.000 187.500 88.500 ;
        RECT 203.000 88.000 244.500 88.500 ;
        RECT 112.500 87.500 175.000 88.000 ;
        RECT 184.000 87.500 186.000 88.000 ;
        RECT 201.000 87.500 244.500 88.000 ;
        RECT 112.000 87.000 174.500 87.500 ;
        RECT 183.500 87.000 184.500 87.500 ;
        RECT 199.500 87.000 244.000 87.500 ;
        RECT 112.000 86.500 174.000 87.000 ;
        RECT 197.500 86.500 243.500 87.000 ;
        RECT 111.500 86.000 173.500 86.500 ;
        RECT 196.000 86.000 243.500 86.500 ;
        RECT 111.000 85.500 172.500 86.000 ;
        RECT 194.000 85.500 243.000 86.000 ;
        RECT 111.000 85.000 171.500 85.500 ;
        RECT 192.500 85.000 243.000 85.500 ;
        RECT 110.500 84.500 170.500 85.000 ;
        RECT 190.500 84.500 242.500 85.000 ;
        RECT 110.000 84.000 169.500 84.500 ;
        RECT 189.000 84.000 242.000 84.500 ;
        RECT 110.000 83.500 168.500 84.000 ;
        RECT 187.500 83.500 241.500 84.000 ;
        RECT 109.500 83.000 167.500 83.500 ;
        RECT 186.000 83.000 241.000 83.500 ;
        RECT 109.000 82.500 166.500 83.000 ;
        RECT 184.500 82.500 241.000 83.000 ;
        RECT 109.000 82.000 165.500 82.500 ;
        RECT 183.000 82.000 240.500 82.500 ;
        RECT 108.500 81.500 164.500 82.000 ;
        RECT 181.500 81.500 240.000 82.000 ;
        RECT 108.000 81.000 163.500 81.500 ;
        RECT 180.000 81.000 239.500 81.500 ;
        RECT 108.000 80.500 162.500 81.000 ;
        RECT 178.500 80.500 239.000 81.000 ;
        RECT 107.500 80.000 161.500 80.500 ;
        RECT 177.000 80.000 238.500 80.500 ;
        RECT 107.000 79.500 160.500 80.000 ;
        RECT 175.500 79.500 238.500 80.000 ;
        RECT 107.000 79.000 160.000 79.500 ;
        RECT 174.500 79.000 238.000 79.500 ;
        RECT 106.500 78.500 159.000 79.000 ;
        RECT 173.000 78.500 237.500 79.000 ;
        RECT 106.000 78.000 158.000 78.500 ;
        RECT 171.500 78.000 237.000 78.500 ;
        RECT 106.000 77.500 157.000 78.000 ;
        RECT 170.500 77.500 236.500 78.000 ;
        RECT 105.500 77.000 156.000 77.500 ;
        RECT 169.000 77.000 236.000 77.500 ;
        RECT 105.000 76.500 155.000 77.000 ;
        RECT 168.000 76.500 235.500 77.000 ;
        RECT 105.000 76.000 154.000 76.500 ;
        RECT 166.500 76.000 235.000 76.500 ;
        RECT 104.500 75.500 153.000 76.000 ;
        RECT 165.500 75.500 234.000 76.000 ;
        RECT 104.000 75.000 152.500 75.500 ;
        RECT 164.000 75.000 233.500 75.500 ;
        RECT 104.000 74.500 151.500 75.000 ;
        RECT 163.000 74.500 233.000 75.000 ;
        RECT 103.500 74.000 150.500 74.500 ;
        RECT 162.000 74.000 232.500 74.500 ;
        RECT 103.000 73.500 149.500 74.000 ;
        RECT 161.000 73.500 232.000 74.000 ;
        RECT 103.000 73.000 148.500 73.500 ;
        RECT 160.000 73.000 231.000 73.500 ;
        RECT 102.500 72.500 147.500 73.000 ;
        RECT 158.500 72.500 230.500 73.000 ;
        RECT 102.000 72.000 147.000 72.500 ;
        RECT 157.500 72.000 230.000 72.500 ;
        RECT 102.000 71.500 146.000 72.000 ;
        RECT 156.500 71.500 229.500 72.000 ;
        RECT 101.500 71.000 145.000 71.500 ;
        RECT 155.500 71.000 228.500 71.500 ;
        RECT 101.500 70.500 144.000 71.000 ;
        RECT 154.500 70.500 228.000 71.000 ;
        RECT 101.000 70.000 143.000 70.500 ;
        RECT 153.500 70.000 227.500 70.500 ;
        RECT 100.500 69.500 142.500 70.000 ;
        RECT 152.500 69.500 226.500 70.000 ;
        RECT 100.500 69.000 141.500 69.500 ;
        RECT 151.500 69.000 226.000 69.500 ;
        RECT 100.000 68.500 140.500 69.000 ;
        RECT 150.500 68.500 225.000 69.000 ;
        RECT 99.500 68.000 139.500 68.500 ;
        RECT 150.000 68.000 224.500 68.500 ;
        RECT 99.500 67.500 139.000 68.000 ;
        RECT 149.000 67.500 224.000 68.000 ;
        RECT 99.000 67.000 138.000 67.500 ;
        RECT 148.000 67.000 223.000 67.500 ;
        RECT 98.500 66.500 137.000 67.000 ;
        RECT 147.000 66.500 222.500 67.000 ;
        RECT 98.500 66.000 136.500 66.500 ;
        RECT 146.500 66.000 221.500 66.500 ;
        RECT 98.000 65.500 135.500 66.000 ;
        RECT 145.500 65.500 221.000 66.000 ;
        RECT 98.000 65.000 134.500 65.500 ;
        RECT 144.500 65.000 220.000 65.500 ;
        RECT 97.500 64.500 134.000 65.000 ;
        RECT 143.500 64.500 219.500 65.000 ;
        RECT 97.000 64.000 133.000 64.500 ;
        RECT 143.000 64.000 218.500 64.500 ;
        RECT 97.000 63.500 132.000 64.000 ;
        RECT 142.000 63.500 217.500 64.000 ;
        RECT 96.500 63.000 131.500 63.500 ;
        RECT 141.500 63.000 217.000 63.500 ;
        RECT 96.000 62.500 130.500 63.000 ;
        RECT 140.500 62.500 216.000 63.000 ;
        RECT 96.000 62.000 130.000 62.500 ;
        RECT 139.500 62.000 215.500 62.500 ;
        RECT 95.500 61.500 129.000 62.000 ;
        RECT 139.000 61.500 214.500 62.000 ;
        RECT 95.500 61.000 128.000 61.500 ;
        RECT 138.000 61.000 214.000 61.500 ;
        RECT 95.000 60.500 127.500 61.000 ;
        RECT 137.500 60.500 213.000 61.000 ;
        RECT 94.500 60.000 126.500 60.500 ;
        RECT 136.500 60.000 212.500 60.500 ;
        RECT 94.500 59.500 126.000 60.000 ;
        RECT 135.500 59.500 211.500 60.000 ;
        RECT 94.000 59.000 125.000 59.500 ;
        RECT 135.000 59.000 210.500 59.500 ;
        RECT 94.000 58.500 124.000 59.000 ;
        RECT 134.000 58.500 210.000 59.000 ;
        RECT 93.500 58.000 123.500 58.500 ;
        RECT 133.500 58.000 209.000 58.500 ;
        RECT 93.000 57.500 122.500 58.000 ;
        RECT 132.500 57.500 208.000 58.000 ;
        RECT 93.000 57.000 122.000 57.500 ;
        RECT 132.000 57.000 207.500 57.500 ;
        RECT 92.500 56.500 121.000 57.000 ;
        RECT 131.000 56.500 206.500 57.000 ;
        RECT 92.000 56.000 120.500 56.500 ;
        RECT 130.500 56.000 205.500 56.500 ;
        RECT 92.000 55.500 119.500 56.000 ;
        RECT 129.500 55.500 205.000 56.000 ;
        RECT 91.500 55.000 119.000 55.500 ;
        RECT 129.000 55.000 204.000 55.500 ;
        RECT 91.500 54.500 118.000 55.000 ;
        RECT 128.000 54.500 203.000 55.000 ;
        RECT 91.000 54.000 117.500 54.500 ;
        RECT 127.500 54.000 202.500 54.500 ;
        RECT 90.500 53.500 116.500 54.000 ;
        RECT 126.500 53.500 201.500 54.000 ;
        RECT 90.500 53.000 116.000 53.500 ;
        RECT 126.000 53.000 200.500 53.500 ;
        RECT 90.000 52.500 115.000 53.000 ;
        RECT 125.000 52.500 200.000 53.000 ;
        RECT 90.000 52.000 114.500 52.500 ;
        RECT 124.500 52.000 199.000 52.500 ;
        RECT 89.500 51.500 114.000 52.000 ;
        RECT 123.500 51.500 198.000 52.000 ;
        RECT 89.500 51.000 113.000 51.500 ;
        RECT 123.000 51.000 197.500 51.500 ;
        RECT 89.000 50.500 112.500 51.000 ;
        RECT 122.000 50.500 196.500 51.000 ;
        RECT 88.500 50.000 111.500 50.500 ;
        RECT 121.500 50.000 195.500 50.500 ;
        RECT 88.500 49.500 111.000 50.000 ;
        RECT 120.500 49.500 195.000 50.000 ;
        RECT 88.000 49.000 110.000 49.500 ;
        RECT 120.000 49.000 194.000 49.500 ;
        RECT 88.000 48.500 109.500 49.000 ;
        RECT 119.000 48.500 193.000 49.000 ;
        RECT 87.500 48.000 109.000 48.500 ;
        RECT 118.500 48.000 192.500 48.500 ;
        RECT 87.000 47.500 108.000 48.000 ;
        RECT 117.500 47.500 191.500 48.000 ;
        RECT 87.000 47.000 107.500 47.500 ;
        RECT 117.000 47.000 190.500 47.500 ;
        RECT 86.500 46.500 106.500 47.000 ;
        RECT 116.000 46.500 190.000 47.000 ;
        RECT 86.500 46.000 106.000 46.500 ;
        RECT 115.500 46.000 189.000 46.500 ;
        RECT 86.000 45.500 105.500 46.000 ;
        RECT 114.500 45.500 188.000 46.000 ;
        RECT 86.000 45.000 104.500 45.500 ;
        RECT 114.000 45.000 187.500 45.500 ;
        RECT 85.500 44.500 104.000 45.000 ;
        RECT 113.000 44.500 186.500 45.000 ;
        RECT 85.500 44.000 103.500 44.500 ;
        RECT 112.500 44.000 185.500 44.500 ;
        RECT 85.000 43.500 102.500 44.000 ;
        RECT 111.500 43.500 185.000 44.000 ;
        RECT 85.000 43.000 102.000 43.500 ;
        RECT 111.000 43.000 184.000 43.500 ;
        RECT 84.500 42.500 101.500 43.000 ;
        RECT 110.000 42.500 183.000 43.000 ;
        RECT 84.000 42.000 100.500 42.500 ;
        RECT 109.500 42.000 182.500 42.500 ;
        RECT 84.000 41.500 100.000 42.000 ;
        RECT 108.500 41.500 181.500 42.000 ;
        RECT 83.500 41.000 99.500 41.500 ;
        RECT 108.000 41.000 180.500 41.500 ;
        RECT 83.500 40.500 99.000 41.000 ;
        RECT 107.000 40.500 180.000 41.000 ;
        RECT 83.000 40.000 98.000 40.500 ;
        RECT 106.500 40.000 179.000 40.500 ;
        RECT 83.000 39.500 97.500 40.000 ;
        RECT 105.500 39.500 178.500 40.000 ;
        RECT 82.500 39.000 97.000 39.500 ;
        RECT 105.000 39.000 177.500 39.500 ;
        RECT 82.500 38.500 96.000 39.000 ;
        RECT 104.500 38.500 176.500 39.000 ;
        RECT 82.000 38.000 95.500 38.500 ;
        RECT 103.500 38.000 175.500 38.500 ;
        RECT 82.000 37.500 95.000 38.000 ;
        RECT 103.000 37.500 174.500 38.000 ;
        RECT 81.500 37.000 94.500 37.500 ;
        RECT 102.000 37.000 173.000 37.500 ;
        RECT 81.500 36.500 93.500 37.000 ;
        RECT 101.500 36.500 172.000 37.000 ;
        RECT 81.000 36.000 93.000 36.500 ;
        RECT 100.500 36.000 170.500 36.500 ;
        RECT 81.000 35.500 92.500 36.000 ;
        RECT 100.000 35.500 169.500 36.000 ;
        RECT 81.000 35.000 92.000 35.500 ;
        RECT 99.500 35.000 168.000 35.500 ;
        RECT 80.500 34.500 91.000 35.000 ;
        RECT 98.500 34.500 166.500 35.000 ;
        RECT 80.500 34.000 90.500 34.500 ;
        RECT 98.000 34.000 165.500 34.500 ;
        RECT 80.000 33.500 90.000 34.000 ;
        RECT 97.000 33.500 164.000 34.000 ;
        RECT 175.000 33.500 176.000 34.000 ;
        RECT 80.000 33.000 89.500 33.500 ;
        RECT 96.500 33.000 163.000 33.500 ;
        RECT 173.500 33.000 175.500 33.500 ;
        RECT 79.500 32.500 88.500 33.000 ;
        RECT 95.500 32.500 161.500 33.000 ;
        RECT 172.500 32.500 175.000 33.000 ;
        RECT 79.500 32.000 88.000 32.500 ;
        RECT 95.000 32.000 160.500 32.500 ;
        RECT 171.000 32.000 174.500 32.500 ;
        RECT 79.500 31.500 87.500 32.000 ;
        RECT 94.500 31.500 159.000 32.000 ;
        RECT 169.500 31.500 174.000 32.000 ;
        RECT 79.000 31.000 86.500 31.500 ;
        RECT 93.500 31.000 158.000 31.500 ;
        RECT 168.500 31.000 173.500 31.500 ;
        RECT 79.000 30.500 86.000 31.000 ;
        RECT 93.000 30.500 156.500 31.000 ;
        RECT 167.000 30.500 173.000 31.000 ;
        RECT 78.500 30.000 85.500 30.500 ;
        RECT 92.500 30.000 155.500 30.500 ;
        RECT 165.500 30.000 172.500 30.500 ;
        RECT 78.500 29.500 85.000 30.000 ;
        RECT 91.500 29.500 154.000 30.000 ;
        RECT 164.500 29.500 172.000 30.000 ;
        RECT 78.500 29.000 84.000 29.500 ;
        RECT 91.000 29.000 153.000 29.500 ;
        RECT 163.000 29.000 171.000 29.500 ;
        RECT 78.000 28.500 83.500 29.000 ;
        RECT 90.000 28.500 151.500 29.000 ;
        RECT 161.500 28.500 170.500 29.000 ;
        RECT 78.000 28.000 83.000 28.500 ;
        RECT 89.500 28.000 150.000 28.500 ;
        RECT 160.000 28.000 170.000 28.500 ;
        RECT 77.500 27.500 82.000 28.000 ;
        RECT 89.000 27.500 149.000 28.000 ;
        RECT 159.000 27.500 169.500 28.000 ;
        RECT 77.500 27.000 81.500 27.500 ;
        RECT 88.000 27.000 147.500 27.500 ;
        RECT 157.500 27.000 169.000 27.500 ;
        RECT 77.500 26.500 81.000 27.000 ;
        RECT 87.500 26.500 146.500 27.000 ;
        RECT 156.000 26.500 168.500 27.000 ;
        RECT 77.000 26.000 80.000 26.500 ;
        RECT 87.000 26.000 145.000 26.500 ;
        RECT 155.000 26.000 168.000 26.500 ;
        RECT 77.000 25.500 79.500 26.000 ;
        RECT 86.000 25.500 144.000 26.000 ;
        RECT 153.500 25.500 167.500 26.000 ;
        RECT 77.000 25.000 79.000 25.500 ;
        RECT 85.500 25.000 142.500 25.500 ;
        RECT 152.000 25.000 167.000 25.500 ;
        RECT 76.500 24.500 78.000 25.000 ;
        RECT 85.000 24.500 141.500 25.000 ;
        RECT 151.000 24.500 166.500 25.000 ;
        RECT 76.500 24.000 77.500 24.500 ;
        RECT 84.000 24.000 140.000 24.500 ;
        RECT 149.500 24.000 165.500 24.500 ;
        RECT 76.000 23.500 77.000 24.000 ;
        RECT 83.500 23.500 103.500 24.000 ;
        RECT 148.000 23.500 165.000 24.000 ;
        RECT 83.000 23.000 100.000 23.500 ;
        RECT 147.000 23.000 164.500 23.500 ;
        RECT 82.000 22.500 98.000 23.000 ;
        RECT 145.500 22.500 164.000 23.000 ;
        RECT 81.500 22.000 96.000 22.500 ;
        RECT 144.000 22.000 163.500 22.500 ;
        RECT 81.000 21.500 95.000 22.000 ;
        RECT 143.000 21.500 163.000 22.000 ;
        RECT 80.500 21.000 93.500 21.500 ;
        RECT 141.500 21.000 162.500 21.500 ;
        RECT 80.000 20.500 92.500 21.000 ;
        RECT 125.500 20.500 161.500 21.000 ;
        RECT 79.000 20.000 91.500 20.500 ;
        RECT 123.500 20.000 161.000 20.500 ;
        RECT 78.500 19.500 90.000 20.000 ;
        RECT 122.000 19.500 160.500 20.000 ;
        RECT 78.000 19.000 89.500 19.500 ;
        RECT 120.000 19.000 159.500 19.500 ;
        RECT 77.500 18.500 88.500 19.000 ;
        RECT 117.500 18.500 159.000 19.000 ;
        RECT 77.000 18.000 87.500 18.500 ;
        RECT 114.500 18.000 158.500 18.500 ;
        RECT 76.500 17.500 86.500 18.000 ;
        RECT 110.500 17.500 158.000 18.000 ;
        RECT 76.000 17.000 86.000 17.500 ;
        RECT 91.000 17.000 97.500 17.500 ;
        RECT 103.500 17.000 157.000 17.500 ;
        RECT 75.500 16.500 85.000 17.000 ;
        RECT 90.500 16.500 156.500 17.000 ;
        RECT 75.000 16.000 84.500 16.500 ;
        RECT 90.000 16.000 155.500 16.500 ;
        RECT 74.500 15.500 83.500 16.000 ;
        RECT 89.000 15.500 155.000 16.000 ;
        RECT 74.000 15.000 83.000 15.500 ;
        RECT 88.500 15.000 154.000 15.500 ;
        RECT 73.500 14.500 82.000 15.000 ;
        RECT 88.000 14.500 153.500 15.000 ;
        RECT 73.500 14.000 81.500 14.500 ;
        RECT 87.500 14.000 152.500 14.500 ;
        RECT 73.000 13.500 81.000 14.000 ;
        RECT 87.000 13.500 152.000 14.000 ;
        RECT 72.500 13.000 80.000 13.500 ;
        RECT 86.000 13.000 151.000 13.500 ;
        RECT 72.500 12.500 79.500 13.000 ;
        RECT 85.500 12.500 150.000 13.000 ;
        RECT 72.000 12.000 79.000 12.500 ;
        RECT 85.000 12.000 149.500 12.500 ;
        RECT 71.500 11.500 78.000 12.000 ;
        RECT 84.500 11.500 148.500 12.000 ;
        RECT 71.500 11.000 77.500 11.500 ;
        RECT 83.500 11.000 147.500 11.500 ;
        RECT 71.000 10.500 77.000 11.000 ;
        RECT 83.000 10.500 146.500 11.000 ;
        RECT 71.000 10.000 76.000 10.500 ;
        RECT 82.500 10.000 145.500 10.500 ;
        RECT 70.500 9.500 75.500 10.000 ;
        RECT 82.000 9.500 144.500 10.000 ;
        RECT 63.500 9.000 64.000 9.500 ;
        RECT 70.500 9.000 74.500 9.500 ;
        RECT 81.000 9.000 143.500 9.500 ;
        RECT 70.000 8.500 74.000 9.000 ;
        RECT 80.500 8.500 142.500 9.000 ;
        RECT 70.000 8.000 73.000 8.500 ;
        RECT 80.000 8.000 141.500 8.500 ;
        RECT 69.500 7.500 72.500 8.000 ;
        RECT 79.500 7.500 140.000 8.000 ;
        RECT 69.500 7.000 71.500 7.500 ;
        RECT 79.000 7.000 139.000 7.500 ;
        RECT 69.000 6.500 70.500 7.000 ;
        RECT 78.000 6.500 137.500 7.000 ;
        RECT 69.000 6.000 70.000 6.500 ;
        RECT 77.500 6.000 136.500 6.500 ;
        RECT 68.500 5.500 69.000 6.000 ;
        RECT 77.000 5.500 135.000 6.000 ;
        RECT 76.500 5.000 133.500 5.500 ;
        RECT 75.500 4.500 132.000 5.000 ;
        RECT 75.000 4.000 130.500 4.500 ;
        RECT 74.500 3.500 128.500 4.000 ;
        RECT 76.500 3.000 127.000 3.500 ;
        RECT 79.500 2.500 125.000 3.000 ;
        RECT 83.000 2.000 122.500 2.500 ;
        RECT 86.000 1.500 120.500 2.000 ;
        RECT 90.000 1.000 117.500 1.500 ;
        RECT 94.000 0.500 114.000 1.000 ;
        RECT 101.000 0.000 107.000 0.500 ;
  END
END avali_logo
END LIBRARY

