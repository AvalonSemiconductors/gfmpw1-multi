magic
tech gf180mcuD
magscale 1 5
timestamp 1698973806
<< obsm1 >>
rect 672 1538 49280 48313
<< metal2 >>
rect 3136 49600 3192 50000
rect 3808 49600 3864 50000
rect 4480 49600 4536 50000
rect 5152 49600 5208 50000
rect 5824 49600 5880 50000
rect 6496 49600 6552 50000
rect 7168 49600 7224 50000
rect 7840 49600 7896 50000
rect 8512 49600 8568 50000
rect 9184 49600 9240 50000
rect 9856 49600 9912 50000
rect 10528 49600 10584 50000
rect 11200 49600 11256 50000
rect 11872 49600 11928 50000
rect 12544 49600 12600 50000
rect 13216 49600 13272 50000
rect 13888 49600 13944 50000
rect 14560 49600 14616 50000
rect 15232 49600 15288 50000
rect 15904 49600 15960 50000
rect 16576 49600 16632 50000
rect 17248 49600 17304 50000
rect 17920 49600 17976 50000
rect 18592 49600 18648 50000
rect 19264 49600 19320 50000
rect 19936 49600 19992 50000
rect 20608 49600 20664 50000
rect 21280 49600 21336 50000
rect 21952 49600 22008 50000
rect 22624 49600 22680 50000
rect 23296 49600 23352 50000
rect 23968 49600 24024 50000
rect 24640 49600 24696 50000
rect 25312 49600 25368 50000
rect 25984 49600 26040 50000
rect 26656 49600 26712 50000
rect 27328 49600 27384 50000
rect 28000 49600 28056 50000
rect 28672 49600 28728 50000
rect 29344 49600 29400 50000
rect 30016 49600 30072 50000
rect 30688 49600 30744 50000
rect 31360 49600 31416 50000
rect 32032 49600 32088 50000
rect 32704 49600 32760 50000
rect 33376 49600 33432 50000
rect 34048 49600 34104 50000
rect 34720 49600 34776 50000
rect 35392 49600 35448 50000
rect 36064 49600 36120 50000
rect 36736 49600 36792 50000
rect 37408 49600 37464 50000
rect 38080 49600 38136 50000
rect 38752 49600 38808 50000
rect 39424 49600 39480 50000
rect 40096 49600 40152 50000
rect 40768 49600 40824 50000
rect 41440 49600 41496 50000
rect 42112 49600 42168 50000
rect 42784 49600 42840 50000
rect 43456 49600 43512 50000
rect 44128 49600 44184 50000
rect 44800 49600 44856 50000
rect 45472 49600 45528 50000
rect 46144 49600 46200 50000
rect 46816 49600 46872 50000
<< obsm2 >>
rect 14 49570 3106 49658
rect 3222 49570 3778 49658
rect 3894 49570 4450 49658
rect 4566 49570 5122 49658
rect 5238 49570 5794 49658
rect 5910 49570 6466 49658
rect 6582 49570 7138 49658
rect 7254 49570 7810 49658
rect 7926 49570 8482 49658
rect 8598 49570 9154 49658
rect 9270 49570 9826 49658
rect 9942 49570 10498 49658
rect 10614 49570 11170 49658
rect 11286 49570 11842 49658
rect 11958 49570 12514 49658
rect 12630 49570 13186 49658
rect 13302 49570 13858 49658
rect 13974 49570 14530 49658
rect 14646 49570 15202 49658
rect 15318 49570 15874 49658
rect 15990 49570 16546 49658
rect 16662 49570 17218 49658
rect 17334 49570 17890 49658
rect 18006 49570 18562 49658
rect 18678 49570 19234 49658
rect 19350 49570 19906 49658
rect 20022 49570 20578 49658
rect 20694 49570 21250 49658
rect 21366 49570 21922 49658
rect 22038 49570 22594 49658
rect 22710 49570 23266 49658
rect 23382 49570 23938 49658
rect 24054 49570 24610 49658
rect 24726 49570 25282 49658
rect 25398 49570 25954 49658
rect 26070 49570 26626 49658
rect 26742 49570 27298 49658
rect 27414 49570 27970 49658
rect 28086 49570 28642 49658
rect 28758 49570 29314 49658
rect 29430 49570 29986 49658
rect 30102 49570 30658 49658
rect 30774 49570 31330 49658
rect 31446 49570 32002 49658
rect 32118 49570 32674 49658
rect 32790 49570 33346 49658
rect 33462 49570 34018 49658
rect 34134 49570 34690 49658
rect 34806 49570 35362 49658
rect 35478 49570 36034 49658
rect 36150 49570 36706 49658
rect 36822 49570 37378 49658
rect 37494 49570 38050 49658
rect 38166 49570 38722 49658
rect 38838 49570 39394 49658
rect 39510 49570 40066 49658
rect 40182 49570 40738 49658
rect 40854 49570 41410 49658
rect 41526 49570 42082 49658
rect 42198 49570 42754 49658
rect 42870 49570 43426 49658
rect 43542 49570 44098 49658
rect 44214 49570 44770 49658
rect 44886 49570 45442 49658
rect 45558 49570 46114 49658
rect 46230 49570 46786 49658
rect 46902 49570 49378 49658
rect 14 569 49378 49570
<< metal3 >>
rect 0 48944 400 49000
rect 0 47488 400 47544
rect 49600 46480 50000 46536
rect 0 46032 400 46088
rect 49600 45696 50000 45752
rect 49600 44912 50000 44968
rect 0 44576 400 44632
rect 49600 44128 50000 44184
rect 49600 43344 50000 43400
rect 0 43120 400 43176
rect 49600 42560 50000 42616
rect 49600 41776 50000 41832
rect 0 41664 400 41720
rect 49600 40992 50000 41048
rect 0 40208 400 40264
rect 49600 40208 50000 40264
rect 49600 39424 50000 39480
rect 0 38752 400 38808
rect 49600 38640 50000 38696
rect 49600 37856 50000 37912
rect 0 37296 400 37352
rect 49600 37072 50000 37128
rect 49600 36288 50000 36344
rect 0 35840 400 35896
rect 49600 35504 50000 35560
rect 49600 34720 50000 34776
rect 0 34384 400 34440
rect 49600 33936 50000 33992
rect 49600 33152 50000 33208
rect 0 32928 400 32984
rect 49600 32368 50000 32424
rect 49600 31584 50000 31640
rect 0 31472 400 31528
rect 49600 30800 50000 30856
rect 0 30016 400 30072
rect 49600 30016 50000 30072
rect 49600 29232 50000 29288
rect 0 28560 400 28616
rect 49600 28448 50000 28504
rect 49600 27664 50000 27720
rect 0 27104 400 27160
rect 49600 26880 50000 26936
rect 49600 26096 50000 26152
rect 0 25648 400 25704
rect 49600 25312 50000 25368
rect 49600 24528 50000 24584
rect 0 24192 400 24248
rect 49600 23744 50000 23800
rect 49600 22960 50000 23016
rect 0 22736 400 22792
rect 49600 22176 50000 22232
rect 49600 21392 50000 21448
rect 0 21280 400 21336
rect 49600 20608 50000 20664
rect 0 19824 400 19880
rect 49600 19824 50000 19880
rect 49600 19040 50000 19096
rect 0 18368 400 18424
rect 49600 18256 50000 18312
rect 49600 17472 50000 17528
rect 0 16912 400 16968
rect 49600 16688 50000 16744
rect 49600 15904 50000 15960
rect 0 15456 400 15512
rect 49600 15120 50000 15176
rect 49600 14336 50000 14392
rect 0 14000 400 14056
rect 49600 13552 50000 13608
rect 49600 12768 50000 12824
rect 0 12544 400 12600
rect 49600 11984 50000 12040
rect 49600 11200 50000 11256
rect 0 11088 400 11144
rect 49600 10416 50000 10472
rect 0 9632 400 9688
rect 49600 9632 50000 9688
rect 49600 8848 50000 8904
rect 0 8176 400 8232
rect 49600 8064 50000 8120
rect 49600 7280 50000 7336
rect 0 6720 400 6776
rect 49600 6496 50000 6552
rect 49600 5712 50000 5768
rect 0 5264 400 5320
rect 49600 4928 50000 4984
rect 49600 4144 50000 4200
rect 0 3808 400 3864
rect 49600 3360 50000 3416
rect 0 2352 400 2408
rect 0 896 400 952
<< obsm3 >>
rect 430 48914 49658 48986
rect 9 47574 49658 48914
rect 430 47458 49658 47574
rect 9 46566 49658 47458
rect 9 46450 49570 46566
rect 9 46118 49658 46450
rect 430 46002 49658 46118
rect 9 45782 49658 46002
rect 9 45666 49570 45782
rect 9 44998 49658 45666
rect 9 44882 49570 44998
rect 9 44662 49658 44882
rect 430 44546 49658 44662
rect 9 44214 49658 44546
rect 9 44098 49570 44214
rect 9 43430 49658 44098
rect 9 43314 49570 43430
rect 9 43206 49658 43314
rect 430 43090 49658 43206
rect 9 42646 49658 43090
rect 9 42530 49570 42646
rect 9 41862 49658 42530
rect 9 41750 49570 41862
rect 430 41746 49570 41750
rect 430 41634 49658 41746
rect 9 41078 49658 41634
rect 9 40962 49570 41078
rect 9 40294 49658 40962
rect 430 40178 49570 40294
rect 9 39510 49658 40178
rect 9 39394 49570 39510
rect 9 38838 49658 39394
rect 430 38726 49658 38838
rect 430 38722 49570 38726
rect 9 38610 49570 38722
rect 9 37942 49658 38610
rect 9 37826 49570 37942
rect 9 37382 49658 37826
rect 430 37266 49658 37382
rect 9 37158 49658 37266
rect 9 37042 49570 37158
rect 9 36374 49658 37042
rect 9 36258 49570 36374
rect 9 35926 49658 36258
rect 430 35810 49658 35926
rect 9 35590 49658 35810
rect 9 35474 49570 35590
rect 9 34806 49658 35474
rect 9 34690 49570 34806
rect 9 34470 49658 34690
rect 430 34354 49658 34470
rect 9 34022 49658 34354
rect 9 33906 49570 34022
rect 9 33238 49658 33906
rect 9 33122 49570 33238
rect 9 33014 49658 33122
rect 430 32898 49658 33014
rect 9 32454 49658 32898
rect 9 32338 49570 32454
rect 9 31670 49658 32338
rect 9 31558 49570 31670
rect 430 31554 49570 31558
rect 430 31442 49658 31554
rect 9 30886 49658 31442
rect 9 30770 49570 30886
rect 9 30102 49658 30770
rect 430 29986 49570 30102
rect 9 29318 49658 29986
rect 9 29202 49570 29318
rect 9 28646 49658 29202
rect 430 28534 49658 28646
rect 430 28530 49570 28534
rect 9 28418 49570 28530
rect 9 27750 49658 28418
rect 9 27634 49570 27750
rect 9 27190 49658 27634
rect 430 27074 49658 27190
rect 9 26966 49658 27074
rect 9 26850 49570 26966
rect 9 26182 49658 26850
rect 9 26066 49570 26182
rect 9 25734 49658 26066
rect 430 25618 49658 25734
rect 9 25398 49658 25618
rect 9 25282 49570 25398
rect 9 24614 49658 25282
rect 9 24498 49570 24614
rect 9 24278 49658 24498
rect 430 24162 49658 24278
rect 9 23830 49658 24162
rect 9 23714 49570 23830
rect 9 23046 49658 23714
rect 9 22930 49570 23046
rect 9 22822 49658 22930
rect 430 22706 49658 22822
rect 9 22262 49658 22706
rect 9 22146 49570 22262
rect 9 21478 49658 22146
rect 9 21366 49570 21478
rect 430 21362 49570 21366
rect 430 21250 49658 21362
rect 9 20694 49658 21250
rect 9 20578 49570 20694
rect 9 19910 49658 20578
rect 430 19794 49570 19910
rect 9 19126 49658 19794
rect 9 19010 49570 19126
rect 9 18454 49658 19010
rect 430 18342 49658 18454
rect 430 18338 49570 18342
rect 9 18226 49570 18338
rect 9 17558 49658 18226
rect 9 17442 49570 17558
rect 9 16998 49658 17442
rect 430 16882 49658 16998
rect 9 16774 49658 16882
rect 9 16658 49570 16774
rect 9 15990 49658 16658
rect 9 15874 49570 15990
rect 9 15542 49658 15874
rect 430 15426 49658 15542
rect 9 15206 49658 15426
rect 9 15090 49570 15206
rect 9 14422 49658 15090
rect 9 14306 49570 14422
rect 9 14086 49658 14306
rect 430 13970 49658 14086
rect 9 13638 49658 13970
rect 9 13522 49570 13638
rect 9 12854 49658 13522
rect 9 12738 49570 12854
rect 9 12630 49658 12738
rect 430 12514 49658 12630
rect 9 12070 49658 12514
rect 9 11954 49570 12070
rect 9 11286 49658 11954
rect 9 11174 49570 11286
rect 430 11170 49570 11174
rect 430 11058 49658 11170
rect 9 10502 49658 11058
rect 9 10386 49570 10502
rect 9 9718 49658 10386
rect 430 9602 49570 9718
rect 9 8934 49658 9602
rect 9 8818 49570 8934
rect 9 8262 49658 8818
rect 430 8150 49658 8262
rect 430 8146 49570 8150
rect 9 8034 49570 8146
rect 9 7366 49658 8034
rect 9 7250 49570 7366
rect 9 6806 49658 7250
rect 430 6690 49658 6806
rect 9 6582 49658 6690
rect 9 6466 49570 6582
rect 9 5798 49658 6466
rect 9 5682 49570 5798
rect 9 5350 49658 5682
rect 430 5234 49658 5350
rect 9 5014 49658 5234
rect 9 4898 49570 5014
rect 9 4230 49658 4898
rect 9 4114 49570 4230
rect 9 3894 49658 4114
rect 430 3778 49658 3894
rect 9 3446 49658 3778
rect 9 3330 49570 3446
rect 9 2438 49658 3330
rect 430 2322 49658 2438
rect 9 982 49658 2322
rect 430 866 49658 982
rect 9 462 49658 866
<< metal4 >>
rect 2224 1538 2384 48246
rect 9904 1538 10064 48246
rect 17584 1538 17744 48246
rect 25264 1538 25424 48246
rect 32944 1538 33104 48246
rect 40624 1538 40784 48246
rect 48304 1538 48464 48246
<< obsm4 >>
rect 1974 48276 48706 48935
rect 1974 1508 2194 48276
rect 2414 1508 9874 48276
rect 10094 1508 17554 48276
rect 17774 1508 25234 48276
rect 25454 1508 32914 48276
rect 33134 1508 40594 48276
rect 40814 1508 48274 48276
rect 48494 1508 48706 48276
rect 1974 457 48706 1508
<< labels >>
rlabel metal3 s 0 3808 400 3864 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 18368 400 18424 6 custom_settings[10]
port 2 nsew signal input
rlabel metal3 s 0 19824 400 19880 6 custom_settings[11]
port 3 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 custom_settings[12]
port 4 nsew signal input
rlabel metal3 s 0 22736 400 22792 6 custom_settings[13]
port 5 nsew signal input
rlabel metal3 s 0 24192 400 24248 6 custom_settings[14]
port 6 nsew signal input
rlabel metal3 s 0 25648 400 25704 6 custom_settings[15]
port 7 nsew signal input
rlabel metal3 s 0 27104 400 27160 6 custom_settings[16]
port 8 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 custom_settings[17]
port 9 nsew signal input
rlabel metal3 s 0 30016 400 30072 6 custom_settings[18]
port 10 nsew signal input
rlabel metal3 s 0 31472 400 31528 6 custom_settings[19]
port 11 nsew signal input
rlabel metal3 s 0 5264 400 5320 6 custom_settings[1]
port 12 nsew signal input
rlabel metal3 s 0 32928 400 32984 6 custom_settings[20]
port 13 nsew signal input
rlabel metal3 s 0 34384 400 34440 6 custom_settings[21]
port 14 nsew signal input
rlabel metal3 s 0 35840 400 35896 6 custom_settings[22]
port 15 nsew signal input
rlabel metal3 s 0 37296 400 37352 6 custom_settings[23]
port 16 nsew signal input
rlabel metal3 s 0 38752 400 38808 6 custom_settings[24]
port 17 nsew signal input
rlabel metal3 s 0 40208 400 40264 6 custom_settings[25]
port 18 nsew signal input
rlabel metal3 s 0 41664 400 41720 6 custom_settings[26]
port 19 nsew signal input
rlabel metal3 s 0 43120 400 43176 6 custom_settings[27]
port 20 nsew signal input
rlabel metal3 s 0 44576 400 44632 6 custom_settings[28]
port 21 nsew signal input
rlabel metal3 s 0 46032 400 46088 6 custom_settings[29]
port 22 nsew signal input
rlabel metal3 s 0 6720 400 6776 6 custom_settings[2]
port 23 nsew signal input
rlabel metal3 s 0 47488 400 47544 6 custom_settings[30]
port 24 nsew signal input
rlabel metal3 s 0 48944 400 49000 6 custom_settings[31]
port 25 nsew signal input
rlabel metal3 s 0 8176 400 8232 6 custom_settings[3]
port 26 nsew signal input
rlabel metal3 s 0 9632 400 9688 6 custom_settings[4]
port 27 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 custom_settings[5]
port 28 nsew signal input
rlabel metal3 s 0 12544 400 12600 6 custom_settings[6]
port 29 nsew signal input
rlabel metal3 s 0 14000 400 14056 6 custom_settings[7]
port 30 nsew signal input
rlabel metal3 s 0 15456 400 15512 6 custom_settings[8]
port 31 nsew signal input
rlabel metal3 s 0 16912 400 16968 6 custom_settings[9]
port 32 nsew signal input
rlabel metal2 s 3136 49600 3192 50000 6 io_in[0]
port 33 nsew signal input
rlabel metal2 s 9856 49600 9912 50000 6 io_in[10]
port 34 nsew signal input
rlabel metal2 s 10528 49600 10584 50000 6 io_in[11]
port 35 nsew signal input
rlabel metal2 s 11200 49600 11256 50000 6 io_in[12]
port 36 nsew signal input
rlabel metal2 s 11872 49600 11928 50000 6 io_in[13]
port 37 nsew signal input
rlabel metal2 s 12544 49600 12600 50000 6 io_in[14]
port 38 nsew signal input
rlabel metal2 s 13216 49600 13272 50000 6 io_in[15]
port 39 nsew signal input
rlabel metal2 s 13888 49600 13944 50000 6 io_in[16]
port 40 nsew signal input
rlabel metal2 s 14560 49600 14616 50000 6 io_in[17]
port 41 nsew signal input
rlabel metal2 s 15232 49600 15288 50000 6 io_in[18]
port 42 nsew signal input
rlabel metal2 s 15904 49600 15960 50000 6 io_in[19]
port 43 nsew signal input
rlabel metal2 s 3808 49600 3864 50000 6 io_in[1]
port 44 nsew signal input
rlabel metal2 s 16576 49600 16632 50000 6 io_in[20]
port 45 nsew signal input
rlabel metal2 s 17248 49600 17304 50000 6 io_in[21]
port 46 nsew signal input
rlabel metal2 s 17920 49600 17976 50000 6 io_in[22]
port 47 nsew signal input
rlabel metal2 s 18592 49600 18648 50000 6 io_in[23]
port 48 nsew signal input
rlabel metal2 s 19264 49600 19320 50000 6 io_in[24]
port 49 nsew signal input
rlabel metal2 s 19936 49600 19992 50000 6 io_in[25]
port 50 nsew signal input
rlabel metal2 s 20608 49600 20664 50000 6 io_in[26]
port 51 nsew signal input
rlabel metal2 s 21280 49600 21336 50000 6 io_in[27]
port 52 nsew signal input
rlabel metal2 s 21952 49600 22008 50000 6 io_in[28]
port 53 nsew signal input
rlabel metal2 s 22624 49600 22680 50000 6 io_in[29]
port 54 nsew signal input
rlabel metal2 s 4480 49600 4536 50000 6 io_in[2]
port 55 nsew signal input
rlabel metal2 s 23296 49600 23352 50000 6 io_in[30]
port 56 nsew signal input
rlabel metal2 s 23968 49600 24024 50000 6 io_in[31]
port 57 nsew signal input
rlabel metal2 s 24640 49600 24696 50000 6 io_in[32]
port 58 nsew signal input
rlabel metal2 s 5152 49600 5208 50000 6 io_in[3]
port 59 nsew signal input
rlabel metal2 s 5824 49600 5880 50000 6 io_in[4]
port 60 nsew signal input
rlabel metal2 s 6496 49600 6552 50000 6 io_in[5]
port 61 nsew signal input
rlabel metal2 s 7168 49600 7224 50000 6 io_in[6]
port 62 nsew signal input
rlabel metal2 s 7840 49600 7896 50000 6 io_in[7]
port 63 nsew signal input
rlabel metal2 s 8512 49600 8568 50000 6 io_in[8]
port 64 nsew signal input
rlabel metal2 s 9184 49600 9240 50000 6 io_in[9]
port 65 nsew signal input
rlabel metal3 s 49600 3360 50000 3416 6 io_oeb[0]
port 66 nsew signal output
rlabel metal3 s 49600 11200 50000 11256 6 io_oeb[10]
port 67 nsew signal output
rlabel metal3 s 49600 11984 50000 12040 6 io_oeb[11]
port 68 nsew signal output
rlabel metal3 s 49600 12768 50000 12824 6 io_oeb[12]
port 69 nsew signal output
rlabel metal3 s 49600 13552 50000 13608 6 io_oeb[13]
port 70 nsew signal output
rlabel metal3 s 49600 14336 50000 14392 6 io_oeb[14]
port 71 nsew signal output
rlabel metal3 s 49600 15120 50000 15176 6 io_oeb[15]
port 72 nsew signal output
rlabel metal3 s 49600 15904 50000 15960 6 io_oeb[16]
port 73 nsew signal output
rlabel metal3 s 49600 16688 50000 16744 6 io_oeb[17]
port 74 nsew signal output
rlabel metal3 s 49600 17472 50000 17528 6 io_oeb[18]
port 75 nsew signal output
rlabel metal3 s 49600 18256 50000 18312 6 io_oeb[19]
port 76 nsew signal output
rlabel metal3 s 49600 4144 50000 4200 6 io_oeb[1]
port 77 nsew signal output
rlabel metal3 s 49600 19040 50000 19096 6 io_oeb[20]
port 78 nsew signal output
rlabel metal3 s 49600 19824 50000 19880 6 io_oeb[21]
port 79 nsew signal output
rlabel metal3 s 49600 20608 50000 20664 6 io_oeb[22]
port 80 nsew signal output
rlabel metal3 s 49600 21392 50000 21448 6 io_oeb[23]
port 81 nsew signal output
rlabel metal3 s 49600 22176 50000 22232 6 io_oeb[24]
port 82 nsew signal output
rlabel metal3 s 49600 22960 50000 23016 6 io_oeb[25]
port 83 nsew signal output
rlabel metal3 s 49600 23744 50000 23800 6 io_oeb[26]
port 84 nsew signal output
rlabel metal3 s 49600 24528 50000 24584 6 io_oeb[27]
port 85 nsew signal output
rlabel metal3 s 49600 25312 50000 25368 6 io_oeb[28]
port 86 nsew signal output
rlabel metal3 s 49600 26096 50000 26152 6 io_oeb[29]
port 87 nsew signal output
rlabel metal3 s 49600 4928 50000 4984 6 io_oeb[2]
port 88 nsew signal output
rlabel metal3 s 49600 26880 50000 26936 6 io_oeb[30]
port 89 nsew signal output
rlabel metal3 s 49600 27664 50000 27720 6 io_oeb[31]
port 90 nsew signal output
rlabel metal3 s 49600 28448 50000 28504 6 io_oeb[32]
port 91 nsew signal output
rlabel metal3 s 49600 5712 50000 5768 6 io_oeb[3]
port 92 nsew signal output
rlabel metal3 s 49600 6496 50000 6552 6 io_oeb[4]
port 93 nsew signal output
rlabel metal3 s 49600 7280 50000 7336 6 io_oeb[5]
port 94 nsew signal output
rlabel metal3 s 49600 8064 50000 8120 6 io_oeb[6]
port 95 nsew signal output
rlabel metal3 s 49600 8848 50000 8904 6 io_oeb[7]
port 96 nsew signal output
rlabel metal3 s 49600 9632 50000 9688 6 io_oeb[8]
port 97 nsew signal output
rlabel metal3 s 49600 10416 50000 10472 6 io_oeb[9]
port 98 nsew signal output
rlabel metal2 s 25312 49600 25368 50000 6 io_out[0]
port 99 nsew signal output
rlabel metal2 s 32032 49600 32088 50000 6 io_out[10]
port 100 nsew signal output
rlabel metal2 s 32704 49600 32760 50000 6 io_out[11]
port 101 nsew signal output
rlabel metal2 s 33376 49600 33432 50000 6 io_out[12]
port 102 nsew signal output
rlabel metal2 s 34048 49600 34104 50000 6 io_out[13]
port 103 nsew signal output
rlabel metal2 s 34720 49600 34776 50000 6 io_out[14]
port 104 nsew signal output
rlabel metal2 s 35392 49600 35448 50000 6 io_out[15]
port 105 nsew signal output
rlabel metal2 s 36064 49600 36120 50000 6 io_out[16]
port 106 nsew signal output
rlabel metal2 s 36736 49600 36792 50000 6 io_out[17]
port 107 nsew signal output
rlabel metal2 s 37408 49600 37464 50000 6 io_out[18]
port 108 nsew signal output
rlabel metal2 s 38080 49600 38136 50000 6 io_out[19]
port 109 nsew signal output
rlabel metal2 s 25984 49600 26040 50000 6 io_out[1]
port 110 nsew signal output
rlabel metal2 s 38752 49600 38808 50000 6 io_out[20]
port 111 nsew signal output
rlabel metal2 s 39424 49600 39480 50000 6 io_out[21]
port 112 nsew signal output
rlabel metal2 s 40096 49600 40152 50000 6 io_out[22]
port 113 nsew signal output
rlabel metal2 s 40768 49600 40824 50000 6 io_out[23]
port 114 nsew signal output
rlabel metal2 s 41440 49600 41496 50000 6 io_out[24]
port 115 nsew signal output
rlabel metal2 s 42112 49600 42168 50000 6 io_out[25]
port 116 nsew signal output
rlabel metal2 s 42784 49600 42840 50000 6 io_out[26]
port 117 nsew signal output
rlabel metal2 s 43456 49600 43512 50000 6 io_out[27]
port 118 nsew signal output
rlabel metal2 s 44128 49600 44184 50000 6 io_out[28]
port 119 nsew signal output
rlabel metal2 s 44800 49600 44856 50000 6 io_out[29]
port 120 nsew signal output
rlabel metal2 s 26656 49600 26712 50000 6 io_out[2]
port 121 nsew signal output
rlabel metal2 s 45472 49600 45528 50000 6 io_out[30]
port 122 nsew signal output
rlabel metal2 s 46144 49600 46200 50000 6 io_out[31]
port 123 nsew signal output
rlabel metal2 s 46816 49600 46872 50000 6 io_out[32]
port 124 nsew signal output
rlabel metal2 s 27328 49600 27384 50000 6 io_out[3]
port 125 nsew signal output
rlabel metal2 s 28000 49600 28056 50000 6 io_out[4]
port 126 nsew signal output
rlabel metal2 s 28672 49600 28728 50000 6 io_out[5]
port 127 nsew signal output
rlabel metal2 s 29344 49600 29400 50000 6 io_out[6]
port 128 nsew signal output
rlabel metal2 s 30016 49600 30072 50000 6 io_out[7]
port 129 nsew signal output
rlabel metal2 s 30688 49600 30744 50000 6 io_out[8]
port 130 nsew signal output
rlabel metal2 s 31360 49600 31416 50000 6 io_out[9]
port 131 nsew signal output
rlabel metal3 s 0 2352 400 2408 6 rst_n
port 132 nsew signal input
rlabel metal3 s 49600 29232 50000 29288 6 sram_addr[0]
port 133 nsew signal output
rlabel metal3 s 49600 30016 50000 30072 6 sram_addr[1]
port 134 nsew signal output
rlabel metal3 s 49600 30800 50000 30856 6 sram_addr[2]
port 135 nsew signal output
rlabel metal3 s 49600 31584 50000 31640 6 sram_addr[3]
port 136 nsew signal output
rlabel metal3 s 49600 32368 50000 32424 6 sram_addr[4]
port 137 nsew signal output
rlabel metal3 s 49600 33152 50000 33208 6 sram_addr[5]
port 138 nsew signal output
rlabel metal3 s 49600 46480 50000 46536 6 sram_gwe
port 139 nsew signal output
rlabel metal3 s 49600 33936 50000 33992 6 sram_in[0]
port 140 nsew signal output
rlabel metal3 s 49600 34720 50000 34776 6 sram_in[1]
port 141 nsew signal output
rlabel metal3 s 49600 35504 50000 35560 6 sram_in[2]
port 142 nsew signal output
rlabel metal3 s 49600 36288 50000 36344 6 sram_in[3]
port 143 nsew signal output
rlabel metal3 s 49600 37072 50000 37128 6 sram_in[4]
port 144 nsew signal output
rlabel metal3 s 49600 37856 50000 37912 6 sram_in[5]
port 145 nsew signal output
rlabel metal3 s 49600 38640 50000 38696 6 sram_in[6]
port 146 nsew signal output
rlabel metal3 s 49600 39424 50000 39480 6 sram_in[7]
port 147 nsew signal output
rlabel metal3 s 49600 40208 50000 40264 6 sram_out[0]
port 148 nsew signal input
rlabel metal3 s 49600 40992 50000 41048 6 sram_out[1]
port 149 nsew signal input
rlabel metal3 s 49600 41776 50000 41832 6 sram_out[2]
port 150 nsew signal input
rlabel metal3 s 49600 42560 50000 42616 6 sram_out[3]
port 151 nsew signal input
rlabel metal3 s 49600 43344 50000 43400 6 sram_out[4]
port 152 nsew signal input
rlabel metal3 s 49600 44128 50000 44184 6 sram_out[5]
port 153 nsew signal input
rlabel metal3 s 49600 44912 50000 44968 6 sram_out[6]
port 154 nsew signal input
rlabel metal3 s 49600 45696 50000 45752 6 sram_out[7]
port 155 nsew signal input
rlabel metal4 s 2224 1538 2384 48246 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 48246 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 48246 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 48246 6 vdd
port 156 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 48246 6 vss
port 157 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 48246 6 vss
port 157 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 48246 6 vss
port 157 nsew ground bidirectional
rlabel metal3 s 0 896 400 952 6 wb_clk_i
port 158 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10532446
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1_group/openlane/wrapped_qcpu/runs/23_11_03_02_02/results/signoff/wrapped_qcpu.magic.gds
string GDS_START 505248
<< end >>

