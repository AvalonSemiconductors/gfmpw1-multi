magic
tech gf180mcuD
magscale 1 10
timestamp 1712520156
<< nwell >>
rect 1258 156423 40798 156448
rect 1258 155609 228678 156423
rect 1258 155584 34764 155609
rect 1258 154855 35956 154880
rect 1258 154041 228678 154855
rect 1258 154016 25720 154041
rect 1258 153287 28217 153312
rect 1258 152473 228678 153287
rect 1258 152448 24782 152473
rect 1258 151719 23663 151744
rect 1258 150905 228678 151719
rect 1258 150880 13981 150905
rect 1258 150151 15878 150176
rect 1258 149337 228678 150151
rect 1258 149312 15225 149337
rect 1258 148583 13064 148608
rect 1258 147769 228678 148583
rect 1258 147744 10908 147769
rect 1258 147015 10502 147040
rect 1258 146201 228678 147015
rect 1258 146176 7823 146201
rect 1258 145447 5896 145472
rect 1258 144633 228678 145447
rect 1258 144608 8024 144633
rect 1258 143879 4799 143904
rect 1258 143065 228678 143879
rect 1258 143040 15103 143065
rect 1258 142311 14870 142336
rect 1258 141497 228678 142311
rect 1258 141472 2760 141497
rect 1258 140743 4140 140768
rect 1258 139929 228678 140743
rect 1258 139904 6680 139929
rect 1258 139175 3180 139200
rect 1258 138361 228678 139175
rect 1258 138336 6358 138361
rect 1258 137607 2437 137632
rect 1258 136793 228678 137607
rect 1258 136768 7030 136793
rect 1258 136039 15710 136064
rect 1258 135225 228678 136039
rect 1258 135200 15206 135225
rect 1258 134471 7478 134496
rect 1258 133657 228678 134471
rect 1258 133632 18342 133657
rect 1258 132903 4239 132928
rect 1258 132089 228678 132903
rect 1258 132064 2662 132089
rect 1258 131335 3117 131360
rect 1258 130521 228678 131335
rect 1258 130496 3166 130521
rect 1258 129767 26415 129792
rect 1258 128953 228678 129767
rect 1258 128928 4734 128953
rect 1258 128199 1887 128224
rect 1258 127385 228678 128199
rect 1258 127360 11293 127385
rect 1258 126631 1878 126656
rect 1258 125817 228678 126631
rect 1258 125792 3455 125817
rect 1258 125063 41983 125088
rect 1258 124249 228678 125063
rect 1258 124224 7646 124249
rect 1258 123495 2893 123520
rect 1258 122681 228678 123495
rect 1258 122656 17343 122681
rect 1258 121927 4622 121952
rect 1258 121113 228678 121927
rect 1258 121088 2895 121113
rect 1258 120359 4118 120384
rect 1258 119545 228678 120359
rect 1258 119520 14197 119545
rect 1258 118791 27414 118816
rect 1258 117977 228678 118791
rect 1258 117952 13638 117977
rect 1258 117223 6582 117248
rect 1258 116409 228678 117223
rect 1258 116384 33013 116409
rect 1258 115655 13750 115680
rect 1258 114841 228678 115655
rect 1258 114816 9942 114841
rect 1258 114087 5631 114112
rect 1258 113273 228678 114087
rect 1258 113248 7870 113273
rect 1258 112519 3404 112544
rect 1258 111705 228678 112519
rect 1258 111680 11454 111705
rect 1258 110951 5483 110976
rect 1258 110137 228678 110951
rect 1258 110112 5927 110137
rect 1258 109383 4461 109408
rect 1258 108569 228678 109383
rect 1258 108544 4174 108569
rect 1258 107815 3592 107840
rect 1258 107001 228678 107815
rect 1258 106976 10493 107001
rect 1258 106247 36701 106272
rect 1258 105433 228678 106247
rect 1258 105408 25277 105433
rect 1258 104679 3592 104704
rect 1258 103865 228678 104679
rect 1258 103840 18440 103865
rect 1258 103111 14189 103136
rect 1258 102297 228678 103111
rect 1258 102272 6589 102297
rect 1258 101543 37949 101568
rect 1258 100729 228678 101543
rect 1258 100704 3565 100729
rect 1258 99975 3592 100000
rect 1258 99161 228678 99975
rect 1258 99136 16653 99161
rect 1258 98407 3278 98432
rect 1258 97593 228678 98407
rect 1258 97568 30541 97593
rect 1258 96839 14366 96864
rect 1258 96025 228678 96839
rect 1258 96000 6652 96025
rect 1258 95271 10421 95296
rect 1258 94457 228678 95271
rect 1258 94432 14268 94457
rect 1258 93703 22951 93728
rect 1258 92889 228678 93703
rect 1258 92864 45614 92889
rect 1258 92135 5901 92160
rect 1258 91321 228678 92135
rect 1258 91296 55069 91321
rect 1258 90567 2541 90592
rect 1258 89753 228678 90567
rect 1258 89728 25165 89753
rect 1258 88999 35469 89024
rect 1258 88185 228678 88999
rect 1258 88160 2765 88185
rect 1258 87431 10334 87456
rect 1258 86617 228678 87431
rect 1258 86592 17032 86617
rect 1258 85863 2942 85888
rect 1258 85049 228678 85863
rect 1258 85024 7142 85049
rect 1258 84295 19909 84320
rect 1258 83481 228678 84295
rect 1258 83456 18583 83481
rect 1258 82727 19272 82752
rect 1258 81913 228678 82727
rect 1258 81888 49478 81913
rect 1258 81159 6573 81184
rect 1258 80345 228678 81159
rect 1258 80320 10045 80345
rect 1258 79591 6573 79616
rect 1258 78777 228678 79591
rect 1258 78752 2989 78777
rect 1258 78023 12397 78048
rect 1258 77209 228678 78023
rect 1258 77184 2541 77209
rect 1258 76455 11544 76480
rect 1258 75641 228678 76455
rect 1258 75616 19272 75641
rect 1258 74887 14749 74912
rect 1258 74073 228678 74887
rect 1258 74048 8271 74073
rect 1258 73319 14982 73344
rect 1258 72505 228678 73319
rect 1258 72480 19014 72505
rect 1258 71751 5250 71776
rect 1258 70937 228678 71751
rect 1258 70912 11902 70937
rect 1258 70183 2214 70208
rect 1258 69369 228678 70183
rect 1258 69344 26014 69369
rect 1258 68615 11566 68640
rect 1258 67801 228678 68615
rect 1258 67776 17119 67801
rect 1258 67047 42142 67072
rect 1258 66233 228678 67047
rect 1258 66208 14254 66233
rect 1258 65479 6701 65504
rect 1258 64665 228678 65479
rect 1258 64640 2214 64665
rect 1258 63911 39678 63936
rect 1258 63097 228678 63911
rect 1258 63072 2214 63097
rect 1258 62343 3894 62368
rect 1258 61529 228678 62343
rect 1258 61504 39501 61529
rect 1258 60775 6694 60800
rect 1258 59961 228678 60775
rect 1258 59936 50520 59961
rect 1258 59207 43569 59232
rect 1258 58393 228678 59207
rect 1258 58368 6358 58393
rect 1258 57639 6703 57664
rect 1258 56825 228678 57639
rect 1258 56800 21836 56825
rect 1258 56071 2326 56096
rect 1258 55257 228678 56071
rect 1258 55232 3351 55257
rect 1258 54503 41741 54528
rect 1258 53689 228678 54503
rect 1258 53664 9718 53689
rect 1258 52935 13984 52960
rect 1258 52121 228678 52935
rect 1258 52096 25977 52121
rect 1258 51367 7758 51392
rect 1258 50553 228678 51367
rect 1258 50528 43457 50553
rect 1258 49799 21693 49824
rect 1258 48985 228678 49799
rect 1258 48960 3592 48985
rect 1258 48231 6461 48256
rect 1258 47417 228678 48231
rect 1258 47392 6461 47417
rect 1258 46663 2541 46688
rect 1258 45849 228678 46663
rect 1258 45824 6461 45849
rect 1258 45095 38312 45120
rect 1258 44281 228678 45095
rect 1258 44256 17101 44281
rect 1258 43527 2541 43552
rect 1258 42713 228678 43527
rect 1258 42688 6461 42713
rect 1258 41959 76828 41984
rect 1258 41145 228678 41959
rect 1258 41120 9821 41145
rect 1258 40391 5789 40416
rect 1258 39577 228678 40391
rect 1258 39552 9597 39577
rect 1258 38823 13069 38848
rect 1258 38009 228678 38823
rect 1258 37984 16653 38009
rect 1258 37255 22072 37280
rect 1258 36441 228678 37255
rect 1258 36416 10829 36441
rect 1258 35687 36296 35712
rect 1258 34873 228678 35687
rect 1258 34848 9752 34873
rect 1258 34119 12285 34144
rect 1258 33305 228678 34119
rect 1258 33280 39725 33305
rect 1258 32551 11501 32576
rect 1258 31737 228678 32551
rect 1258 31712 7469 31737
rect 1258 30983 27965 31008
rect 1258 30169 228678 30983
rect 1258 30144 9261 30169
rect 1258 29415 27414 29440
rect 1258 28601 228678 29415
rect 1258 28576 6461 28601
rect 1258 27847 10381 27872
rect 1258 27033 228678 27847
rect 1258 27008 35400 27033
rect 1258 26279 27741 26304
rect 1258 25465 228678 26279
rect 1258 25440 9933 25465
rect 1258 24711 30429 24736
rect 1258 23897 228678 24711
rect 1258 23872 7736 23897
rect 1258 23143 18221 23168
rect 1258 22329 228678 23143
rect 1258 22304 14301 22329
rect 1258 21575 18557 21600
rect 1258 20761 228678 21575
rect 1258 20736 14525 20761
rect 1258 20007 12621 20032
rect 1258 19193 228678 20007
rect 1258 19168 32781 19193
rect 1258 18439 14637 18464
rect 1258 17625 228678 18439
rect 1258 17600 25320 17625
rect 1258 16871 62840 16896
rect 1258 16057 228678 16871
rect 1258 16032 11880 16057
rect 1258 15303 28749 15328
rect 1258 14489 228678 15303
rect 1258 14464 23057 14489
rect 1258 13735 14189 13760
rect 1258 12921 228678 13735
rect 1258 12896 17101 12921
rect 1258 12167 62280 12192
rect 1258 11353 228678 12167
rect 1258 11328 16653 11353
rect 1258 10599 20237 10624
rect 1258 9785 228678 10599
rect 1258 9760 38420 9785
rect 1258 9031 20125 9056
rect 1258 8217 228678 9031
rect 1258 8192 32669 8217
rect 1258 7463 27965 7488
rect 1258 6649 228678 7463
rect 1258 6624 18669 6649
rect 1258 5895 22589 5920
rect 1258 5081 228678 5895
rect 1258 5056 39277 5081
rect 1258 4327 36365 4352
rect 1258 3513 228678 4327
rect 1258 3488 82509 3513
<< pwell >>
rect 1258 156448 228678 156886
rect 1258 154880 228678 155584
rect 1258 153312 228678 154016
rect 1258 151744 228678 152448
rect 1258 150176 228678 150880
rect 1258 148608 228678 149312
rect 1258 147040 228678 147744
rect 1258 145472 228678 146176
rect 1258 143904 228678 144608
rect 1258 142336 228678 143040
rect 1258 140768 228678 141472
rect 1258 139200 228678 139904
rect 1258 137632 228678 138336
rect 1258 136064 228678 136768
rect 1258 134496 228678 135200
rect 1258 132928 228678 133632
rect 1258 131360 228678 132064
rect 1258 129792 228678 130496
rect 1258 128224 228678 128928
rect 1258 126656 228678 127360
rect 1258 125088 228678 125792
rect 1258 123520 228678 124224
rect 1258 121952 228678 122656
rect 1258 120384 228678 121088
rect 1258 118816 228678 119520
rect 1258 117248 228678 117952
rect 1258 115680 228678 116384
rect 1258 114112 228678 114816
rect 1258 112544 228678 113248
rect 1258 110976 228678 111680
rect 1258 109408 228678 110112
rect 1258 107840 228678 108544
rect 1258 106272 228678 106976
rect 1258 104704 228678 105408
rect 1258 103136 228678 103840
rect 1258 101568 228678 102272
rect 1258 100000 228678 100704
rect 1258 98432 228678 99136
rect 1258 96864 228678 97568
rect 1258 95296 228678 96000
rect 1258 93728 228678 94432
rect 1258 92160 228678 92864
rect 1258 90592 228678 91296
rect 1258 89024 228678 89728
rect 1258 87456 228678 88160
rect 1258 85888 228678 86592
rect 1258 84320 228678 85024
rect 1258 82752 228678 83456
rect 1258 81184 228678 81888
rect 1258 79616 228678 80320
rect 1258 78048 228678 78752
rect 1258 76480 228678 77184
rect 1258 74912 228678 75616
rect 1258 73344 228678 74048
rect 1258 71776 228678 72480
rect 1258 70208 228678 70912
rect 1258 68640 228678 69344
rect 1258 67072 228678 67776
rect 1258 65504 228678 66208
rect 1258 63936 228678 64640
rect 1258 62368 228678 63072
rect 1258 60800 228678 61504
rect 1258 59232 228678 59936
rect 1258 57664 228678 58368
rect 1258 56096 228678 56800
rect 1258 54528 228678 55232
rect 1258 52960 228678 53664
rect 1258 51392 228678 52096
rect 1258 49824 228678 50528
rect 1258 48256 228678 48960
rect 1258 46688 228678 47392
rect 1258 45120 228678 45824
rect 1258 43552 228678 44256
rect 1258 41984 228678 42688
rect 1258 40416 228678 41120
rect 1258 38848 228678 39552
rect 1258 37280 228678 37984
rect 1258 35712 228678 36416
rect 1258 34144 228678 34848
rect 1258 32576 228678 33280
rect 1258 31008 228678 31712
rect 1258 29440 228678 30144
rect 1258 27872 228678 28576
rect 1258 26304 228678 27008
rect 1258 24736 228678 25440
rect 1258 23168 228678 23872
rect 1258 21600 228678 22304
rect 1258 20032 228678 20736
rect 1258 18464 228678 19168
rect 1258 16896 228678 17600
rect 1258 15328 228678 16032
rect 1258 13760 228678 14464
rect 1258 12192 228678 12896
rect 1258 10624 228678 11328
rect 1258 9056 228678 9760
rect 1258 7488 228678 8192
rect 1258 5920 228678 6624
rect 1258 4352 228678 5056
rect 1258 3050 228678 3488
<< obsm1 >>
rect 1344 3076 228592 156860
<< metal2 >>
rect 114912 159200 115024 160000
rect 57344 0 57456 800
rect 172256 0 172368 800
<< obsm2 >>
rect 1484 159140 114852 159200
rect 115084 159140 228564 159200
rect 1484 860 228564 159140
rect 1484 700 57284 860
rect 57516 700 172196 860
rect 172428 700 228564 860
<< metal3 >>
rect 229200 157024 230000 157136
rect 229200 154112 230000 154224
rect 229200 151200 230000 151312
rect 229200 148288 230000 148400
rect 229200 145376 230000 145488
rect 229200 142464 230000 142576
rect 229200 139552 230000 139664
rect 229200 136640 230000 136752
rect 229200 133728 230000 133840
rect 229200 130816 230000 130928
rect 229200 127904 230000 128016
rect 229200 124992 230000 125104
rect 229200 122080 230000 122192
rect 229200 119168 230000 119280
rect 229200 116256 230000 116368
rect 229200 113344 230000 113456
rect 229200 110432 230000 110544
rect 229200 107520 230000 107632
rect 229200 104608 230000 104720
rect 229200 101696 230000 101808
rect 229200 98784 230000 98896
rect 229200 95872 230000 95984
rect 229200 92960 230000 93072
rect 229200 90048 230000 90160
rect 229200 87136 230000 87248
rect 229200 84224 230000 84336
rect 229200 81312 230000 81424
rect 229200 78400 230000 78512
rect 229200 75488 230000 75600
rect 229200 72576 230000 72688
rect 229200 69664 230000 69776
rect 229200 66752 230000 66864
rect 229200 63840 230000 63952
rect 229200 60928 230000 61040
rect 229200 58016 230000 58128
rect 229200 55104 230000 55216
rect 229200 52192 230000 52304
rect 229200 49280 230000 49392
rect 229200 46368 230000 46480
rect 229200 43456 230000 43568
rect 229200 40544 230000 40656
rect 229200 37632 230000 37744
rect 229200 34720 230000 34832
rect 229200 31808 230000 31920
rect 229200 28896 230000 29008
rect 229200 25984 230000 26096
rect 229200 23072 230000 23184
rect 229200 20160 230000 20272
rect 229200 17248 230000 17360
rect 229200 14336 230000 14448
rect 229200 11424 230000 11536
rect 229200 8512 230000 8624
rect 229200 5600 230000 5712
rect 229200 2688 230000 2800
<< obsm3 >>
rect 1474 157196 229200 158676
rect 1474 156964 229140 157196
rect 1474 154284 229200 156964
rect 1474 154052 229140 154284
rect 1474 151372 229200 154052
rect 1474 151140 229140 151372
rect 1474 148460 229200 151140
rect 1474 148228 229140 148460
rect 1474 145548 229200 148228
rect 1474 145316 229140 145548
rect 1474 142636 229200 145316
rect 1474 142404 229140 142636
rect 1474 139724 229200 142404
rect 1474 139492 229140 139724
rect 1474 136812 229200 139492
rect 1474 136580 229140 136812
rect 1474 133900 229200 136580
rect 1474 133668 229140 133900
rect 1474 130988 229200 133668
rect 1474 130756 229140 130988
rect 1474 128076 229200 130756
rect 1474 127844 229140 128076
rect 1474 125164 229200 127844
rect 1474 124932 229140 125164
rect 1474 122252 229200 124932
rect 1474 122020 229140 122252
rect 1474 119340 229200 122020
rect 1474 119108 229140 119340
rect 1474 116428 229200 119108
rect 1474 116196 229140 116428
rect 1474 113516 229200 116196
rect 1474 113284 229140 113516
rect 1474 110604 229200 113284
rect 1474 110372 229140 110604
rect 1474 107692 229200 110372
rect 1474 107460 229140 107692
rect 1474 104780 229200 107460
rect 1474 104548 229140 104780
rect 1474 101868 229200 104548
rect 1474 101636 229140 101868
rect 1474 98956 229200 101636
rect 1474 98724 229140 98956
rect 1474 96044 229200 98724
rect 1474 95812 229140 96044
rect 1474 93132 229200 95812
rect 1474 92900 229140 93132
rect 1474 90220 229200 92900
rect 1474 89988 229140 90220
rect 1474 87308 229200 89988
rect 1474 87076 229140 87308
rect 1474 84396 229200 87076
rect 1474 84164 229140 84396
rect 1474 81484 229200 84164
rect 1474 81252 229140 81484
rect 1474 78572 229200 81252
rect 1474 78340 229140 78572
rect 1474 75660 229200 78340
rect 1474 75428 229140 75660
rect 1474 72748 229200 75428
rect 1474 72516 229140 72748
rect 1474 69836 229200 72516
rect 1474 69604 229140 69836
rect 1474 66924 229200 69604
rect 1474 66692 229140 66924
rect 1474 64012 229200 66692
rect 1474 63780 229140 64012
rect 1474 61100 229200 63780
rect 1474 60868 229140 61100
rect 1474 58188 229200 60868
rect 1474 57956 229140 58188
rect 1474 55276 229200 57956
rect 1474 55044 229140 55276
rect 1474 52364 229200 55044
rect 1474 52132 229140 52364
rect 1474 49452 229200 52132
rect 1474 49220 229140 49452
rect 1474 46540 229200 49220
rect 1474 46308 229140 46540
rect 1474 43628 229200 46308
rect 1474 43396 229140 43628
rect 1474 40716 229200 43396
rect 1474 40484 229140 40716
rect 1474 37804 229200 40484
rect 1474 37572 229140 37804
rect 1474 34892 229200 37572
rect 1474 34660 229140 34892
rect 1474 31980 229200 34660
rect 1474 31748 229140 31980
rect 1474 29068 229200 31748
rect 1474 28836 229140 29068
rect 1474 26156 229200 28836
rect 1474 25924 229140 26156
rect 1474 23244 229200 25924
rect 1474 23012 229140 23244
rect 1474 20332 229200 23012
rect 1474 20100 229140 20332
rect 1474 17420 229200 20100
rect 1474 17188 229140 17420
rect 1474 14508 229200 17188
rect 1474 14276 229140 14508
rect 1474 11596 229200 14276
rect 1474 11364 229140 11596
rect 1474 8684 229200 11364
rect 1474 8452 229140 8684
rect 1474 5772 229200 8452
rect 1474 5540 229140 5772
rect 1474 2860 229200 5540
rect 1474 2628 229140 2860
rect 1474 812 229200 2628
<< metal4 >>
rect 4448 3076 4768 156860
rect 19808 3076 20128 156860
rect 35168 3076 35488 156860
rect 50528 3076 50848 156860
rect 65888 3076 66208 156860
rect 81248 3076 81568 156860
rect 96608 3076 96928 156860
rect 111968 3076 112288 156860
rect 127328 3076 127648 156860
rect 142688 3076 143008 156860
rect 158048 3076 158368 156860
rect 173408 3076 173728 156860
rect 188768 3076 189088 156860
rect 204128 3076 204448 156860
rect 219488 3076 219808 156860
<< obsm4 >>
rect 4284 156920 226772 158462
rect 4284 3016 4388 156920
rect 4828 3016 19748 156920
rect 20188 3016 35108 156920
rect 35548 3016 50468 156920
rect 50908 3016 65828 156920
rect 66268 3016 81188 156920
rect 81628 3016 96548 156920
rect 96988 3016 111908 156920
rect 112348 3016 127268 156920
rect 127708 3016 142628 156920
rect 143068 3016 157988 156920
rect 158428 3016 173348 156920
rect 173788 3016 188708 156920
rect 189148 3016 204068 156920
rect 204508 3016 219428 156920
rect 219868 3016 226772 156920
rect 4284 1026 226772 3016
<< labels >>
rlabel metal3 s 229200 2688 230000 2800 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 229200 31808 230000 31920 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 229200 34720 230000 34832 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 229200 37632 230000 37744 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 229200 40544 230000 40656 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 229200 43456 230000 43568 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 229200 46368 230000 46480 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 229200 49280 230000 49392 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 229200 52192 230000 52304 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 229200 55104 230000 55216 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 229200 58016 230000 58128 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 229200 5600 230000 5712 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 229200 60928 230000 61040 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 229200 63840 230000 63952 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 229200 66752 230000 66864 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 229200 69664 230000 69776 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 229200 72576 230000 72688 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 229200 75488 230000 75600 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 229200 78400 230000 78512 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 229200 81312 230000 81424 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 229200 84224 230000 84336 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 229200 87136 230000 87248 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 229200 8512 230000 8624 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 229200 90048 230000 90160 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 229200 92960 230000 93072 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 229200 95872 230000 95984 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 229200 11424 230000 11536 6 io_in[3]
port 27 nsew signal input
rlabel metal3 s 229200 14336 230000 14448 6 io_in[4]
port 28 nsew signal input
rlabel metal3 s 229200 17248 230000 17360 6 io_in[5]
port 29 nsew signal input
rlabel metal3 s 229200 20160 230000 20272 6 io_in[6]
port 30 nsew signal input
rlabel metal3 s 229200 23072 230000 23184 6 io_in[7]
port 31 nsew signal input
rlabel metal3 s 229200 25984 230000 26096 6 io_in[8]
port 32 nsew signal input
rlabel metal3 s 229200 28896 230000 29008 6 io_in[9]
port 33 nsew signal input
rlabel metal2 s 114912 159200 115024 160000 6 io_oeb
port 34 nsew signal output
rlabel metal3 s 229200 98784 230000 98896 6 io_out[0]
port 35 nsew signal output
rlabel metal3 s 229200 127904 230000 128016 6 io_out[10]
port 36 nsew signal output
rlabel metal3 s 229200 130816 230000 130928 6 io_out[11]
port 37 nsew signal output
rlabel metal3 s 229200 133728 230000 133840 6 io_out[12]
port 38 nsew signal output
rlabel metal3 s 229200 136640 230000 136752 6 io_out[13]
port 39 nsew signal output
rlabel metal3 s 229200 139552 230000 139664 6 io_out[14]
port 40 nsew signal output
rlabel metal3 s 229200 142464 230000 142576 6 io_out[15]
port 41 nsew signal output
rlabel metal3 s 229200 145376 230000 145488 6 io_out[16]
port 42 nsew signal output
rlabel metal3 s 229200 148288 230000 148400 6 io_out[17]
port 43 nsew signal output
rlabel metal3 s 229200 151200 230000 151312 6 io_out[18]
port 44 nsew signal output
rlabel metal3 s 229200 154112 230000 154224 6 io_out[19]
port 45 nsew signal output
rlabel metal3 s 229200 101696 230000 101808 6 io_out[1]
port 46 nsew signal output
rlabel metal3 s 229200 157024 230000 157136 6 io_out[20]
port 47 nsew signal output
rlabel metal3 s 229200 104608 230000 104720 6 io_out[2]
port 48 nsew signal output
rlabel metal3 s 229200 107520 230000 107632 6 io_out[3]
port 49 nsew signal output
rlabel metal3 s 229200 110432 230000 110544 6 io_out[4]
port 50 nsew signal output
rlabel metal3 s 229200 113344 230000 113456 6 io_out[5]
port 51 nsew signal output
rlabel metal3 s 229200 116256 230000 116368 6 io_out[6]
port 52 nsew signal output
rlabel metal3 s 229200 119168 230000 119280 6 io_out[7]
port 53 nsew signal output
rlabel metal3 s 229200 122080 230000 122192 6 io_out[8]
port 54 nsew signal output
rlabel metal3 s 229200 124992 230000 125104 6 io_out[9]
port 55 nsew signal output
rlabel metal2 s 172256 0 172368 800 6 rst_n
port 56 nsew signal input
rlabel metal4 s 4448 3076 4768 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 156860 6 vdd
port 57 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 156860 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 156860 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 156860 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 156860 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 156860 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 156860 6 vss
port 58 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 156860 6 vss
port 58 nsew ground bidirectional
rlabel metal2 s 57344 0 57456 800 6 wb_clk_i
port 59 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 230000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30451236
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_sid/runs/24_04_07_21_29/results/signoff/wrapped_sid.magic.gds
string GDS_START 541024
<< end >>

