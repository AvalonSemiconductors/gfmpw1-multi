VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avali_logo
  CLASS BLOCK ;
  FOREIGN avali_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 469.600 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 150.400 322.400 172.000 323.200 ;
        RECT 142.400 321.600 182.400 322.400 ;
        RECT 136.000 320.800 190.400 321.600 ;
        RECT 132.000 320.000 196.000 320.800 ;
        RECT 128.000 319.200 196.000 320.000 ;
        RECT 124.000 318.400 195.200 319.200 ;
        RECT 120.800 317.600 195.200 318.400 ;
        RECT 118.400 316.800 194.400 317.600 ;
        RECT 115.200 316.000 194.400 316.800 ;
        RECT 112.800 315.200 193.600 316.000 ;
        RECT 110.400 314.400 193.600 315.200 ;
        RECT 108.000 313.600 192.800 314.400 ;
        RECT 105.600 312.800 192.000 313.600 ;
        RECT 104.000 312.000 192.000 312.800 ;
        RECT 101.600 311.200 191.200 312.000 ;
        RECT 100.000 310.400 191.200 311.200 ;
        RECT 97.600 309.600 190.400 310.400 ;
        RECT 96.000 308.800 190.400 309.600 ;
        RECT 94.400 308.000 189.600 308.800 ;
        RECT 92.800 307.200 189.600 308.000 ;
        RECT 91.200 306.400 188.800 307.200 ;
        RECT 89.600 305.600 188.800 306.400 ;
        RECT 88.000 304.800 188.000 305.600 ;
        RECT 86.400 304.000 188.000 304.800 ;
        RECT 84.800 303.200 187.200 304.000 ;
        RECT 83.200 302.400 186.400 303.200 ;
        RECT 81.600 301.600 186.400 302.400 ;
        RECT 80.000 300.800 185.600 301.600 ;
        RECT 79.200 300.000 185.600 300.800 ;
        RECT 77.600 299.200 184.800 300.000 ;
        RECT 76.800 298.400 184.800 299.200 ;
        RECT 75.200 297.600 184.000 298.400 ;
        RECT 73.600 296.800 184.000 297.600 ;
        RECT 72.800 296.000 183.200 296.800 ;
        RECT 71.200 295.200 183.200 296.000 ;
        RECT 70.400 294.400 148.800 295.200 ;
        RECT 176.800 294.400 182.400 295.200 ;
        RECT 68.800 293.600 142.400 294.400 ;
        RECT 68.000 292.800 137.600 293.600 ;
        RECT 67.200 292.000 133.600 292.800 ;
        RECT 65.600 291.200 130.400 292.000 ;
        RECT 64.800 290.400 127.200 291.200 ;
        RECT 64.000 289.600 124.000 290.400 ;
        RECT 62.400 288.800 121.600 289.600 ;
        RECT 61.600 288.000 119.200 288.800 ;
        RECT 60.800 287.200 116.800 288.000 ;
        RECT 59.200 286.400 114.400 287.200 ;
        RECT 58.400 285.600 112.800 286.400 ;
        RECT 57.600 284.800 110.400 285.600 ;
        RECT 56.800 284.000 108.800 284.800 ;
        RECT 56.000 283.200 107.200 284.000 ;
        RECT 55.200 282.400 104.800 283.200 ;
        RECT 53.600 281.600 103.200 282.400 ;
        RECT 52.800 280.800 101.600 281.600 ;
        RECT 52.000 280.000 100.000 280.800 ;
        RECT 51.200 279.200 98.400 280.000 ;
        RECT 50.400 278.400 97.600 279.200 ;
        RECT 49.600 277.600 96.000 278.400 ;
        RECT 48.800 276.800 94.400 277.600 ;
        RECT 48.000 276.000 92.800 276.800 ;
        RECT 47.200 275.200 92.000 276.000 ;
        RECT 46.400 274.400 90.400 275.200 ;
        RECT 45.600 273.600 89.600 274.400 ;
        RECT 44.800 272.800 88.000 273.600 ;
        RECT 44.000 272.000 86.400 272.800 ;
        RECT 43.200 271.200 85.600 272.000 ;
        RECT 42.400 270.400 84.800 271.200 ;
        RECT 41.600 269.600 83.200 270.400 ;
        RECT 41.600 268.800 82.400 269.600 ;
        RECT 40.800 268.000 80.800 268.800 ;
        RECT 40.000 267.200 80.000 268.000 ;
        RECT 39.200 266.400 79.200 267.200 ;
        RECT 38.400 265.600 78.400 266.400 ;
        RECT 37.600 264.800 76.800 265.600 ;
        RECT 36.800 264.000 76.000 264.800 ;
        RECT 36.800 263.200 75.200 264.000 ;
        RECT 36.000 262.400 74.400 263.200 ;
        RECT 35.200 261.600 73.600 262.400 ;
        RECT 34.400 260.800 72.800 261.600 ;
        RECT 33.600 260.000 71.200 260.800 ;
        RECT 33.600 259.200 70.400 260.000 ;
        RECT 32.800 258.400 69.600 259.200 ;
        RECT 32.000 257.600 68.800 258.400 ;
        RECT 31.200 256.800 68.000 257.600 ;
        RECT 31.200 256.000 67.200 256.800 ;
        RECT 30.400 255.200 66.400 256.000 ;
        RECT 29.600 254.400 65.600 255.200 ;
        RECT 29.600 253.600 64.800 254.400 ;
        RECT 28.800 252.800 64.000 253.600 ;
        RECT 28.000 252.000 63.200 252.800 ;
        RECT 27.200 250.400 62.400 252.000 ;
        RECT 26.400 249.600 61.600 250.400 ;
        RECT 26.400 248.800 60.800 249.600 ;
        RECT 25.600 248.000 60.000 248.800 ;
        RECT 24.800 247.200 59.200 248.000 ;
        RECT 24.800 246.400 58.400 247.200 ;
        RECT 24.000 245.600 57.600 246.400 ;
        RECT 23.200 244.800 57.600 245.600 ;
        RECT 23.200 244.000 56.800 244.800 ;
        RECT 22.400 243.200 56.000 244.000 ;
        RECT 22.400 242.400 55.200 243.200 ;
        RECT 21.600 241.600 55.200 242.400 ;
        RECT 20.800 240.800 54.400 241.600 ;
        RECT 20.800 240.000 53.600 240.800 ;
        RECT 20.000 238.400 52.800 240.000 ;
        RECT 19.200 237.600 52.000 238.400 ;
        RECT 19.200 236.800 51.200 237.600 ;
        RECT 18.400 236.000 51.200 236.800 ;
        RECT 18.400 235.200 50.400 236.000 ;
        RECT 17.600 233.600 49.600 235.200 ;
        RECT 16.800 232.800 48.800 233.600 ;
        RECT 16.800 232.000 48.000 232.800 ;
        RECT 16.000 231.200 48.000 232.000 ;
        RECT 16.000 230.400 47.200 231.200 ;
        RECT 15.200 228.800 46.400 230.400 ;
        RECT 14.400 227.200 45.600 228.800 ;
        RECT 13.600 225.600 44.800 227.200 ;
        RECT 13.600 224.800 44.000 225.600 ;
        RECT 12.800 224.000 44.000 224.800 ;
        RECT 12.800 223.200 43.200 224.000 ;
        RECT 12.000 222.400 43.200 223.200 ;
        RECT 12.000 221.600 42.400 222.400 ;
        RECT 11.200 220.800 42.400 221.600 ;
        RECT 11.200 219.200 41.600 220.800 ;
        RECT 10.400 217.600 40.800 219.200 ;
        RECT 10.400 216.800 40.000 217.600 ;
        RECT 9.600 216.000 40.000 216.800 ;
        RECT 9.600 215.200 39.200 216.000 ;
        RECT 8.800 214.400 39.200 215.200 ;
        RECT 8.800 212.800 38.400 214.400 ;
        RECT 8.000 210.400 37.600 212.800 ;
        RECT 7.200 208.000 36.800 210.400 ;
        RECT 7.200 207.200 36.000 208.000 ;
        RECT 6.400 206.400 36.000 207.200 ;
        RECT 6.400 204.800 35.200 206.400 ;
        RECT 5.600 204.000 35.200 204.800 ;
        RECT 5.600 201.600 34.400 204.000 ;
        RECT 4.800 198.400 33.600 201.600 ;
        RECT 4.000 196.000 32.800 198.400 ;
        RECT 4.000 194.400 32.000 196.000 ;
        RECT 3.200 192.800 32.000 194.400 ;
        RECT 3.200 190.400 31.200 192.800 ;
        RECT 2.400 188.800 31.200 190.400 ;
        RECT 2.400 185.600 30.400 188.800 ;
        RECT 1.600 184.800 30.400 185.600 ;
        RECT 1.600 180.000 29.600 184.800 ;
        RECT 0.800 179.200 29.600 180.000 ;
        RECT 0.800 172.000 28.800 179.200 ;
        RECT 0.800 170.400 28.000 172.000 ;
        RECT 0.000 152.800 28.000 170.400 ;
        RECT 0.800 151.200 28.000 152.800 ;
        RECT 0.800 143.200 28.800 151.200 ;
        RECT 1.600 138.400 29.600 143.200 ;
        RECT 1.600 137.600 30.400 138.400 ;
        RECT 2.400 134.400 30.400 137.600 ;
        RECT 2.400 132.800 31.200 134.400 ;
        RECT 3.200 130.400 31.200 132.800 ;
        RECT 3.200 128.000 32.000 130.400 ;
        RECT 4.000 127.200 32.000 128.000 ;
        RECT 4.000 124.800 32.800 127.200 ;
        RECT 4.800 121.600 33.600 124.800 ;
        RECT 5.600 119.200 34.400 121.600 ;
        RECT 5.600 118.400 35.200 119.200 ;
        RECT 6.400 116.800 35.200 118.400 ;
        RECT 6.400 116.000 36.000 116.800 ;
        RECT 7.200 115.200 36.000 116.000 ;
        RECT 7.200 112.800 36.800 115.200 ;
        RECT 8.000 110.400 37.600 112.800 ;
        RECT 8.800 108.800 38.400 110.400 ;
        RECT 8.800 108.000 39.200 108.800 ;
        RECT 9.600 107.200 39.200 108.000 ;
        RECT 9.600 106.400 40.000 107.200 ;
        RECT 10.400 105.600 40.000 106.400 ;
        RECT 10.400 104.000 40.800 105.600 ;
        RECT 11.200 103.200 40.800 104.000 ;
        RECT 11.200 101.600 41.600 103.200 ;
        RECT 12.000 100.000 42.400 101.600 ;
        RECT 12.800 98.400 43.200 100.000 ;
        RECT 12.800 97.600 44.000 98.400 ;
        RECT 13.600 96.000 44.800 97.600 ;
        RECT 14.400 94.400 45.600 96.000 ;
        RECT 15.200 92.800 46.400 94.400 ;
        RECT 16.000 92.000 47.200 92.800 ;
        RECT 16.000 91.200 48.000 92.000 ;
        RECT 16.800 90.400 48.000 91.200 ;
        RECT 16.800 89.600 48.800 90.400 ;
        RECT 17.600 88.000 49.600 89.600 ;
        RECT 18.400 86.400 50.400 88.000 ;
        RECT 19.200 85.600 51.200 86.400 ;
        RECT 19.200 84.800 52.000 85.600 ;
        RECT 20.000 83.200 52.800 84.800 ;
        RECT 20.800 82.400 53.600 83.200 ;
        RECT 20.800 81.600 54.400 82.400 ;
        RECT 21.600 80.800 54.400 81.600 ;
        RECT 22.400 80.000 55.200 80.800 ;
        RECT 22.400 79.200 56.000 80.000 ;
        RECT 23.200 78.400 56.800 79.200 ;
        RECT 23.200 77.600 57.600 78.400 ;
        RECT 24.000 76.800 57.600 77.600 ;
        RECT 24.800 76.000 58.400 76.800 ;
        RECT 24.800 75.200 59.200 76.000 ;
        RECT 25.600 74.400 60.000 75.200 ;
        RECT 25.600 73.600 60.800 74.400 ;
        RECT 26.400 72.800 61.600 73.600 ;
        RECT 27.200 72.000 61.600 72.800 ;
        RECT 27.200 71.200 62.400 72.000 ;
        RECT 28.000 70.400 63.200 71.200 ;
        RECT 28.800 69.600 64.000 70.400 ;
        RECT 28.800 68.800 64.800 69.600 ;
        RECT 29.600 68.000 65.600 68.800 ;
        RECT 30.400 67.200 66.400 68.000 ;
        RECT 31.200 66.400 67.200 67.200 ;
        RECT 31.200 65.600 68.000 66.400 ;
        RECT 32.000 64.800 68.800 65.600 ;
        RECT 32.800 64.000 69.600 64.800 ;
        RECT 33.600 63.200 70.400 64.000 ;
        RECT 33.600 62.400 71.200 63.200 ;
        RECT 34.400 61.600 72.000 62.400 ;
        RECT 35.200 60.800 73.600 61.600 ;
        RECT 36.000 60.000 74.400 60.800 ;
        RECT 36.000 59.200 75.200 60.000 ;
        RECT 36.800 58.400 76.000 59.200 ;
        RECT 37.600 57.600 76.800 58.400 ;
        RECT 38.400 56.800 77.600 57.600 ;
        RECT 39.200 56.000 79.200 56.800 ;
        RECT 40.000 55.200 80.000 56.000 ;
        RECT 40.800 54.400 80.800 55.200 ;
        RECT 40.800 53.600 81.600 54.400 ;
        RECT 41.600 52.800 83.200 53.600 ;
        RECT 42.400 52.000 84.000 52.800 ;
        RECT 43.200 51.200 84.800 52.000 ;
        RECT 44.000 50.400 86.400 51.200 ;
        RECT 44.800 49.600 87.200 50.400 ;
        RECT 45.600 48.800 88.800 49.600 ;
        RECT 46.400 48.000 89.600 48.800 ;
        RECT 47.200 47.200 91.200 48.000 ;
        RECT 48.000 46.400 92.000 47.200 ;
        RECT 48.800 45.600 93.600 46.400 ;
        RECT 49.600 44.800 95.200 45.600 ;
        RECT 50.400 44.000 96.800 44.800 ;
        RECT 51.200 43.200 98.400 44.000 ;
        RECT 52.000 42.400 98.400 43.200 ;
        RECT 52.800 41.600 98.400 42.400 ;
        RECT 53.600 40.800 98.400 41.600 ;
        RECT 54.400 40.000 98.400 40.800 ;
        RECT 56.000 39.200 98.400 40.000 ;
        RECT 56.800 38.400 98.400 39.200 ;
        RECT 57.600 37.600 98.400 38.400 ;
        RECT 58.400 36.800 98.400 37.600 ;
        RECT 59.200 36.000 97.600 36.800 ;
        RECT 60.800 35.200 97.600 36.000 ;
        RECT 61.600 34.400 97.600 35.200 ;
        RECT 62.400 33.600 97.600 34.400 ;
        RECT 63.200 32.800 97.600 33.600 ;
        RECT 64.800 32.000 97.600 32.800 ;
        RECT 65.600 31.200 97.600 32.000 ;
        RECT 66.400 30.400 97.600 31.200 ;
        RECT 68.000 29.600 97.600 30.400 ;
        RECT 68.800 28.800 96.800 29.600 ;
        RECT 70.400 28.000 96.800 28.800 ;
        RECT 71.200 27.200 96.800 28.000 ;
        RECT 72.000 26.400 96.800 27.200 ;
        RECT 73.600 25.600 96.800 26.400 ;
        RECT 75.200 24.800 96.800 25.600 ;
        RECT 76.000 24.000 96.800 24.800 ;
        RECT 77.600 23.200 96.800 24.000 ;
        RECT 78.400 22.400 96.000 23.200 ;
        RECT 80.000 21.600 96.000 22.400 ;
        RECT 81.600 20.800 96.000 21.600 ;
        RECT 82.400 20.000 96.000 20.800 ;
        RECT 84.000 19.200 96.000 20.000 ;
        RECT 85.600 18.400 96.000 19.200 ;
        RECT 87.200 17.600 96.000 18.400 ;
        RECT 88.800 16.800 96.000 17.600 ;
        RECT 89.600 16.000 95.200 16.800 ;
        RECT 91.200 15.200 95.200 16.000 ;
        RECT 92.800 14.400 95.200 15.200 ;
        RECT 94.400 13.600 95.200 14.400 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 313.600 468.000 315.200 468.800 ;
        RECT 312.800 467.200 315.200 468.000 ;
        RECT 312.000 465.600 315.200 467.200 ;
        RECT 311.200 464.800 316.000 465.600 ;
        RECT 310.400 464.000 316.000 464.800 ;
        RECT 309.600 463.200 316.000 464.000 ;
        RECT 308.800 462.400 316.000 463.200 ;
        RECT 308.000 460.800 316.800 462.400 ;
        RECT 307.200 460.000 316.800 460.800 ;
        RECT 306.400 459.200 317.600 460.000 ;
        RECT 305.600 458.400 317.600 459.200 ;
        RECT 304.800 456.800 317.600 458.400 ;
        RECT 304.000 456.000 318.400 456.800 ;
        RECT 303.200 455.200 318.400 456.000 ;
        RECT 302.400 454.400 318.400 455.200 ;
        RECT 301.600 453.600 318.400 454.400 ;
        RECT 300.800 452.000 319.200 453.600 ;
        RECT 300.000 451.200 319.200 452.000 ;
        RECT 299.200 450.400 319.200 451.200 ;
        RECT 298.400 449.600 320.000 450.400 ;
        RECT 297.600 448.000 320.000 449.600 ;
        RECT 296.800 447.200 320.000 448.000 ;
        RECT 296.000 446.400 320.800 447.200 ;
        RECT 295.200 445.600 320.800 446.400 ;
        RECT 294.400 444.000 320.800 445.600 ;
        RECT 293.600 443.200 321.600 444.000 ;
        RECT 292.800 442.400 321.600 443.200 ;
        RECT 292.000 441.600 321.600 442.400 ;
        RECT 291.200 440.800 321.600 441.600 ;
        RECT 291.200 440.000 322.400 440.800 ;
        RECT 290.400 439.200 322.400 440.000 ;
        RECT 289.600 438.400 322.400 439.200 ;
        RECT 288.800 437.600 322.400 438.400 ;
        RECT 288.000 436.800 322.400 437.600 ;
        RECT 288.000 436.000 323.200 436.800 ;
        RECT 287.200 435.200 323.200 436.000 ;
        RECT 286.400 434.400 323.200 435.200 ;
        RECT 285.600 433.600 323.200 434.400 ;
        RECT 284.800 432.800 323.200 433.600 ;
        RECT 284.800 432.000 324.000 432.800 ;
        RECT 284.000 431.200 324.000 432.000 ;
        RECT 283.200 430.400 324.000 431.200 ;
        RECT 282.400 429.600 324.000 430.400 ;
        RECT 281.600 428.800 324.000 429.600 ;
        RECT 281.600 428.000 324.800 428.800 ;
        RECT 280.800 427.200 324.800 428.000 ;
        RECT 280.000 426.400 324.800 427.200 ;
        RECT 279.200 425.600 324.800 426.400 ;
        RECT 278.400 424.000 324.800 425.600 ;
        RECT 277.600 423.200 324.800 424.000 ;
        RECT 276.800 422.400 325.600 423.200 ;
        RECT 276.000 421.600 325.600 422.400 ;
        RECT 275.200 420.000 325.600 421.600 ;
        RECT 274.400 419.200 325.600 420.000 ;
        RECT 273.600 418.400 325.600 419.200 ;
        RECT 272.800 416.800 325.600 418.400 ;
        RECT 272.000 416.000 325.600 416.800 ;
        RECT 271.200 415.200 325.600 416.000 ;
        RECT 270.400 414.400 325.600 415.200 ;
        RECT 269.600 412.800 325.600 414.400 ;
        RECT 268.800 412.000 326.400 412.800 ;
        RECT 268.000 411.200 326.400 412.000 ;
        RECT 267.200 409.600 326.400 411.200 ;
        RECT 266.400 408.800 326.400 409.600 ;
        RECT 265.600 408.000 325.600 408.800 ;
        RECT 264.800 406.400 325.600 408.000 ;
        RECT 264.000 405.600 325.600 406.400 ;
        RECT 263.200 404.800 325.600 405.600 ;
        RECT 262.400 404.000 325.600 404.800 ;
        RECT 261.600 402.400 325.600 404.000 ;
        RECT 260.800 401.600 325.600 402.400 ;
        RECT 260.000 400.800 325.600 401.600 ;
        RECT 259.200 399.200 325.600 400.800 ;
        RECT 258.400 398.400 324.800 399.200 ;
        RECT 257.600 397.600 324.800 398.400 ;
        RECT 256.800 396.000 324.800 397.600 ;
        RECT 256.000 395.200 324.800 396.000 ;
        RECT 255.200 394.400 324.800 395.200 ;
        RECT 254.400 392.800 324.000 394.400 ;
        RECT 253.600 392.000 324.000 392.800 ;
        RECT 252.800 391.200 324.000 392.000 ;
        RECT 252.000 389.600 324.000 391.200 ;
        RECT 251.200 388.800 323.200 389.600 ;
        RECT 250.400 388.000 323.200 388.800 ;
        RECT 249.600 386.400 323.200 388.000 ;
        RECT 248.800 385.600 322.400 386.400 ;
        RECT 248.000 384.000 322.400 385.600 ;
        RECT 247.200 383.200 322.400 384.000 ;
        RECT 246.400 382.400 321.600 383.200 ;
        RECT 245.600 380.800 321.600 382.400 ;
        RECT 244.800 380.000 321.600 380.800 ;
        RECT 244.000 379.200 320.800 380.000 ;
        RECT 243.200 377.600 320.800 379.200 ;
        RECT 242.400 376.800 320.800 377.600 ;
        RECT 241.600 375.200 320.000 376.800 ;
        RECT 240.800 374.400 320.000 375.200 ;
        RECT 240.000 373.600 319.200 374.400 ;
        RECT 239.200 372.000 319.200 373.600 ;
        RECT 238.400 371.200 318.400 372.000 ;
        RECT 237.600 369.600 318.400 371.200 ;
        RECT 236.800 368.800 318.400 369.600 ;
        RECT 236.000 368.000 317.600 368.800 ;
        RECT 235.200 366.400 317.600 368.000 ;
        RECT 234.400 365.600 316.800 366.400 ;
        RECT 233.600 364.000 316.800 365.600 ;
        RECT 232.800 363.200 316.000 364.000 ;
        RECT 232.000 361.600 316.000 363.200 ;
        RECT 231.200 360.800 315.200 361.600 ;
        RECT 230.400 359.200 315.200 360.800 ;
        RECT 229.600 358.400 314.400 359.200 ;
        RECT 228.800 357.600 314.400 358.400 ;
        RECT 228.000 356.800 314.400 357.600 ;
        RECT 228.000 356.000 313.600 356.800 ;
        RECT 227.200 355.200 313.600 356.000 ;
        RECT 226.400 354.400 313.600 355.200 ;
        RECT 226.400 353.600 312.800 354.400 ;
        RECT 225.600 352.800 312.800 353.600 ;
        RECT 224.800 352.000 312.800 352.800 ;
        RECT 224.800 351.200 312.000 352.000 ;
        RECT 224.000 350.400 312.000 351.200 ;
        RECT 223.200 349.600 312.000 350.400 ;
        RECT 223.200 348.800 311.200 349.600 ;
        RECT 222.400 348.000 311.200 348.800 ;
        RECT 221.600 347.200 311.200 348.000 ;
        RECT 221.600 346.400 310.400 347.200 ;
        RECT 220.800 345.600 310.400 346.400 ;
        RECT 220.000 344.000 309.600 345.600 ;
        RECT 219.200 343.200 309.600 344.000 ;
        RECT 218.400 341.600 308.800 343.200 ;
        RECT 217.600 340.800 308.800 341.600 ;
        RECT 217.600 340.000 308.000 340.800 ;
        RECT 216.800 339.200 308.000 340.000 ;
        RECT 216.000 337.600 307.200 339.200 ;
        RECT 215.200 336.800 307.200 337.600 ;
        RECT 214.400 335.200 306.400 336.800 ;
        RECT 213.600 334.400 306.400 335.200 ;
        RECT 212.800 332.800 305.600 334.400 ;
        RECT 212.000 331.200 304.800 332.800 ;
        RECT 211.200 330.400 304.800 331.200 ;
        RECT 210.400 328.800 304.000 330.400 ;
        RECT 209.600 328.000 304.000 328.800 ;
        RECT 208.800 326.400 303.200 328.000 ;
        RECT 208.000 324.800 302.400 326.400 ;
        RECT 207.200 324.000 302.400 324.800 ;
        RECT 206.400 322.400 301.600 324.000 ;
        RECT 205.600 320.800 300.800 322.400 ;
        RECT 204.800 320.000 300.800 320.800 ;
        RECT 204.000 318.400 300.000 320.000 ;
        RECT 203.200 316.800 299.200 318.400 ;
        RECT 202.400 316.000 299.200 316.800 ;
        RECT 201.600 314.400 298.400 316.000 ;
        RECT 200.800 312.800 297.600 314.400 ;
        RECT 200.000 312.000 297.600 312.800 ;
        RECT 199.200 310.400 296.800 312.000 ;
        RECT 198.400 308.800 296.000 310.400 ;
        RECT 197.600 308.000 296.000 308.800 ;
        RECT 197.600 307.200 295.200 308.000 ;
        RECT 196.800 306.400 295.200 307.200 ;
        RECT 196.800 305.600 294.400 306.400 ;
        RECT 196.000 304.800 294.400 305.600 ;
        RECT 195.200 304.000 294.400 304.800 ;
        RECT 195.200 303.200 293.600 304.000 ;
        RECT 194.400 302.400 293.600 303.200 ;
        RECT 194.400 301.600 292.800 302.400 ;
        RECT 193.600 300.800 292.800 301.600 ;
        RECT 193.600 300.000 292.000 300.800 ;
        RECT 192.800 298.400 292.000 300.000 ;
        RECT 192.000 297.600 291.200 298.400 ;
        RECT 191.200 296.800 291.200 297.600 ;
        RECT 191.200 296.000 290.400 296.800 ;
        RECT 190.400 294.400 290.400 296.000 ;
        RECT 189.600 292.800 289.600 294.400 ;
        RECT 188.800 291.200 288.800 292.800 ;
        RECT 188.000 289.600 288.000 291.200 ;
        RECT 187.200 288.800 288.000 289.600 ;
        RECT 187.200 288.000 287.200 288.800 ;
        RECT 186.400 287.200 287.200 288.000 ;
        RECT 186.400 286.400 286.400 287.200 ;
        RECT 185.600 284.800 286.400 286.400 ;
        RECT 184.800 283.200 285.600 284.800 ;
        RECT 184.000 281.600 284.800 283.200 ;
        RECT 183.200 280.000 284.000 281.600 ;
        RECT 182.400 279.200 284.000 280.000 ;
        RECT 182.400 278.400 283.200 279.200 ;
        RECT 181.600 277.600 283.200 278.400 ;
        RECT 181.600 276.800 282.400 277.600 ;
        RECT 180.800 276.000 282.400 276.800 ;
        RECT 180.800 275.200 281.600 276.000 ;
        RECT 180.000 273.600 281.600 275.200 ;
        RECT 179.200 272.000 280.800 273.600 ;
        RECT 178.400 270.400 280.000 272.000 ;
        RECT 177.600 268.800 279.200 270.400 ;
        RECT 176.800 268.000 279.200 268.800 ;
        RECT 176.800 267.200 278.400 268.000 ;
        RECT 176.000 266.400 278.400 267.200 ;
        RECT 176.000 264.800 277.600 266.400 ;
        RECT 175.200 263.200 276.800 264.800 ;
        RECT 174.400 262.400 276.800 263.200 ;
        RECT 174.400 261.600 276.000 262.400 ;
        RECT 173.600 260.800 276.000 261.600 ;
        RECT 173.600 260.000 275.200 260.800 ;
        RECT 172.800 259.200 275.200 260.000 ;
        RECT 172.800 257.600 274.400 259.200 ;
        RECT 172.000 256.800 273.600 257.600 ;
        RECT 172.000 256.000 272.800 256.800 ;
        RECT 171.200 255.200 272.000 256.000 ;
        RECT 171.200 254.400 271.200 255.200 ;
        RECT 170.400 253.600 270.400 254.400 ;
        RECT 170.400 252.800 269.600 253.600 ;
        RECT 169.600 252.000 268.800 252.800 ;
        RECT 169.600 251.200 268.000 252.000 ;
        RECT 169.600 250.400 267.200 251.200 ;
        RECT 168.800 249.600 266.400 250.400 ;
        RECT 168.800 248.800 265.600 249.600 ;
        RECT 168.000 248.000 264.800 248.800 ;
        RECT 168.000 247.200 264.000 248.000 ;
        RECT 168.000 246.400 263.200 247.200 ;
        RECT 167.200 245.600 262.400 246.400 ;
        RECT 167.200 244.800 261.600 245.600 ;
        RECT 166.400 244.000 260.800 244.800 ;
        RECT 166.400 243.200 260.000 244.000 ;
        RECT 165.600 242.400 259.200 243.200 ;
        RECT 165.600 241.600 258.400 242.400 ;
        RECT 165.600 240.800 257.600 241.600 ;
        RECT 164.800 239.200 256.800 240.800 ;
        RECT 164.000 238.400 256.000 239.200 ;
        RECT 164.000 237.600 255.200 238.400 ;
        RECT 164.000 236.800 254.400 237.600 ;
        RECT 163.200 236.000 253.600 236.800 ;
        RECT 163.200 235.200 252.800 236.000 ;
        RECT 162.400 234.400 252.000 235.200 ;
        RECT 162.400 233.600 251.200 234.400 ;
        RECT 162.400 232.800 250.400 233.600 ;
        RECT 161.600 232.000 249.600 232.800 ;
        RECT 161.600 231.200 248.800 232.000 ;
        RECT 160.800 230.400 248.000 231.200 ;
        RECT 160.800 229.600 247.200 230.400 ;
        RECT 160.800 228.800 246.400 229.600 ;
        RECT 160.000 228.000 245.600 228.800 ;
        RECT 160.000 227.200 244.800 228.000 ;
        RECT 159.200 226.400 244.000 227.200 ;
        RECT 159.200 225.600 243.200 226.400 ;
        RECT 159.200 224.800 242.400 225.600 ;
        RECT 158.400 224.000 241.600 224.800 ;
        RECT 158.400 223.200 240.800 224.000 ;
        RECT 158.400 222.400 240.000 223.200 ;
        RECT 157.600 221.600 239.200 222.400 ;
        RECT 157.600 220.800 238.400 221.600 ;
        RECT 156.800 220.000 237.600 220.800 ;
        RECT 156.800 219.200 236.800 220.000 ;
        RECT 156.800 218.400 236.000 219.200 ;
        RECT 156.000 217.600 235.200 218.400 ;
        RECT 156.000 216.800 234.400 217.600 ;
        RECT 156.000 216.000 233.600 216.800 ;
        RECT 155.200 215.200 233.600 216.000 ;
        RECT 155.200 214.400 232.800 215.200 ;
        RECT 154.400 213.600 232.000 214.400 ;
        RECT 154.400 212.800 231.200 213.600 ;
        RECT 154.400 212.000 230.400 212.800 ;
        RECT 153.600 211.200 229.600 212.000 ;
        RECT 153.600 210.400 228.800 211.200 ;
        RECT 153.600 209.600 228.000 210.400 ;
        RECT 152.800 208.800 227.200 209.600 ;
        RECT 152.800 208.000 226.400 208.800 ;
        RECT 152.800 207.200 225.600 208.000 ;
        RECT 152.000 206.400 224.800 207.200 ;
        RECT 152.000 205.600 224.000 206.400 ;
        RECT 151.200 204.000 223.200 205.600 ;
        RECT 151.200 203.200 222.400 204.000 ;
        RECT 150.400 202.400 221.600 203.200 ;
        RECT 150.400 201.600 220.800 202.400 ;
        RECT 150.400 200.800 220.000 201.600 ;
        RECT 149.600 200.000 219.200 200.800 ;
        RECT 149.600 199.200 218.400 200.000 ;
        RECT 149.600 198.400 217.600 199.200 ;
        RECT 148.800 197.600 217.600 198.400 ;
        RECT 148.800 196.800 216.800 197.600 ;
        RECT 148.800 196.000 216.000 196.800 ;
        RECT 148.000 195.200 215.200 196.000 ;
        RECT 148.000 194.400 214.400 195.200 ;
        RECT 148.000 193.600 213.600 194.400 ;
        RECT 147.200 192.000 212.800 193.600 ;
        RECT 147.200 191.200 212.000 192.000 ;
        RECT 146.400 190.400 211.200 191.200 ;
        RECT 146.400 189.600 210.400 190.400 ;
        RECT 146.400 188.800 209.600 189.600 ;
        RECT 145.600 187.200 208.800 188.800 ;
        RECT 145.600 186.400 208.000 187.200 ;
        RECT 144.800 185.600 207.200 186.400 ;
        RECT 144.800 184.800 206.400 185.600 ;
        RECT 144.800 184.000 205.600 184.800 ;
        RECT 144.000 182.400 204.800 184.000 ;
        RECT 144.000 181.600 204.000 182.400 ;
        RECT 143.200 180.800 203.200 181.600 ;
        RECT 143.200 180.000 202.400 180.800 ;
        RECT 143.200 178.400 201.600 180.000 ;
        RECT 142.400 177.600 200.800 178.400 ;
        RECT 142.400 176.800 200.000 177.600 ;
        RECT 142.400 176.000 199.200 176.800 ;
        RECT 141.600 175.200 199.200 176.000 ;
        RECT 141.600 174.400 198.400 175.200 ;
        RECT 141.600 173.600 197.600 174.400 ;
        RECT 140.800 172.800 196.800 173.600 ;
        RECT 140.800 171.200 196.000 172.800 ;
        RECT 140.000 170.400 195.200 171.200 ;
        RECT 140.000 169.600 194.400 170.400 ;
        RECT 140.000 168.800 193.600 169.600 ;
        RECT 139.200 168.000 193.600 168.800 ;
        RECT 139.200 167.200 192.800 168.000 ;
        RECT 139.200 166.400 192.000 167.200 ;
        RECT 139.200 165.600 191.200 166.400 ;
        RECT 138.400 164.800 191.200 165.600 ;
        RECT 138.400 164.000 190.400 164.800 ;
        RECT 138.400 163.200 189.600 164.000 ;
        RECT 137.600 161.600 188.800 163.200 ;
        RECT 137.600 160.800 188.000 161.600 ;
        RECT 136.800 160.000 187.200 160.800 ;
        RECT 136.800 158.400 186.400 160.000 ;
        RECT 136.800 157.600 185.600 158.400 ;
        RECT 136.000 156.000 184.800 157.600 ;
        RECT 136.000 155.200 184.000 156.000 ;
        RECT 135.200 154.400 183.200 155.200 ;
        RECT 135.200 152.800 182.400 154.400 ;
        RECT 135.200 152.000 181.600 152.800 ;
        RECT 134.400 151.200 180.800 152.000 ;
        RECT 134.400 149.600 180.000 151.200 ;
        RECT 133.600 148.800 179.200 149.600 ;
        RECT 133.600 147.200 178.400 148.800 ;
        RECT 132.800 146.400 177.600 147.200 ;
        RECT 132.800 145.600 176.800 146.400 ;
        RECT 132.800 144.000 176.000 145.600 ;
        RECT 132.000 143.200 175.200 144.000 ;
        RECT 132.000 142.400 174.400 143.200 ;
        RECT 132.000 141.600 173.600 142.400 ;
        RECT 131.200 140.800 173.600 141.600 ;
        RECT 131.200 140.000 172.800 140.800 ;
        RECT 131.200 138.400 172.000 140.000 ;
        RECT 130.400 137.600 171.200 138.400 ;
        RECT 130.400 136.000 170.400 137.600 ;
        RECT 129.600 135.200 169.600 136.000 ;
        RECT 129.600 134.400 168.800 135.200 ;
        RECT 129.600 132.800 168.000 134.400 ;
        RECT 128.800 132.000 167.200 132.800 ;
        RECT 128.800 130.400 166.400 132.000 ;
        RECT 128.000 129.600 165.600 130.400 ;
        RECT 128.000 128.000 164.800 129.600 ;
        RECT 128.000 127.200 164.000 128.000 ;
        RECT 127.200 125.600 163.200 127.200 ;
        RECT 127.200 124.800 162.400 125.600 ;
        RECT 126.400 123.200 161.600 124.800 ;
        RECT 126.400 122.400 160.800 123.200 ;
        RECT 126.400 121.600 160.000 122.400 ;
        RECT 125.600 120.800 160.000 121.600 ;
        RECT 125.600 120.000 159.200 120.800 ;
        RECT 125.600 119.200 158.400 120.000 ;
        RECT 124.800 118.400 158.400 119.200 ;
        RECT 124.800 117.600 157.600 118.400 ;
        RECT 124.800 116.000 156.800 117.600 ;
        RECT 124.000 115.200 156.000 116.000 ;
        RECT 124.000 113.600 155.200 115.200 ;
        RECT 123.200 112.800 154.400 113.600 ;
        RECT 123.200 111.200 153.600 112.800 ;
        RECT 123.200 110.400 152.800 111.200 ;
        RECT 122.400 108.800 152.000 110.400 ;
        RECT 122.400 108.000 151.200 108.800 ;
        RECT 122.400 107.200 150.400 108.000 ;
        RECT 121.600 106.400 150.400 107.200 ;
        RECT 121.600 104.800 149.600 106.400 ;
        RECT 121.600 104.000 148.800 104.800 ;
        RECT 120.800 102.400 148.000 104.000 ;
        RECT 120.800 101.600 147.200 102.400 ;
        RECT 120.000 100.800 147.200 101.600 ;
        RECT 120.000 100.000 146.400 100.800 ;
        RECT 120.000 98.400 145.600 100.000 ;
        RECT 119.200 97.600 144.800 98.400 ;
        RECT 119.200 96.000 144.000 97.600 ;
        RECT 119.200 95.200 143.200 96.000 ;
        RECT 118.400 94.400 143.200 95.200 ;
        RECT 118.400 92.800 142.400 94.400 ;
        RECT 118.400 92.000 141.600 92.800 ;
        RECT 117.600 90.400 140.800 92.000 ;
        RECT 117.600 88.800 140.000 90.400 ;
        RECT 116.800 87.200 139.200 88.800 ;
        RECT 116.800 86.400 138.400 87.200 ;
        RECT 116.800 85.600 137.600 86.400 ;
        RECT 116.000 84.800 137.600 85.600 ;
        RECT 116.000 83.200 136.800 84.800 ;
        RECT 116.000 82.400 136.000 83.200 ;
        RECT 115.200 81.600 136.000 82.400 ;
        RECT 115.200 80.000 135.200 81.600 ;
        RECT 115.200 78.400 134.400 80.000 ;
        RECT 114.400 77.600 133.600 78.400 ;
        RECT 114.400 76.000 132.800 77.600 ;
        RECT 114.400 75.200 132.000 76.000 ;
        RECT 113.600 74.400 132.000 75.200 ;
        RECT 113.600 72.800 131.200 74.400 ;
        RECT 113.600 71.200 130.400 72.800 ;
        RECT 112.800 69.600 129.600 71.200 ;
        RECT 112.800 68.000 128.800 69.600 ;
        RECT 112.000 66.400 128.000 68.000 ;
        RECT 112.000 64.800 127.200 66.400 ;
        RECT 112.000 64.000 126.400 64.800 ;
        RECT 111.200 63.200 126.400 64.000 ;
        RECT 111.200 61.600 125.600 63.200 ;
        RECT 111.200 60.000 124.800 61.600 ;
        RECT 110.400 58.400 124.000 60.000 ;
        RECT 110.400 56.800 123.200 58.400 ;
        RECT 110.400 56.000 122.400 56.800 ;
        RECT 109.600 55.200 122.400 56.000 ;
        RECT 109.600 53.600 121.600 55.200 ;
        RECT 109.600 52.800 120.800 53.600 ;
        RECT 108.800 52.000 120.800 52.800 ;
        RECT 108.800 50.400 120.000 52.000 ;
        RECT 108.800 48.800 119.200 50.400 ;
        RECT 108.000 47.200 118.400 48.800 ;
        RECT 108.000 45.600 117.600 47.200 ;
        RECT 108.000 44.000 116.800 45.600 ;
        RECT 107.200 42.400 116.000 44.000 ;
        RECT 107.200 40.800 115.200 42.400 ;
        RECT 107.200 40.000 114.400 40.800 ;
        RECT 106.400 39.200 114.400 40.000 ;
        RECT 106.400 37.600 113.600 39.200 ;
        RECT 106.400 36.000 112.800 37.600 ;
        RECT 105.600 34.400 112.000 36.000 ;
        RECT 105.600 32.800 111.200 34.400 ;
        RECT 105.600 32.000 110.400 32.800 ;
        RECT 104.800 31.200 110.400 32.000 ;
        RECT 104.800 29.600 109.600 31.200 ;
        RECT 104.800 28.000 108.800 29.600 ;
        RECT 104.000 27.200 108.800 28.000 ;
        RECT 104.000 25.600 108.000 27.200 ;
        RECT 104.000 24.000 107.200 25.600 ;
        RECT 104.000 23.200 106.400 24.000 ;
        RECT 103.200 22.400 106.400 23.200 ;
        RECT 103.200 20.800 105.600 22.400 ;
        RECT 103.200 19.200 104.800 20.800 ;
        RECT 102.400 17.600 104.000 19.200 ;
        RECT 102.400 16.000 103.200 17.600 ;
    END
  END vdd
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 400.000 469.600 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 400.000 469.600 ;
      LAYER Metal4 ;
        RECT 389.600 334.400 390.400 335.200 ;
        RECT 388.800 333.600 390.400 334.400 ;
        RECT 387.200 332.800 390.400 333.600 ;
        RECT 386.400 332.000 390.400 332.800 ;
        RECT 384.800 331.200 390.400 332.000 ;
        RECT 384.000 330.400 390.400 331.200 ;
        RECT 382.400 329.600 390.400 330.400 ;
        RECT 381.600 328.800 390.400 329.600 ;
        RECT 380.000 328.000 390.400 328.800 ;
        RECT 378.400 327.200 390.400 328.000 ;
        RECT 377.600 326.400 390.400 327.200 ;
        RECT 376.000 325.600 390.400 326.400 ;
        RECT 375.200 324.800 390.400 325.600 ;
        RECT 373.600 324.000 390.400 324.800 ;
        RECT 372.800 323.200 390.400 324.000 ;
        RECT 371.200 322.400 390.400 323.200 ;
        RECT 370.400 321.600 390.400 322.400 ;
        RECT 368.800 320.800 390.400 321.600 ;
        RECT 368.000 320.000 390.400 320.800 ;
        RECT 366.400 319.200 390.400 320.000 ;
        RECT 365.600 318.400 390.400 319.200 ;
        RECT 364.000 317.600 390.400 318.400 ;
        RECT 363.200 316.800 390.400 317.600 ;
        RECT 361.600 316.000 390.400 316.800 ;
        RECT 360.800 315.200 390.400 316.000 ;
        RECT 360.000 314.400 390.400 315.200 ;
        RECT 358.400 313.600 390.400 314.400 ;
        RECT 357.600 312.800 390.400 313.600 ;
        RECT 356.000 312.000 390.400 312.800 ;
        RECT 355.200 311.200 390.400 312.000 ;
        RECT 353.600 310.400 390.400 311.200 ;
        RECT 352.800 309.600 390.400 310.400 ;
        RECT 352.000 308.800 390.400 309.600 ;
        RECT 350.400 308.000 390.400 308.800 ;
        RECT 349.600 307.200 390.400 308.000 ;
        RECT 348.000 306.400 390.400 307.200 ;
        RECT 347.200 305.600 390.400 306.400 ;
        RECT 346.400 304.800 390.400 305.600 ;
        RECT 344.800 304.000 390.400 304.800 ;
        RECT 344.000 303.200 390.400 304.000 ;
        RECT 343.200 302.400 390.400 303.200 ;
        RECT 341.600 301.600 389.600 302.400 ;
        RECT 340.800 300.800 389.600 301.600 ;
        RECT 340.000 300.000 389.600 300.800 ;
        RECT 338.400 299.200 389.600 300.000 ;
        RECT 337.600 298.400 389.600 299.200 ;
        RECT 336.800 297.600 389.600 298.400 ;
        RECT 335.200 296.800 389.600 297.600 ;
        RECT 334.400 296.000 389.600 296.800 ;
        RECT 333.600 295.200 388.800 296.000 ;
        RECT 332.000 294.400 388.800 295.200 ;
        RECT 331.200 293.600 388.800 294.400 ;
        RECT 330.400 292.800 388.800 293.600 ;
        RECT 328.800 292.000 388.800 292.800 ;
        RECT 328.000 291.200 388.000 292.000 ;
        RECT 327.200 290.400 388.000 291.200 ;
        RECT 326.400 289.600 388.000 290.400 ;
        RECT 324.800 288.800 388.000 289.600 ;
        RECT 324.000 288.000 387.200 288.800 ;
        RECT 323.200 287.200 387.200 288.000 ;
        RECT 321.600 286.400 387.200 287.200 ;
        RECT 320.800 285.600 387.200 286.400 ;
        RECT 320.000 284.800 386.400 285.600 ;
        RECT 319.200 284.000 386.400 284.800 ;
        RECT 318.400 283.200 386.400 284.000 ;
        RECT 316.800 282.400 386.400 283.200 ;
        RECT 316.000 281.600 385.600 282.400 ;
        RECT 315.200 280.800 385.600 281.600 ;
        RECT 314.400 280.000 384.800 280.800 ;
        RECT 312.800 279.200 384.800 280.000 ;
        RECT 312.000 278.400 384.000 279.200 ;
        RECT 311.200 277.600 384.000 278.400 ;
        RECT 310.400 276.800 384.000 277.600 ;
        RECT 308.800 276.000 383.200 276.800 ;
        RECT 308.000 275.200 383.200 276.000 ;
        RECT 307.200 274.400 382.400 275.200 ;
        RECT 306.400 273.600 382.400 274.400 ;
        RECT 305.600 272.800 381.600 273.600 ;
        RECT 304.000 272.000 381.600 272.800 ;
        RECT 303.200 271.200 381.600 272.000 ;
        RECT 302.400 270.400 380.800 271.200 ;
        RECT 301.600 269.600 380.800 270.400 ;
        RECT 300.800 268.800 380.000 269.600 ;
        RECT 300.000 268.000 379.200 268.800 ;
        RECT 298.400 267.200 379.200 268.000 ;
        RECT 297.600 266.400 378.400 267.200 ;
        RECT 296.800 265.600 378.400 266.400 ;
        RECT 296.000 264.800 377.600 265.600 ;
        RECT 295.200 264.000 376.800 264.800 ;
        RECT 293.600 263.200 376.800 264.000 ;
        RECT 292.800 262.400 376.000 263.200 ;
        RECT 292.000 261.600 376.000 262.400 ;
        RECT 291.200 260.800 375.200 261.600 ;
        RECT 290.400 260.000 374.400 260.800 ;
        RECT 289.600 259.200 374.400 260.000 ;
        RECT 288.800 258.400 373.600 259.200 ;
        RECT 288.000 257.600 373.600 258.400 ;
        RECT 286.400 256.800 372.800 257.600 ;
        RECT 285.600 256.000 372.000 256.800 ;
        RECT 284.800 255.200 372.000 256.000 ;
        RECT 284.000 254.400 371.200 255.200 ;
        RECT 283.200 253.600 370.400 254.400 ;
        RECT 282.400 252.800 370.400 253.600 ;
        RECT 281.600 252.000 369.600 252.800 ;
        RECT 280.800 251.200 368.800 252.000 ;
        RECT 279.200 250.400 368.000 251.200 ;
        RECT 278.400 249.600 368.000 250.400 ;
        RECT 277.600 248.800 367.200 249.600 ;
        RECT 276.800 248.000 366.400 248.800 ;
        RECT 276.000 247.200 366.400 248.000 ;
        RECT 275.200 246.400 365.600 247.200 ;
        RECT 274.400 245.600 364.800 246.400 ;
        RECT 273.600 244.800 364.000 245.600 ;
        RECT 272.800 244.000 364.000 244.800 ;
        RECT 272.000 243.200 363.200 244.000 ;
        RECT 271.200 242.400 362.400 243.200 ;
        RECT 269.600 241.600 362.400 242.400 ;
        RECT 268.800 240.800 361.600 241.600 ;
        RECT 268.000 240.000 360.800 240.800 ;
        RECT 267.200 239.200 360.000 240.000 ;
        RECT 266.400 238.400 359.200 239.200 ;
        RECT 265.600 237.600 359.200 238.400 ;
        RECT 264.800 236.800 358.400 237.600 ;
        RECT 264.000 236.000 357.600 236.800 ;
        RECT 263.200 235.200 356.800 236.000 ;
        RECT 262.400 234.400 356.800 235.200 ;
        RECT 261.600 233.600 356.000 234.400 ;
        RECT 260.800 232.800 355.200 233.600 ;
        RECT 260.000 232.000 354.400 232.800 ;
        RECT 259.200 231.200 353.600 232.000 ;
        RECT 258.400 230.400 353.600 231.200 ;
        RECT 257.600 229.600 352.800 230.400 ;
        RECT 256.800 228.800 352.000 229.600 ;
        RECT 256.000 228.000 351.200 228.800 ;
        RECT 254.400 227.200 351.200 228.000 ;
        RECT 253.600 226.400 350.400 227.200 ;
        RECT 252.800 225.600 349.600 226.400 ;
        RECT 252.000 224.800 348.800 225.600 ;
        RECT 251.200 224.000 348.000 224.800 ;
        RECT 250.400 223.200 348.000 224.000 ;
        RECT 249.600 222.400 347.200 223.200 ;
        RECT 248.800 221.600 346.400 222.400 ;
        RECT 248.000 220.800 345.600 221.600 ;
        RECT 247.200 220.000 344.800 220.800 ;
        RECT 246.400 219.200 344.800 220.000 ;
        RECT 245.600 218.400 344.000 219.200 ;
        RECT 244.800 217.600 343.200 218.400 ;
        RECT 244.000 216.800 342.400 217.600 ;
        RECT 243.200 216.000 341.600 216.800 ;
        RECT 242.400 215.200 341.600 216.000 ;
        RECT 241.600 214.400 340.800 215.200 ;
        RECT 240.800 213.600 340.000 214.400 ;
        RECT 240.000 212.800 339.200 213.600 ;
        RECT 239.200 212.000 338.400 212.800 ;
        RECT 238.400 211.200 337.600 212.000 ;
        RECT 237.600 210.400 337.600 211.200 ;
        RECT 236.800 209.600 336.800 210.400 ;
        RECT 236.000 208.800 336.000 209.600 ;
        RECT 235.200 208.000 335.200 208.800 ;
        RECT 234.400 207.200 334.400 208.000 ;
        RECT 233.600 206.400 334.400 207.200 ;
        RECT 232.800 205.600 333.600 206.400 ;
        RECT 232.000 204.800 332.800 205.600 ;
        RECT 231.200 204.000 332.000 204.800 ;
        RECT 231.200 203.200 331.200 204.000 ;
        RECT 230.400 202.400 331.200 203.200 ;
        RECT 229.600 201.600 330.400 202.400 ;
        RECT 228.800 200.800 329.600 201.600 ;
        RECT 228.000 200.000 328.800 200.800 ;
        RECT 227.200 199.200 328.000 200.000 ;
        RECT 226.400 198.400 328.000 199.200 ;
        RECT 225.600 197.600 327.200 198.400 ;
        RECT 224.800 196.800 326.400 197.600 ;
        RECT 224.000 196.000 325.600 196.800 ;
        RECT 223.200 195.200 324.800 196.000 ;
        RECT 222.400 194.400 324.000 195.200 ;
        RECT 221.600 193.600 324.000 194.400 ;
        RECT 220.800 192.800 323.200 193.600 ;
        RECT 220.000 192.000 322.400 192.800 ;
        RECT 220.000 191.200 321.600 192.000 ;
        RECT 219.200 190.400 320.800 191.200 ;
        RECT 218.400 189.600 320.800 190.400 ;
        RECT 217.600 188.800 320.000 189.600 ;
        RECT 216.800 188.000 319.200 188.800 ;
        RECT 216.000 187.200 318.400 188.000 ;
        RECT 215.200 186.400 317.600 187.200 ;
        RECT 214.400 185.600 317.600 186.400 ;
        RECT 213.600 184.800 316.800 185.600 ;
        RECT 213.600 184.000 316.000 184.800 ;
        RECT 212.800 183.200 315.200 184.000 ;
        RECT 212.000 182.400 314.400 183.200 ;
        RECT 211.200 181.600 313.600 182.400 ;
        RECT 210.400 180.800 313.600 181.600 ;
        RECT 321.600 180.800 322.400 181.600 ;
        RECT 209.600 180.000 312.800 180.800 ;
        RECT 320.800 180.000 322.400 180.800 ;
        RECT 209.600 179.200 312.000 180.000 ;
        RECT 320.000 179.200 323.200 180.000 ;
        RECT 208.800 178.400 311.200 179.200 ;
        RECT 319.200 178.400 323.200 179.200 ;
        RECT 208.000 177.600 310.400 178.400 ;
        RECT 318.400 177.600 323.200 178.400 ;
        RECT 207.200 176.800 310.400 177.600 ;
        RECT 206.400 176.000 309.600 176.800 ;
        RECT 317.600 176.000 323.200 177.600 ;
        RECT 205.600 175.200 308.800 176.000 ;
        RECT 316.800 175.200 323.200 176.000 ;
        RECT 205.600 174.400 308.000 175.200 ;
        RECT 316.000 174.400 324.000 175.200 ;
        RECT 204.800 173.600 307.200 174.400 ;
        RECT 315.200 173.600 324.000 174.400 ;
        RECT 204.000 172.800 306.400 173.600 ;
        RECT 314.400 172.800 324.000 173.600 ;
        RECT 203.200 172.000 306.400 172.800 ;
        RECT 313.600 172.000 324.000 172.800 ;
        RECT 202.400 171.200 305.600 172.000 ;
        RECT 202.400 170.400 304.800 171.200 ;
        RECT 312.800 170.400 324.000 172.000 ;
        RECT 201.600 169.600 304.000 170.400 ;
        RECT 312.000 169.600 324.000 170.400 ;
        RECT 200.800 168.800 303.200 169.600 ;
        RECT 311.200 168.800 324.000 169.600 ;
        RECT 200.000 168.000 303.200 168.800 ;
        RECT 310.400 168.000 324.000 168.800 ;
        RECT 200.000 167.200 302.400 168.000 ;
        RECT 309.600 167.200 324.000 168.000 ;
        RECT 199.200 166.400 301.600 167.200 ;
        RECT 308.800 166.400 324.000 167.200 ;
        RECT 198.400 165.600 300.800 166.400 ;
        RECT 308.000 165.600 324.000 166.400 ;
        RECT 197.600 164.800 300.000 165.600 ;
        RECT 196.800 164.000 300.000 164.800 ;
        RECT 307.200 164.000 324.000 165.600 ;
        RECT 196.800 163.200 299.200 164.000 ;
        RECT 306.400 163.200 324.000 164.000 ;
        RECT 196.000 162.400 298.400 163.200 ;
        RECT 305.600 162.400 324.000 163.200 ;
        RECT 195.200 161.600 297.600 162.400 ;
        RECT 304.800 161.600 324.000 162.400 ;
        RECT 194.400 160.800 296.800 161.600 ;
        RECT 304.000 160.800 324.000 161.600 ;
        RECT 194.400 160.000 296.000 160.800 ;
        RECT 303.200 160.000 324.000 160.800 ;
        RECT 193.600 159.200 296.000 160.000 ;
        RECT 302.400 159.200 324.000 160.000 ;
        RECT 396.800 159.200 400.000 160.000 ;
        RECT 192.800 158.400 295.200 159.200 ;
        RECT 192.800 157.600 294.400 158.400 ;
        RECT 301.600 157.600 324.000 159.200 ;
        RECT 393.600 158.400 399.200 159.200 ;
        RECT 390.400 157.600 399.200 158.400 ;
        RECT 192.000 156.800 293.600 157.600 ;
        RECT 300.800 156.800 324.000 157.600 ;
        RECT 387.200 156.800 398.400 157.600 ;
        RECT 191.200 156.000 292.800 156.800 ;
        RECT 300.000 156.000 324.000 156.800 ;
        RECT 383.200 156.000 398.400 156.800 ;
        RECT 190.400 155.200 292.800 156.000 ;
        RECT 299.200 155.200 324.000 156.000 ;
        RECT 380.000 155.200 398.400 156.000 ;
        RECT 190.400 154.400 292.000 155.200 ;
        RECT 298.400 154.400 324.000 155.200 ;
        RECT 376.800 154.400 397.600 155.200 ;
        RECT 189.600 153.600 291.200 154.400 ;
        RECT 297.600 153.600 324.000 154.400 ;
        RECT 373.600 153.600 397.600 154.400 ;
        RECT 188.800 152.800 290.400 153.600 ;
        RECT 296.800 152.800 324.000 153.600 ;
        RECT 370.400 152.800 396.800 153.600 ;
        RECT 188.000 152.000 289.600 152.800 ;
        RECT 296.800 152.000 323.200 152.800 ;
        RECT 367.200 152.000 396.800 152.800 ;
        RECT 188.000 151.200 288.800 152.000 ;
        RECT 296.000 151.200 323.200 152.000 ;
        RECT 364.000 151.200 396.800 152.000 ;
        RECT 187.200 150.400 288.800 151.200 ;
        RECT 295.200 150.400 323.200 151.200 ;
        RECT 360.800 150.400 396.000 151.200 ;
        RECT 186.400 149.600 288.000 150.400 ;
        RECT 294.400 149.600 323.200 150.400 ;
        RECT 357.600 149.600 396.000 150.400 ;
        RECT 186.400 148.800 287.200 149.600 ;
        RECT 294.400 148.800 321.600 149.600 ;
        RECT 354.400 148.800 395.200 149.600 ;
        RECT 185.600 148.000 286.400 148.800 ;
        RECT 294.400 148.000 319.200 148.800 ;
        RECT 351.200 148.000 395.200 148.800 ;
        RECT 184.800 146.400 285.600 148.000 ;
        RECT 294.400 147.200 317.600 148.000 ;
        RECT 348.000 147.200 394.400 148.000 ;
        RECT 294.400 146.400 315.200 147.200 ;
        RECT 345.600 146.400 394.400 147.200 ;
        RECT 184.000 145.600 284.800 146.400 ;
        RECT 294.400 145.600 312.800 146.400 ;
        RECT 342.400 145.600 393.600 146.400 ;
        RECT 183.200 144.800 284.000 145.600 ;
        RECT 294.400 144.800 311.200 145.600 ;
        RECT 339.200 144.800 393.600 145.600 ;
        RECT 182.400 144.000 283.200 144.800 ;
        RECT 294.400 144.000 308.800 144.800 ;
        RECT 336.000 144.000 392.800 144.800 ;
        RECT 182.400 143.200 282.400 144.000 ;
        RECT 294.400 143.200 306.400 144.000 ;
        RECT 333.600 143.200 392.800 144.000 ;
        RECT 181.600 142.400 281.600 143.200 ;
        RECT 180.800 141.600 281.600 142.400 ;
        RECT 294.400 142.400 304.000 143.200 ;
        RECT 330.400 142.400 392.000 143.200 ;
        RECT 294.400 141.600 302.400 142.400 ;
        RECT 327.200 141.600 392.000 142.400 ;
        RECT 180.800 140.800 280.800 141.600 ;
        RECT 294.400 140.800 300.000 141.600 ;
        RECT 324.800 140.800 391.200 141.600 ;
        RECT 180.000 140.000 280.000 140.800 ;
        RECT 294.400 140.000 297.600 140.800 ;
        RECT 321.600 140.000 391.200 140.800 ;
        RECT 179.200 139.200 279.200 140.000 ;
        RECT 293.600 139.200 295.200 140.000 ;
        RECT 319.200 139.200 390.400 140.000 ;
        RECT 179.200 138.400 278.400 139.200 ;
        RECT 316.000 138.400 389.600 139.200 ;
        RECT 178.400 137.600 277.600 138.400 ;
        RECT 313.600 137.600 389.600 138.400 ;
        RECT 177.600 136.800 276.000 137.600 ;
        RECT 310.400 136.800 388.800 137.600 ;
        RECT 177.600 136.000 274.400 136.800 ;
        RECT 308.000 136.000 388.800 136.800 ;
        RECT 176.800 135.200 272.800 136.000 ;
        RECT 304.800 135.200 388.000 136.000 ;
        RECT 176.000 134.400 271.200 135.200 ;
        RECT 302.400 134.400 387.200 135.200 ;
        RECT 176.000 133.600 269.600 134.400 ;
        RECT 300.000 133.600 386.400 134.400 ;
        RECT 175.200 132.800 268.000 133.600 ;
        RECT 297.600 132.800 385.600 133.600 ;
        RECT 174.400 132.000 266.400 132.800 ;
        RECT 295.200 132.000 385.600 132.800 ;
        RECT 174.400 131.200 264.800 132.000 ;
        RECT 292.800 131.200 384.800 132.000 ;
        RECT 173.600 130.400 263.200 131.200 ;
        RECT 290.400 130.400 384.000 131.200 ;
        RECT 172.800 129.600 261.600 130.400 ;
        RECT 288.000 129.600 383.200 130.400 ;
        RECT 172.800 128.800 260.000 129.600 ;
        RECT 285.600 128.800 382.400 129.600 ;
        RECT 172.000 128.000 258.400 128.800 ;
        RECT 283.200 128.000 381.600 128.800 ;
        RECT 171.200 127.200 256.800 128.000 ;
        RECT 280.800 127.200 381.600 128.000 ;
        RECT 171.200 126.400 256.000 127.200 ;
        RECT 279.200 126.400 380.800 127.200 ;
        RECT 170.400 125.600 254.400 126.400 ;
        RECT 276.800 125.600 380.000 126.400 ;
        RECT 169.600 124.800 252.800 125.600 ;
        RECT 274.400 124.800 379.200 125.600 ;
        RECT 169.600 124.000 251.200 124.800 ;
        RECT 272.800 124.000 378.400 124.800 ;
        RECT 168.800 123.200 249.600 124.000 ;
        RECT 270.400 123.200 377.600 124.000 ;
        RECT 168.000 122.400 248.000 123.200 ;
        RECT 268.800 122.400 376.800 123.200 ;
        RECT 168.000 121.600 246.400 122.400 ;
        RECT 266.400 121.600 376.000 122.400 ;
        RECT 167.200 120.800 244.800 121.600 ;
        RECT 264.800 120.800 374.400 121.600 ;
        RECT 166.400 120.000 244.000 120.800 ;
        RECT 262.400 120.000 373.600 120.800 ;
        RECT 166.400 119.200 242.400 120.000 ;
        RECT 260.800 119.200 372.800 120.000 ;
        RECT 165.600 118.400 240.800 119.200 ;
        RECT 259.200 118.400 372.000 119.200 ;
        RECT 164.800 117.600 239.200 118.400 ;
        RECT 257.600 117.600 371.200 118.400 ;
        RECT 164.800 116.800 237.600 117.600 ;
        RECT 256.000 116.800 369.600 117.600 ;
        RECT 164.000 116.000 236.000 116.800 ;
        RECT 253.600 116.000 368.800 116.800 ;
        RECT 163.200 115.200 235.200 116.000 ;
        RECT 252.000 115.200 368.000 116.000 ;
        RECT 163.200 114.400 233.600 115.200 ;
        RECT 250.400 114.400 367.200 115.200 ;
        RECT 162.400 113.600 232.000 114.400 ;
        RECT 248.800 113.600 365.600 114.400 ;
        RECT 162.400 112.800 230.400 113.600 ;
        RECT 247.200 112.800 364.800 113.600 ;
        RECT 161.600 112.000 228.800 112.800 ;
        RECT 245.600 112.000 364.000 112.800 ;
        RECT 160.800 111.200 228.000 112.000 ;
        RECT 244.000 111.200 362.400 112.000 ;
        RECT 160.800 110.400 226.400 111.200 ;
        RECT 242.400 110.400 361.600 111.200 ;
        RECT 160.000 109.600 224.800 110.400 ;
        RECT 240.800 109.600 360.000 110.400 ;
        RECT 159.200 108.800 223.200 109.600 ;
        RECT 240.000 108.800 359.200 109.600 ;
        RECT 159.200 108.000 222.400 108.800 ;
        RECT 238.400 108.000 358.400 108.800 ;
        RECT 158.400 107.200 220.800 108.000 ;
        RECT 236.800 107.200 356.800 108.000 ;
        RECT 157.600 106.400 219.200 107.200 ;
        RECT 235.200 106.400 356.000 107.200 ;
        RECT 157.600 105.600 218.400 106.400 ;
        RECT 234.400 105.600 354.400 106.400 ;
        RECT 156.800 104.800 216.800 105.600 ;
        RECT 232.800 104.800 353.600 105.600 ;
        RECT 156.800 104.000 215.200 104.800 ;
        RECT 231.200 104.000 352.000 104.800 ;
        RECT 156.000 103.200 214.400 104.000 ;
        RECT 229.600 103.200 351.200 104.000 ;
        RECT 155.200 102.400 212.800 103.200 ;
        RECT 228.800 102.400 349.600 103.200 ;
        RECT 155.200 101.600 211.200 102.400 ;
        RECT 227.200 101.600 348.000 102.400 ;
        RECT 154.400 100.800 210.400 101.600 ;
        RECT 226.400 100.800 347.200 101.600 ;
        RECT 153.600 100.000 208.800 100.800 ;
        RECT 224.800 100.000 345.600 100.800 ;
        RECT 153.600 99.200 208.000 100.000 ;
        RECT 223.200 99.200 344.800 100.000 ;
        RECT 152.800 98.400 206.400 99.200 ;
        RECT 222.400 98.400 343.200 99.200 ;
        RECT 152.800 97.600 204.800 98.400 ;
        RECT 220.800 97.600 342.400 98.400 ;
        RECT 152.000 96.800 204.000 97.600 ;
        RECT 220.000 96.800 340.800 97.600 ;
        RECT 151.200 96.000 202.400 96.800 ;
        RECT 218.400 96.000 340.000 96.800 ;
        RECT 151.200 95.200 201.600 96.000 ;
        RECT 216.800 95.200 338.400 96.000 ;
        RECT 150.400 94.400 200.000 95.200 ;
        RECT 216.000 94.400 336.800 95.200 ;
        RECT 150.400 93.600 198.400 94.400 ;
        RECT 214.400 93.600 336.000 94.400 ;
        RECT 149.600 92.800 197.600 93.600 ;
        RECT 213.600 92.800 334.400 93.600 ;
        RECT 148.800 92.000 196.000 92.800 ;
        RECT 212.000 92.000 332.800 92.800 ;
        RECT 148.800 91.200 195.200 92.000 ;
        RECT 211.200 91.200 332.000 92.000 ;
        RECT 148.000 90.400 193.600 91.200 ;
        RECT 209.600 90.400 330.400 91.200 ;
        RECT 147.200 89.600 192.800 90.400 ;
        RECT 208.800 89.600 328.800 90.400 ;
        RECT 147.200 88.800 191.200 89.600 ;
        RECT 207.200 88.800 328.000 89.600 ;
        RECT 146.400 88.000 190.400 88.800 ;
        RECT 206.400 88.000 326.400 88.800 ;
        RECT 146.400 87.200 188.800 88.000 ;
        RECT 204.800 87.200 324.800 88.000 ;
        RECT 145.600 86.400 188.000 87.200 ;
        RECT 204.000 86.400 324.000 87.200 ;
        RECT 144.800 85.600 186.400 86.400 ;
        RECT 202.400 85.600 322.400 86.400 ;
        RECT 144.800 84.800 185.600 85.600 ;
        RECT 201.600 84.800 320.800 85.600 ;
        RECT 144.000 84.000 184.000 84.800 ;
        RECT 200.000 84.000 320.000 84.800 ;
        RECT 144.000 83.200 183.200 84.000 ;
        RECT 199.200 83.200 318.400 84.000 ;
        RECT 143.200 82.400 182.400 83.200 ;
        RECT 197.600 82.400 316.800 83.200 ;
        RECT 143.200 81.600 180.800 82.400 ;
        RECT 196.800 81.600 316.000 82.400 ;
        RECT 142.400 80.800 180.000 81.600 ;
        RECT 195.200 80.800 314.400 81.600 ;
        RECT 141.600 80.000 178.400 80.800 ;
        RECT 194.400 80.000 312.800 80.800 ;
        RECT 141.600 79.200 177.600 80.000 ;
        RECT 192.800 79.200 312.000 80.000 ;
        RECT 140.800 78.400 176.000 79.200 ;
        RECT 192.000 78.400 310.400 79.200 ;
        RECT 140.800 77.600 175.200 78.400 ;
        RECT 190.400 77.600 308.800 78.400 ;
        RECT 140.000 76.800 174.400 77.600 ;
        RECT 189.600 76.800 308.000 77.600 ;
        RECT 139.200 76.000 172.800 76.800 ;
        RECT 188.000 76.000 306.400 76.800 ;
        RECT 139.200 75.200 172.000 76.000 ;
        RECT 187.200 75.200 304.800 76.000 ;
        RECT 138.400 74.400 170.400 75.200 ;
        RECT 185.600 74.400 304.000 75.200 ;
        RECT 138.400 73.600 169.600 74.400 ;
        RECT 184.800 73.600 302.400 74.400 ;
        RECT 137.600 72.800 168.800 73.600 ;
        RECT 183.200 72.800 300.800 73.600 ;
        RECT 137.600 72.000 167.200 72.800 ;
        RECT 182.400 72.000 300.000 72.800 ;
        RECT 136.800 71.200 166.400 72.000 ;
        RECT 180.800 71.200 298.400 72.000 ;
        RECT 136.800 70.400 165.600 71.200 ;
        RECT 180.000 70.400 296.800 71.200 ;
        RECT 136.000 69.600 164.000 70.400 ;
        RECT 178.400 69.600 296.000 70.400 ;
        RECT 136.000 68.800 163.200 69.600 ;
        RECT 177.600 68.800 294.400 69.600 ;
        RECT 135.200 68.000 162.400 68.800 ;
        RECT 176.000 68.000 292.800 68.800 ;
        RECT 134.400 67.200 160.800 68.000 ;
        RECT 175.200 67.200 292.000 68.000 ;
        RECT 134.400 66.400 160.000 67.200 ;
        RECT 173.600 66.400 290.400 67.200 ;
        RECT 133.600 65.600 159.200 66.400 ;
        RECT 172.800 65.600 288.800 66.400 ;
        RECT 133.600 64.800 158.400 65.600 ;
        RECT 171.200 64.800 288.000 65.600 ;
        RECT 132.800 64.000 156.800 64.800 ;
        RECT 170.400 64.000 286.400 64.800 ;
        RECT 132.800 63.200 156.000 64.000 ;
        RECT 168.800 63.200 285.600 64.000 ;
        RECT 132.000 62.400 155.200 63.200 ;
        RECT 168.000 62.400 284.000 63.200 ;
        RECT 132.000 61.600 153.600 62.400 ;
        RECT 167.200 61.600 282.400 62.400 ;
        RECT 131.200 60.800 152.800 61.600 ;
        RECT 165.600 60.800 280.800 61.600 ;
        RECT 131.200 60.000 152.000 60.800 ;
        RECT 164.800 60.000 279.200 60.800 ;
        RECT 130.400 59.200 151.200 60.000 ;
        RECT 163.200 59.200 276.800 60.000 ;
        RECT 130.400 58.400 149.600 59.200 ;
        RECT 162.400 58.400 275.200 59.200 ;
        RECT 129.600 57.600 148.800 58.400 ;
        RECT 160.800 57.600 272.800 58.400 ;
        RECT 129.600 56.800 148.000 57.600 ;
        RECT 160.000 56.800 271.200 57.600 ;
        RECT 129.600 56.000 147.200 56.800 ;
        RECT 159.200 56.000 268.800 56.800 ;
        RECT 128.800 55.200 145.600 56.000 ;
        RECT 157.600 55.200 266.400 56.000 ;
        RECT 128.800 54.400 144.800 55.200 ;
        RECT 156.800 54.400 264.800 55.200 ;
        RECT 128.000 53.600 144.000 54.400 ;
        RECT 155.200 53.600 262.400 54.400 ;
        RECT 280.000 53.600 281.600 54.400 ;
        RECT 128.000 52.800 143.200 53.600 ;
        RECT 154.400 52.800 260.800 53.600 ;
        RECT 277.600 52.800 280.800 53.600 ;
        RECT 127.200 52.000 141.600 52.800 ;
        RECT 152.800 52.000 258.400 52.800 ;
        RECT 276.000 52.000 280.000 52.800 ;
        RECT 127.200 51.200 140.800 52.000 ;
        RECT 152.000 51.200 256.800 52.000 ;
        RECT 273.600 51.200 279.200 52.000 ;
        RECT 127.200 50.400 140.000 51.200 ;
        RECT 151.200 50.400 254.400 51.200 ;
        RECT 271.200 50.400 278.400 51.200 ;
        RECT 126.400 49.600 138.400 50.400 ;
        RECT 149.600 49.600 252.800 50.400 ;
        RECT 269.600 49.600 277.600 50.400 ;
        RECT 126.400 48.800 137.600 49.600 ;
        RECT 148.800 48.800 250.400 49.600 ;
        RECT 267.200 48.800 276.800 49.600 ;
        RECT 125.600 48.000 136.800 48.800 ;
        RECT 148.000 48.000 248.800 48.800 ;
        RECT 264.800 48.000 276.000 48.800 ;
        RECT 125.600 47.200 136.000 48.000 ;
        RECT 146.400 47.200 246.400 48.000 ;
        RECT 263.200 47.200 275.200 48.000 ;
        RECT 125.600 46.400 134.400 47.200 ;
        RECT 145.600 46.400 244.800 47.200 ;
        RECT 260.800 46.400 273.600 47.200 ;
        RECT 124.800 45.600 133.600 46.400 ;
        RECT 144.000 45.600 242.400 46.400 ;
        RECT 258.400 45.600 272.800 46.400 ;
        RECT 124.800 44.800 132.800 45.600 ;
        RECT 143.200 44.800 240.000 45.600 ;
        RECT 256.000 44.800 272.000 45.600 ;
        RECT 124.000 44.000 131.200 44.800 ;
        RECT 142.400 44.000 238.400 44.800 ;
        RECT 254.400 44.000 271.200 44.800 ;
        RECT 124.000 43.200 130.400 44.000 ;
        RECT 140.800 43.200 236.000 44.000 ;
        RECT 252.000 43.200 270.400 44.000 ;
        RECT 124.000 42.400 129.600 43.200 ;
        RECT 140.000 42.400 234.400 43.200 ;
        RECT 249.600 42.400 269.600 43.200 ;
        RECT 123.200 41.600 128.000 42.400 ;
        RECT 139.200 41.600 232.000 42.400 ;
        RECT 248.000 41.600 268.800 42.400 ;
        RECT 123.200 40.800 127.200 41.600 ;
        RECT 137.600 40.800 230.400 41.600 ;
        RECT 245.600 40.800 268.000 41.600 ;
        RECT 123.200 40.000 126.400 40.800 ;
        RECT 136.800 40.000 228.000 40.800 ;
        RECT 243.200 40.000 267.200 40.800 ;
        RECT 122.400 39.200 124.800 40.000 ;
        RECT 136.000 39.200 226.400 40.000 ;
        RECT 241.600 39.200 266.400 40.000 ;
        RECT 122.400 38.400 124.000 39.200 ;
        RECT 134.400 38.400 224.000 39.200 ;
        RECT 239.200 38.400 264.800 39.200 ;
        RECT 121.600 37.600 123.200 38.400 ;
        RECT 133.600 37.600 165.600 38.400 ;
        RECT 236.800 37.600 264.000 38.400 ;
        RECT 132.800 36.800 160.000 37.600 ;
        RECT 235.200 36.800 263.200 37.600 ;
        RECT 131.200 36.000 156.800 36.800 ;
        RECT 232.800 36.000 262.400 36.800 ;
        RECT 130.400 35.200 153.600 36.000 ;
        RECT 230.400 35.200 261.600 36.000 ;
        RECT 129.600 34.400 152.000 35.200 ;
        RECT 228.800 34.400 260.800 35.200 ;
        RECT 128.800 33.600 149.600 34.400 ;
        RECT 226.400 33.600 260.000 34.400 ;
        RECT 128.000 32.800 148.000 33.600 ;
        RECT 200.800 32.800 258.400 33.600 ;
        RECT 126.400 32.000 146.400 32.800 ;
        RECT 197.600 32.000 257.600 32.800 ;
        RECT 125.600 31.200 144.000 32.000 ;
        RECT 195.200 31.200 256.800 32.000 ;
        RECT 124.800 30.400 143.200 31.200 ;
        RECT 192.000 30.400 255.200 31.200 ;
        RECT 124.000 29.600 141.600 30.400 ;
        RECT 188.000 29.600 254.400 30.400 ;
        RECT 123.200 28.800 140.000 29.600 ;
        RECT 183.200 28.800 253.600 29.600 ;
        RECT 122.400 28.000 138.400 28.800 ;
        RECT 176.800 28.000 252.800 28.800 ;
        RECT 121.600 27.200 137.600 28.000 ;
        RECT 145.600 27.200 156.000 28.000 ;
        RECT 165.600 27.200 251.200 28.000 ;
        RECT 120.800 26.400 136.000 27.200 ;
        RECT 144.800 26.400 250.400 27.200 ;
        RECT 120.000 25.600 135.200 26.400 ;
        RECT 144.000 25.600 248.800 26.400 ;
        RECT 119.200 24.800 133.600 25.600 ;
        RECT 142.400 24.800 248.000 25.600 ;
        RECT 118.400 24.000 132.800 24.800 ;
        RECT 141.600 24.000 246.400 24.800 ;
        RECT 117.600 23.200 131.200 24.000 ;
        RECT 140.800 23.200 245.600 24.000 ;
        RECT 117.600 22.400 130.400 23.200 ;
        RECT 140.000 22.400 244.000 23.200 ;
        RECT 116.800 21.600 129.600 22.400 ;
        RECT 139.200 21.600 243.200 22.400 ;
        RECT 116.000 20.800 128.000 21.600 ;
        RECT 137.600 20.800 241.600 21.600 ;
        RECT 116.000 20.000 127.200 20.800 ;
        RECT 136.800 20.000 240.000 20.800 ;
        RECT 115.200 19.200 126.400 20.000 ;
        RECT 136.000 19.200 239.200 20.000 ;
        RECT 114.400 18.400 124.800 19.200 ;
        RECT 135.200 18.400 237.600 19.200 ;
        RECT 114.400 17.600 124.000 18.400 ;
        RECT 133.600 17.600 236.000 18.400 ;
        RECT 113.600 16.800 123.200 17.600 ;
        RECT 132.800 16.800 234.400 17.600 ;
        RECT 113.600 16.000 121.600 16.800 ;
        RECT 132.000 16.000 232.800 16.800 ;
        RECT 112.800 15.200 120.800 16.000 ;
        RECT 131.200 15.200 231.200 16.000 ;
        RECT 112.800 14.400 119.200 15.200 ;
        RECT 129.600 14.400 229.600 15.200 ;
        RECT 112.000 13.600 118.400 14.400 ;
        RECT 128.800 13.600 228.000 14.400 ;
        RECT 112.000 12.800 116.800 13.600 ;
        RECT 128.000 12.800 226.400 13.600 ;
        RECT 111.200 12.000 116.000 12.800 ;
        RECT 127.200 12.000 224.000 12.800 ;
        RECT 111.200 11.200 114.400 12.000 ;
        RECT 126.400 11.200 222.400 12.000 ;
        RECT 110.400 10.400 112.800 11.200 ;
        RECT 124.800 10.400 220.000 11.200 ;
        RECT 110.400 9.600 112.000 10.400 ;
        RECT 124.000 9.600 218.400 10.400 ;
        RECT 123.200 8.800 216.000 9.600 ;
        RECT 122.400 8.000 213.600 8.800 ;
        RECT 120.800 7.200 211.200 8.000 ;
        RECT 120.000 6.400 208.800 7.200 ;
        RECT 119.200 5.600 205.600 6.400 ;
        RECT 122.400 4.800 203.200 5.600 ;
        RECT 127.200 4.000 200.000 4.800 ;
        RECT 132.800 3.200 196.000 4.000 ;
        RECT 137.600 2.400 192.800 3.200 ;
        RECT 144.000 1.600 188.000 2.400 ;
        RECT 150.400 0.800 182.400 1.600 ;
        RECT 161.600 0.000 171.200 0.800 ;
  END
END avali_logo
END LIBRARY

