magic
tech gf180mcuD
magscale 1 10
timestamp 1699362100
<< metal1 >>
rect 1344 22762 24640 22796
rect 1344 22710 4126 22762
rect 4178 22710 4230 22762
rect 4282 22710 4334 22762
rect 4386 22710 9950 22762
rect 10002 22710 10054 22762
rect 10106 22710 10158 22762
rect 10210 22710 15774 22762
rect 15826 22710 15878 22762
rect 15930 22710 15982 22762
rect 16034 22710 21598 22762
rect 21650 22710 21702 22762
rect 21754 22710 21806 22762
rect 21858 22710 24640 22762
rect 1344 22676 24640 22710
rect 22430 22594 22482 22606
rect 22430 22530 22482 22542
rect 12686 22482 12738 22494
rect 12686 22418 12738 22430
rect 13134 22370 13186 22382
rect 13134 22306 13186 22318
rect 19630 22370 19682 22382
rect 19954 22318 19966 22370
rect 20018 22318 20030 22370
rect 20850 22318 20862 22370
rect 20914 22318 20926 22370
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 19630 22306 19682 22318
rect 13470 22146 13522 22158
rect 13470 22082 13522 22094
rect 20190 22146 20242 22158
rect 20190 22082 20242 22094
rect 21086 22146 21138 22158
rect 21086 22082 21138 22094
rect 1344 21978 24800 22012
rect 1344 21926 7038 21978
rect 7090 21926 7142 21978
rect 7194 21926 7246 21978
rect 7298 21926 12862 21978
rect 12914 21926 12966 21978
rect 13018 21926 13070 21978
rect 13122 21926 18686 21978
rect 18738 21926 18790 21978
rect 18842 21926 18894 21978
rect 18946 21926 24510 21978
rect 24562 21926 24614 21978
rect 24666 21926 24718 21978
rect 24770 21926 24800 21978
rect 1344 21892 24800 21926
rect 8542 21698 8594 21710
rect 8542 21634 8594 21646
rect 5058 21534 5070 21586
rect 5122 21534 5134 21586
rect 8306 21534 8318 21586
rect 8370 21534 8382 21586
rect 9874 21534 9886 21586
rect 9938 21534 9950 21586
rect 13234 21534 13246 21586
rect 13298 21534 13310 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 21074 21534 21086 21586
rect 21138 21534 21150 21586
rect 5730 21422 5742 21474
rect 5794 21422 5806 21474
rect 7858 21422 7870 21474
rect 7922 21422 7934 21474
rect 10658 21422 10670 21474
rect 10722 21422 10734 21474
rect 12786 21422 12798 21474
rect 12850 21422 12862 21474
rect 13906 21422 13918 21474
rect 13970 21422 13982 21474
rect 16034 21422 16046 21474
rect 16098 21422 16110 21474
rect 18610 21422 18622 21474
rect 18674 21422 18686 21474
rect 20738 21422 20750 21474
rect 20802 21422 20814 21474
rect 21858 21422 21870 21474
rect 21922 21422 21934 21474
rect 23986 21422 23998 21474
rect 24050 21422 24062 21474
rect 1344 21194 24640 21228
rect 1344 21142 4126 21194
rect 4178 21142 4230 21194
rect 4282 21142 4334 21194
rect 4386 21142 9950 21194
rect 10002 21142 10054 21194
rect 10106 21142 10158 21194
rect 10210 21142 15774 21194
rect 15826 21142 15878 21194
rect 15930 21142 15982 21194
rect 16034 21142 21598 21194
rect 21650 21142 21702 21194
rect 21754 21142 21806 21194
rect 21858 21142 24640 21194
rect 1344 21108 24640 21142
rect 10222 21026 10274 21038
rect 9090 20974 9102 21026
rect 9154 20974 9166 21026
rect 21186 20974 21198 21026
rect 21250 21023 21262 21026
rect 21522 21023 21534 21026
rect 21250 20977 21534 21023
rect 21250 20974 21262 20977
rect 21522 20974 21534 20977
rect 21586 20974 21598 21026
rect 10222 20962 10274 20974
rect 21534 20914 21586 20926
rect 18386 20862 18398 20914
rect 18450 20862 18462 20914
rect 23986 20862 23998 20914
rect 24050 20862 24062 20914
rect 21534 20850 21586 20862
rect 7982 20802 8034 20814
rect 10110 20802 10162 20814
rect 8418 20750 8430 20802
rect 8482 20750 8494 20802
rect 8866 20750 8878 20802
rect 8930 20750 8942 20802
rect 9538 20750 9550 20802
rect 9602 20750 9614 20802
rect 7982 20738 8034 20750
rect 10110 20738 10162 20750
rect 10670 20802 10722 20814
rect 19294 20802 19346 20814
rect 15586 20750 15598 20802
rect 15650 20750 15662 20802
rect 19730 20750 19742 20802
rect 19794 20750 19806 20802
rect 22082 20750 22094 20802
rect 22146 20750 22158 20802
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 23650 20750 23662 20802
rect 23714 20750 23726 20802
rect 10670 20738 10722 20750
rect 19294 20738 19346 20750
rect 7870 20690 7922 20702
rect 10222 20690 10274 20702
rect 8530 20638 8542 20690
rect 8594 20638 8606 20690
rect 7870 20626 7922 20638
rect 10222 20626 10274 20638
rect 10782 20690 10834 20702
rect 20190 20690 20242 20702
rect 16258 20638 16270 20690
rect 16322 20638 16334 20690
rect 10782 20626 10834 20638
rect 20190 20626 20242 20638
rect 21870 20690 21922 20702
rect 21870 20626 21922 20638
rect 23214 20690 23266 20702
rect 23214 20626 23266 20638
rect 1344 20410 24800 20444
rect 1344 20358 7038 20410
rect 7090 20358 7142 20410
rect 7194 20358 7246 20410
rect 7298 20358 12862 20410
rect 12914 20358 12966 20410
rect 13018 20358 13070 20410
rect 13122 20358 18686 20410
rect 18738 20358 18790 20410
rect 18842 20358 18894 20410
rect 18946 20358 24510 20410
rect 24562 20358 24614 20410
rect 24666 20358 24718 20410
rect 24770 20358 24800 20410
rect 1344 20324 24800 20358
rect 8766 20242 8818 20254
rect 8766 20178 8818 20190
rect 14030 20242 14082 20254
rect 14030 20178 14082 20190
rect 17502 20242 17554 20254
rect 17502 20178 17554 20190
rect 6974 20130 7026 20142
rect 6974 20066 7026 20078
rect 9550 20130 9602 20142
rect 9550 20066 9602 20078
rect 9998 20130 10050 20142
rect 9998 20066 10050 20078
rect 14254 20130 14306 20142
rect 14254 20066 14306 20078
rect 14926 20130 14978 20142
rect 14926 20066 14978 20078
rect 16494 20130 16546 20142
rect 16494 20066 16546 20078
rect 16606 20130 16658 20142
rect 16606 20066 16658 20078
rect 17726 20130 17778 20142
rect 17726 20066 17778 20078
rect 19630 20130 19682 20142
rect 19630 20066 19682 20078
rect 19854 20130 19906 20142
rect 19854 20066 19906 20078
rect 20302 20130 20354 20142
rect 20302 20066 20354 20078
rect 21198 20130 21250 20142
rect 21198 20066 21250 20078
rect 21310 20130 21362 20142
rect 21310 20066 21362 20078
rect 21422 20130 21474 20142
rect 21422 20066 21474 20078
rect 21982 20130 22034 20142
rect 21982 20066 22034 20078
rect 22206 20130 22258 20142
rect 22206 20066 22258 20078
rect 8654 20018 8706 20030
rect 13918 20018 13970 20030
rect 3490 19966 3502 20018
rect 3554 19966 3566 20018
rect 4162 19966 4174 20018
rect 4226 19966 4238 20018
rect 7970 19966 7982 20018
rect 8034 19966 8046 20018
rect 9762 19966 9774 20018
rect 9826 19966 9838 20018
rect 8654 19954 8706 19966
rect 13918 19954 13970 19966
rect 14366 20018 14418 20030
rect 16830 20018 16882 20030
rect 15138 19966 15150 20018
rect 15202 19966 15214 20018
rect 16034 19966 16046 20018
rect 16098 19966 16110 20018
rect 14366 19954 14418 19966
rect 16830 19954 16882 19966
rect 17390 20018 17442 20030
rect 17390 19954 17442 19966
rect 20078 20018 20130 20030
rect 20078 19954 20130 19966
rect 20414 20018 20466 20030
rect 23214 20018 23266 20030
rect 21746 19966 21758 20018
rect 21810 19966 21822 20018
rect 23538 19966 23550 20018
rect 23602 19966 23614 20018
rect 20414 19954 20466 19966
rect 23214 19954 23266 19966
rect 6862 19906 6914 19918
rect 6290 19854 6302 19906
rect 6354 19854 6366 19906
rect 6862 19842 6914 19854
rect 7310 19906 7362 19918
rect 22878 19906 22930 19918
rect 8194 19854 8206 19906
rect 8258 19854 8270 19906
rect 16482 19854 16494 19906
rect 16546 19854 16558 19906
rect 19506 19854 19518 19906
rect 19570 19854 19582 19906
rect 22082 19854 22094 19906
rect 22146 19854 22158 19906
rect 7310 19842 7362 19854
rect 22878 19842 22930 19854
rect 24110 19906 24162 19918
rect 24110 19842 24162 19854
rect 8766 19794 8818 19806
rect 8766 19730 8818 19742
rect 9886 19794 9938 19806
rect 9886 19730 9938 19742
rect 1344 19626 24640 19660
rect 1344 19574 4126 19626
rect 4178 19574 4230 19626
rect 4282 19574 4334 19626
rect 4386 19574 9950 19626
rect 10002 19574 10054 19626
rect 10106 19574 10158 19626
rect 10210 19574 15774 19626
rect 15826 19574 15878 19626
rect 15930 19574 15982 19626
rect 16034 19574 21598 19626
rect 21650 19574 21702 19626
rect 21754 19574 21806 19626
rect 21858 19574 24640 19626
rect 1344 19540 24640 19574
rect 4958 19458 5010 19470
rect 4958 19394 5010 19406
rect 12014 19458 12066 19470
rect 12014 19394 12066 19406
rect 10334 19346 10386 19358
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 10334 19282 10386 19294
rect 14366 19346 14418 19358
rect 21646 19346 21698 19358
rect 20290 19294 20302 19346
rect 20354 19294 20366 19346
rect 14366 19282 14418 19294
rect 21646 19282 21698 19294
rect 8206 19234 8258 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 7970 19182 7982 19234
rect 8034 19182 8046 19234
rect 8206 19170 8258 19182
rect 8318 19234 8370 19246
rect 8318 19170 8370 19182
rect 10558 19234 10610 19246
rect 10558 19170 10610 19182
rect 11230 19234 11282 19246
rect 11230 19170 11282 19182
rect 12014 19234 12066 19246
rect 12014 19170 12066 19182
rect 12462 19234 12514 19246
rect 12462 19170 12514 19182
rect 12686 19234 12738 19246
rect 12686 19170 12738 19182
rect 14254 19234 14306 19246
rect 14254 19170 14306 19182
rect 14926 19234 14978 19246
rect 14926 19170 14978 19182
rect 15038 19234 15090 19246
rect 15038 19170 15090 19182
rect 15262 19234 15314 19246
rect 15262 19170 15314 19182
rect 15598 19234 15650 19246
rect 15598 19170 15650 19182
rect 16046 19234 16098 19246
rect 16046 19170 16098 19182
rect 17166 19234 17218 19246
rect 22542 19234 22594 19246
rect 17490 19182 17502 19234
rect 17554 19182 17566 19234
rect 21970 19182 21982 19234
rect 22034 19182 22046 19234
rect 17166 19170 17218 19182
rect 22542 19170 22594 19182
rect 22654 19234 22706 19246
rect 22978 19182 22990 19234
rect 23042 19182 23054 19234
rect 22654 19170 22706 19182
rect 5070 19122 5122 19134
rect 2482 19070 2494 19122
rect 2546 19070 2558 19122
rect 5070 19058 5122 19070
rect 9102 19122 9154 19134
rect 9102 19058 9154 19070
rect 9214 19122 9266 19134
rect 9214 19058 9266 19070
rect 11902 19122 11954 19134
rect 11902 19058 11954 19070
rect 13806 19122 13858 19134
rect 13806 19058 13858 19070
rect 14478 19122 14530 19134
rect 14478 19058 14530 19070
rect 15486 19122 15538 19134
rect 24222 19122 24274 19134
rect 18162 19070 18174 19122
rect 18226 19070 18238 19122
rect 15486 19058 15538 19070
rect 24222 19058 24274 19070
rect 7758 19010 7810 19022
rect 9438 19010 9490 19022
rect 8754 18958 8766 19010
rect 8818 18958 8830 19010
rect 7758 18946 7810 18958
rect 9438 18946 9490 18958
rect 10110 19010 10162 19022
rect 11342 19010 11394 19022
rect 10882 18958 10894 19010
rect 10946 18958 10958 19010
rect 10110 18946 10162 18958
rect 11342 18946 11394 18958
rect 11566 19010 11618 19022
rect 11566 18946 11618 18958
rect 13918 19010 13970 19022
rect 13918 18946 13970 18958
rect 16158 19010 16210 19022
rect 16158 18946 16210 18958
rect 16494 19010 16546 19022
rect 16494 18946 16546 18958
rect 16606 19010 16658 19022
rect 16606 18946 16658 18958
rect 16830 19010 16882 19022
rect 16830 18946 16882 18958
rect 22206 19010 22258 19022
rect 22206 18946 22258 18958
rect 23886 19010 23938 19022
rect 23886 18946 23938 18958
rect 1344 18842 24800 18876
rect 1344 18790 7038 18842
rect 7090 18790 7142 18842
rect 7194 18790 7246 18842
rect 7298 18790 12862 18842
rect 12914 18790 12966 18842
rect 13018 18790 13070 18842
rect 13122 18790 18686 18842
rect 18738 18790 18790 18842
rect 18842 18790 18894 18842
rect 18946 18790 24510 18842
rect 24562 18790 24614 18842
rect 24666 18790 24718 18842
rect 24770 18790 24800 18842
rect 1344 18756 24800 18790
rect 8206 18674 8258 18686
rect 8206 18610 8258 18622
rect 8430 18674 8482 18686
rect 8430 18610 8482 18622
rect 8990 18674 9042 18686
rect 8990 18610 9042 18622
rect 11566 18674 11618 18686
rect 11566 18610 11618 18622
rect 13358 18674 13410 18686
rect 13358 18610 13410 18622
rect 14814 18674 14866 18686
rect 14814 18610 14866 18622
rect 15486 18674 15538 18686
rect 15486 18610 15538 18622
rect 18174 18674 18226 18686
rect 18174 18610 18226 18622
rect 20190 18674 20242 18686
rect 20190 18610 20242 18622
rect 3390 18562 3442 18574
rect 6190 18562 6242 18574
rect 8094 18562 8146 18574
rect 10446 18562 10498 18574
rect 5618 18510 5630 18562
rect 5682 18510 5694 18562
rect 7074 18510 7086 18562
rect 7138 18510 7150 18562
rect 8642 18510 8654 18562
rect 8706 18510 8718 18562
rect 3390 18498 3442 18510
rect 6190 18498 6242 18510
rect 8094 18498 8146 18510
rect 10446 18498 10498 18510
rect 11342 18562 11394 18574
rect 11342 18498 11394 18510
rect 11790 18562 11842 18574
rect 12674 18510 12686 18562
rect 12738 18510 12750 18562
rect 13682 18510 13694 18562
rect 13746 18510 13758 18562
rect 17378 18510 17390 18562
rect 17442 18510 17454 18562
rect 19730 18510 19742 18562
rect 19794 18510 19806 18562
rect 11790 18498 11842 18510
rect 3950 18450 4002 18462
rect 9774 18450 9826 18462
rect 3602 18398 3614 18450
rect 3666 18398 3678 18450
rect 4386 18398 4398 18450
rect 4450 18398 4462 18450
rect 4834 18398 4846 18450
rect 4898 18398 4910 18450
rect 5506 18398 5518 18450
rect 5570 18398 5582 18450
rect 7298 18398 7310 18450
rect 7362 18398 7374 18450
rect 3950 18386 4002 18398
rect 9774 18386 9826 18398
rect 10782 18450 10834 18462
rect 10782 18386 10834 18398
rect 11006 18450 11058 18462
rect 11006 18386 11058 18398
rect 12238 18450 12290 18462
rect 14702 18450 14754 18462
rect 18062 18450 18114 18462
rect 12898 18398 12910 18450
rect 12962 18398 12974 18450
rect 15698 18398 15710 18450
rect 15762 18398 15774 18450
rect 17602 18398 17614 18450
rect 17666 18398 17678 18450
rect 18386 18398 18398 18450
rect 18450 18398 18462 18450
rect 19506 18398 19518 18450
rect 19570 18398 19582 18450
rect 20962 18398 20974 18450
rect 21026 18398 21038 18450
rect 12238 18386 12290 18398
rect 14702 18386 14754 18398
rect 18062 18386 18114 18398
rect 9550 18338 9602 18350
rect 9550 18274 9602 18286
rect 10558 18338 10610 18350
rect 10558 18274 10610 18286
rect 14926 18338 14978 18350
rect 20066 18286 20078 18338
rect 20130 18286 20142 18338
rect 21746 18286 21758 18338
rect 21810 18286 21822 18338
rect 23874 18286 23886 18338
rect 23938 18286 23950 18338
rect 14926 18274 14978 18286
rect 3278 18226 3330 18238
rect 3278 18162 3330 18174
rect 4062 18226 4114 18238
rect 4062 18162 4114 18174
rect 6526 18226 6578 18238
rect 11454 18226 11506 18238
rect 10098 18174 10110 18226
rect 10162 18174 10174 18226
rect 6526 18162 6578 18174
rect 11454 18162 11506 18174
rect 12126 18226 12178 18238
rect 12126 18162 12178 18174
rect 14366 18226 14418 18238
rect 14366 18162 14418 18174
rect 14478 18226 14530 18238
rect 14478 18162 14530 18174
rect 15374 18226 15426 18238
rect 15374 18162 15426 18174
rect 20414 18226 20466 18238
rect 20414 18162 20466 18174
rect 1344 18058 24640 18092
rect 1344 18006 4126 18058
rect 4178 18006 4230 18058
rect 4282 18006 4334 18058
rect 4386 18006 9950 18058
rect 10002 18006 10054 18058
rect 10106 18006 10158 18058
rect 10210 18006 15774 18058
rect 15826 18006 15878 18058
rect 15930 18006 15982 18058
rect 16034 18006 21598 18058
rect 21650 18006 21702 18058
rect 21754 18006 21806 18058
rect 21858 18006 24640 18058
rect 1344 17972 24640 18006
rect 2942 17890 2994 17902
rect 2942 17826 2994 17838
rect 3614 17890 3666 17902
rect 3614 17826 3666 17838
rect 4622 17890 4674 17902
rect 4622 17826 4674 17838
rect 14254 17890 14306 17902
rect 14254 17826 14306 17838
rect 16494 17890 16546 17902
rect 22206 17890 22258 17902
rect 21298 17838 21310 17890
rect 21362 17838 21374 17890
rect 16494 17826 16546 17838
rect 22206 17826 22258 17838
rect 22318 17890 22370 17902
rect 22318 17826 22370 17838
rect 22654 17890 22706 17902
rect 22654 17826 22706 17838
rect 3838 17778 3890 17790
rect 3838 17714 3890 17726
rect 6302 17778 6354 17790
rect 7186 17726 7198 17778
rect 7250 17726 7262 17778
rect 8866 17726 8878 17778
rect 8930 17726 8942 17778
rect 20290 17726 20302 17778
rect 20354 17726 20366 17778
rect 6302 17714 6354 17726
rect 2830 17666 2882 17678
rect 2370 17614 2382 17666
rect 2434 17614 2446 17666
rect 2830 17602 2882 17614
rect 4734 17666 4786 17678
rect 14142 17666 14194 17678
rect 5730 17614 5742 17666
rect 5794 17614 5806 17666
rect 6738 17614 6750 17666
rect 6802 17614 6814 17666
rect 12674 17614 12686 17666
rect 12738 17614 12750 17666
rect 4734 17602 4786 17614
rect 14142 17602 14194 17614
rect 16158 17666 16210 17678
rect 21646 17666 21698 17678
rect 17490 17614 17502 17666
rect 17554 17614 17566 17666
rect 16158 17602 16210 17614
rect 21646 17602 21698 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 22542 17666 22594 17678
rect 22542 17602 22594 17614
rect 23214 17666 23266 17678
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 23214 17602 23266 17614
rect 4622 17554 4674 17566
rect 4622 17490 4674 17502
rect 15934 17554 15986 17566
rect 15934 17490 15986 17502
rect 16830 17554 16882 17566
rect 23102 17554 23154 17566
rect 18162 17502 18174 17554
rect 18226 17502 18238 17554
rect 16830 17490 16882 17502
rect 23102 17490 23154 17502
rect 14254 17442 14306 17454
rect 2146 17390 2158 17442
rect 2210 17390 2222 17442
rect 3266 17390 3278 17442
rect 3330 17390 3342 17442
rect 5954 17390 5966 17442
rect 6018 17390 6030 17442
rect 14254 17378 14306 17390
rect 16942 17442 16994 17454
rect 16942 17378 16994 17390
rect 17166 17442 17218 17454
rect 17166 17378 17218 17390
rect 1344 17274 24800 17308
rect 1344 17222 7038 17274
rect 7090 17222 7142 17274
rect 7194 17222 7246 17274
rect 7298 17222 12862 17274
rect 12914 17222 12966 17274
rect 13018 17222 13070 17274
rect 13122 17222 18686 17274
rect 18738 17222 18790 17274
rect 18842 17222 18894 17274
rect 18946 17222 24510 17274
rect 24562 17222 24614 17274
rect 24666 17222 24718 17274
rect 24770 17222 24800 17274
rect 1344 17188 24800 17222
rect 5966 17106 6018 17118
rect 5966 17042 6018 17054
rect 6302 17106 6354 17118
rect 6302 17042 6354 17054
rect 5182 16994 5234 17006
rect 8542 16994 8594 17006
rect 5618 16942 5630 16994
rect 5682 16942 5694 16994
rect 7298 16942 7310 16994
rect 7362 16942 7374 16994
rect 5182 16930 5234 16942
rect 8542 16930 8594 16942
rect 14142 16994 14194 17006
rect 14142 16930 14194 16942
rect 16270 16994 16322 17006
rect 20962 16942 20974 16994
rect 21026 16942 21038 16994
rect 16270 16930 16322 16942
rect 6638 16882 6690 16894
rect 6638 16818 6690 16830
rect 7646 16882 7698 16894
rect 7646 16818 7698 16830
rect 8094 16882 8146 16894
rect 8094 16818 8146 16830
rect 9438 16882 9490 16894
rect 9438 16818 9490 16830
rect 10110 16882 10162 16894
rect 10110 16818 10162 16830
rect 10334 16882 10386 16894
rect 16606 16882 16658 16894
rect 22878 16882 22930 16894
rect 10882 16830 10894 16882
rect 10946 16830 10958 16882
rect 17378 16830 17390 16882
rect 17442 16830 17454 16882
rect 10334 16818 10386 16830
rect 16606 16818 16658 16830
rect 22878 16818 22930 16830
rect 23102 16882 23154 16894
rect 23102 16818 23154 16830
rect 23438 16882 23490 16894
rect 23438 16818 23490 16830
rect 23550 16882 23602 16894
rect 23550 16818 23602 16830
rect 9886 16770 9938 16782
rect 11666 16718 11678 16770
rect 11730 16718 11742 16770
rect 13794 16718 13806 16770
rect 13858 16718 13870 16770
rect 9886 16706 9938 16718
rect 5294 16658 5346 16670
rect 5294 16594 5346 16606
rect 7982 16658 8034 16670
rect 7982 16594 8034 16606
rect 14254 16658 14306 16670
rect 23986 16606 23998 16658
rect 24050 16606 24062 16658
rect 14254 16594 14306 16606
rect 1344 16490 24640 16524
rect 1344 16438 4126 16490
rect 4178 16438 4230 16490
rect 4282 16438 4334 16490
rect 4386 16438 9950 16490
rect 10002 16438 10054 16490
rect 10106 16438 10158 16490
rect 10210 16438 15774 16490
rect 15826 16438 15878 16490
rect 15930 16438 15982 16490
rect 16034 16438 21598 16490
rect 21650 16438 21702 16490
rect 21754 16438 21806 16490
rect 21858 16438 24640 16490
rect 1344 16404 24640 16438
rect 2830 16322 2882 16334
rect 21298 16270 21310 16322
rect 21362 16270 21374 16322
rect 2830 16258 2882 16270
rect 12686 16210 12738 16222
rect 10210 16158 10222 16210
rect 10274 16158 10286 16210
rect 23426 16158 23438 16210
rect 23490 16158 23502 16210
rect 12686 16146 12738 16158
rect 11566 16098 11618 16110
rect 4834 16046 4846 16098
rect 4898 16046 4910 16098
rect 5842 16046 5854 16098
rect 5906 16046 5918 16098
rect 6066 16046 6078 16098
rect 6130 16046 6142 16098
rect 7410 16046 7422 16098
rect 7474 16046 7486 16098
rect 11566 16034 11618 16046
rect 11902 16098 11954 16110
rect 16718 16098 16770 16110
rect 14578 16046 14590 16098
rect 14642 16046 14654 16098
rect 11902 16034 11954 16046
rect 16718 16034 16770 16046
rect 19070 16098 19122 16110
rect 19070 16034 19122 16046
rect 21646 16098 21698 16110
rect 21646 16034 21698 16046
rect 21870 16098 21922 16110
rect 23202 16046 23214 16098
rect 23266 16046 23278 16098
rect 24210 16046 24222 16098
rect 24274 16046 24286 16098
rect 21870 16034 21922 16046
rect 4062 15986 4114 15998
rect 3154 15934 3166 15986
rect 3218 15934 3230 15986
rect 3602 15934 3614 15986
rect 3666 15934 3678 15986
rect 4062 15922 4114 15934
rect 4286 15986 4338 15998
rect 4286 15922 4338 15934
rect 4398 15986 4450 15998
rect 11230 15986 11282 15998
rect 8082 15934 8094 15986
rect 8146 15934 8158 15986
rect 4398 15922 4450 15934
rect 11230 15922 11282 15934
rect 12126 15986 12178 15998
rect 12126 15922 12178 15934
rect 12238 15986 12290 15998
rect 17726 15986 17778 15998
rect 14690 15934 14702 15986
rect 14754 15934 14766 15986
rect 22530 15934 22542 15986
rect 22594 15934 22606 15986
rect 24098 15934 24110 15986
rect 24162 15934 24174 15986
rect 12238 15922 12290 15934
rect 17726 15922 17778 15934
rect 2494 15874 2546 15886
rect 2494 15810 2546 15822
rect 4174 15874 4226 15886
rect 4174 15810 4226 15822
rect 6302 15874 6354 15886
rect 6302 15810 6354 15822
rect 6414 15874 6466 15886
rect 18274 15822 18286 15874
rect 18338 15822 18350 15874
rect 18722 15822 18734 15874
rect 18786 15822 18798 15874
rect 6414 15810 6466 15822
rect 1344 15706 24800 15740
rect 1344 15654 7038 15706
rect 7090 15654 7142 15706
rect 7194 15654 7246 15706
rect 7298 15654 12862 15706
rect 12914 15654 12966 15706
rect 13018 15654 13070 15706
rect 13122 15654 18686 15706
rect 18738 15654 18790 15706
rect 18842 15654 18894 15706
rect 18946 15654 24510 15706
rect 24562 15654 24614 15706
rect 24666 15654 24718 15706
rect 24770 15654 24800 15706
rect 1344 15620 24800 15654
rect 8542 15538 8594 15550
rect 2930 15486 2942 15538
rect 2994 15486 3006 15538
rect 5954 15486 5966 15538
rect 6018 15486 6030 15538
rect 8082 15486 8094 15538
rect 8146 15486 8158 15538
rect 8542 15474 8594 15486
rect 13022 15538 13074 15550
rect 13022 15474 13074 15486
rect 16494 15538 16546 15550
rect 16494 15474 16546 15486
rect 18510 15538 18562 15550
rect 21410 15486 21422 15538
rect 21474 15486 21486 15538
rect 18510 15474 18562 15486
rect 2046 15426 2098 15438
rect 2046 15362 2098 15374
rect 2270 15426 2322 15438
rect 8654 15426 8706 15438
rect 2818 15374 2830 15426
rect 2882 15374 2894 15426
rect 3826 15374 3838 15426
rect 3890 15374 3902 15426
rect 5282 15374 5294 15426
rect 5346 15374 5358 15426
rect 5842 15374 5854 15426
rect 5906 15374 5918 15426
rect 7410 15374 7422 15426
rect 7474 15374 7486 15426
rect 2270 15362 2322 15374
rect 8654 15362 8706 15374
rect 13806 15426 13858 15438
rect 13806 15362 13858 15374
rect 14142 15426 14194 15438
rect 17614 15426 17666 15438
rect 16146 15374 16158 15426
rect 16210 15374 16222 15426
rect 14142 15362 14194 15374
rect 17614 15362 17666 15374
rect 18846 15426 18898 15438
rect 18846 15362 18898 15374
rect 19518 15426 19570 15438
rect 19518 15362 19570 15374
rect 21534 15426 21586 15438
rect 21534 15362 21586 15374
rect 22990 15426 23042 15438
rect 22990 15362 23042 15374
rect 2606 15314 2658 15326
rect 13358 15314 13410 15326
rect 3378 15262 3390 15314
rect 3442 15262 3454 15314
rect 4386 15262 4398 15314
rect 4450 15262 4462 15314
rect 4722 15262 4734 15314
rect 4786 15262 4798 15314
rect 6402 15262 6414 15314
rect 6466 15262 6478 15314
rect 6738 15262 6750 15314
rect 6802 15262 6814 15314
rect 7858 15262 7870 15314
rect 7922 15262 7934 15314
rect 13122 15262 13134 15314
rect 13186 15262 13198 15314
rect 2606 15250 2658 15262
rect 13358 15250 13410 15262
rect 13470 15314 13522 15326
rect 13470 15250 13522 15262
rect 14254 15314 14306 15326
rect 15598 15314 15650 15326
rect 17726 15314 17778 15326
rect 14578 15262 14590 15314
rect 14642 15262 14654 15314
rect 15810 15262 15822 15314
rect 15874 15262 15886 15314
rect 17378 15262 17390 15314
rect 17442 15262 17454 15314
rect 14254 15250 14306 15262
rect 15598 15250 15650 15262
rect 17726 15250 17778 15262
rect 19630 15314 19682 15326
rect 19630 15250 19682 15262
rect 19854 15314 19906 15326
rect 24110 15314 24162 15326
rect 20402 15262 20414 15314
rect 20466 15262 20478 15314
rect 19854 15250 19906 15262
rect 24110 15250 24162 15262
rect 2158 15202 2210 15214
rect 15486 15202 15538 15214
rect 4834 15150 4846 15202
rect 4898 15150 4910 15202
rect 2158 15138 2210 15150
rect 15486 15138 15538 15150
rect 3054 15090 3106 15102
rect 3054 15026 3106 15038
rect 8542 15090 8594 15102
rect 19966 15090 20018 15102
rect 18162 15038 18174 15090
rect 18226 15038 18238 15090
rect 8542 15026 8594 15038
rect 19966 15026 20018 15038
rect 1344 14922 24640 14956
rect 1344 14870 4126 14922
rect 4178 14870 4230 14922
rect 4282 14870 4334 14922
rect 4386 14870 9950 14922
rect 10002 14870 10054 14922
rect 10106 14870 10158 14922
rect 10210 14870 15774 14922
rect 15826 14870 15878 14922
rect 15930 14870 15982 14922
rect 16034 14870 21598 14922
rect 21650 14870 21702 14922
rect 21754 14870 21806 14922
rect 21858 14870 24640 14922
rect 1344 14836 24640 14870
rect 2270 14754 2322 14766
rect 2270 14690 2322 14702
rect 12910 14754 12962 14766
rect 12910 14690 12962 14702
rect 20078 14754 20130 14766
rect 20078 14690 20130 14702
rect 20414 14754 20466 14766
rect 20414 14690 20466 14702
rect 20750 14754 20802 14766
rect 20750 14690 20802 14702
rect 22094 14754 22146 14766
rect 22094 14690 22146 14702
rect 2830 14642 2882 14654
rect 7870 14642 7922 14654
rect 12798 14642 12850 14654
rect 19966 14642 20018 14654
rect 23550 14642 23602 14654
rect 6290 14590 6302 14642
rect 6354 14590 6366 14642
rect 12002 14590 12014 14642
rect 12066 14590 12078 14642
rect 17154 14590 17166 14642
rect 17218 14590 17230 14642
rect 22642 14590 22654 14642
rect 22706 14590 22718 14642
rect 2830 14578 2882 14590
rect 7870 14578 7922 14590
rect 12798 14578 12850 14590
rect 19966 14578 20018 14590
rect 23550 14578 23602 14590
rect 3278 14530 3330 14542
rect 2594 14478 2606 14530
rect 2658 14478 2670 14530
rect 3278 14466 3330 14478
rect 3614 14530 3666 14542
rect 3614 14466 3666 14478
rect 4174 14530 4226 14542
rect 4174 14466 4226 14478
rect 4622 14530 4674 14542
rect 4622 14466 4674 14478
rect 4846 14530 4898 14542
rect 8094 14530 8146 14542
rect 12574 14530 12626 14542
rect 22318 14530 22370 14542
rect 6514 14478 6526 14530
rect 6578 14478 6590 14530
rect 9202 14478 9214 14530
rect 9266 14478 9278 14530
rect 13458 14478 13470 14530
rect 13522 14478 13534 14530
rect 19282 14478 19294 14530
rect 19346 14478 19358 14530
rect 23090 14478 23102 14530
rect 23154 14478 23166 14530
rect 4846 14466 4898 14478
rect 8094 14466 8146 14478
rect 12574 14466 12626 14478
rect 22318 14466 22370 14478
rect 2718 14418 2770 14430
rect 2718 14354 2770 14366
rect 3502 14418 3554 14430
rect 3502 14354 3554 14366
rect 7198 14418 7250 14430
rect 19854 14418 19906 14430
rect 9874 14366 9886 14418
rect 9938 14366 9950 14418
rect 7198 14354 7250 14366
rect 19854 14354 19906 14366
rect 20638 14418 20690 14430
rect 20638 14354 20690 14366
rect 21758 14418 21810 14430
rect 21758 14354 21810 14366
rect 23886 14418 23938 14430
rect 23886 14354 23938 14366
rect 24222 14418 24274 14430
rect 24222 14354 24274 14366
rect 2942 14306 2994 14318
rect 2942 14242 2994 14254
rect 4398 14306 4450 14318
rect 19070 14306 19122 14318
rect 8418 14254 8430 14306
rect 8482 14254 8494 14306
rect 4398 14242 4450 14254
rect 19070 14242 19122 14254
rect 21534 14306 21586 14318
rect 21534 14242 21586 14254
rect 21982 14306 22034 14318
rect 21982 14242 22034 14254
rect 1344 14138 24800 14172
rect 1344 14086 7038 14138
rect 7090 14086 7142 14138
rect 7194 14086 7246 14138
rect 7298 14086 12862 14138
rect 12914 14086 12966 14138
rect 13018 14086 13070 14138
rect 13122 14086 18686 14138
rect 18738 14086 18790 14138
rect 18842 14086 18894 14138
rect 18946 14086 24510 14138
rect 24562 14086 24614 14138
rect 24666 14086 24718 14138
rect 24770 14086 24800 14138
rect 1344 14052 24800 14086
rect 5966 13970 6018 13982
rect 5966 13906 6018 13918
rect 9886 13970 9938 13982
rect 9886 13906 9938 13918
rect 14702 13970 14754 13982
rect 14702 13906 14754 13918
rect 16494 13970 16546 13982
rect 16494 13906 16546 13918
rect 4958 13858 5010 13870
rect 15374 13858 15426 13870
rect 23886 13858 23938 13870
rect 2482 13806 2494 13858
rect 2546 13806 2558 13858
rect 12114 13806 12126 13858
rect 12178 13806 12190 13858
rect 18162 13806 18174 13858
rect 18226 13806 18238 13858
rect 4958 13794 5010 13806
rect 15374 13794 15426 13806
rect 23886 13794 23938 13806
rect 24222 13858 24274 13870
rect 24222 13794 24274 13806
rect 5182 13746 5234 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 5182 13682 5234 13694
rect 6078 13746 6130 13758
rect 6078 13682 6130 13694
rect 6302 13746 6354 13758
rect 6302 13682 6354 13694
rect 9550 13746 9602 13758
rect 15598 13746 15650 13758
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 14914 13694 14926 13746
rect 14978 13694 14990 13746
rect 17490 13694 17502 13746
rect 17554 13694 17566 13746
rect 20626 13694 20638 13746
rect 20690 13694 20702 13746
rect 9550 13682 9602 13694
rect 15598 13682 15650 13694
rect 16382 13634 16434 13646
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 14242 13582 14254 13634
rect 14306 13582 14318 13634
rect 20290 13582 20302 13634
rect 20354 13582 20366 13634
rect 21410 13582 21422 13634
rect 21474 13582 21486 13634
rect 23538 13582 23550 13634
rect 23602 13582 23614 13634
rect 16382 13570 16434 13582
rect 5518 13522 5570 13534
rect 5518 13458 5570 13470
rect 5966 13522 6018 13534
rect 5966 13458 6018 13470
rect 14590 13522 14642 13534
rect 14590 13458 14642 13470
rect 15934 13522 15986 13534
rect 15934 13458 15986 13470
rect 1344 13354 24640 13388
rect 1344 13302 4126 13354
rect 4178 13302 4230 13354
rect 4282 13302 4334 13354
rect 4386 13302 9950 13354
rect 10002 13302 10054 13354
rect 10106 13302 10158 13354
rect 10210 13302 15774 13354
rect 15826 13302 15878 13354
rect 15930 13302 15982 13354
rect 16034 13302 21598 13354
rect 21650 13302 21702 13354
rect 21754 13302 21806 13354
rect 21858 13302 24640 13354
rect 1344 13268 24640 13302
rect 3054 13186 3106 13198
rect 3054 13122 3106 13134
rect 20862 13186 20914 13198
rect 20862 13122 20914 13134
rect 14030 13074 14082 13086
rect 19406 13074 19458 13086
rect 8642 13022 8654 13074
rect 8706 13022 8718 13074
rect 10770 13022 10782 13074
rect 10834 13022 10846 13074
rect 14354 13022 14366 13074
rect 14418 13022 14430 13074
rect 14030 13010 14082 13022
rect 19406 13010 19458 13022
rect 22430 13074 22482 13086
rect 23314 13022 23326 13074
rect 23378 13022 23390 13074
rect 22430 13010 22482 13022
rect 6190 12962 6242 12974
rect 19854 12962 19906 12974
rect 3378 12910 3390 12962
rect 3442 12910 3454 12962
rect 4946 12910 4958 12962
rect 5010 12910 5022 12962
rect 7858 12910 7870 12962
rect 7922 12910 7934 12962
rect 13570 12910 13582 12962
rect 13634 12910 13646 12962
rect 17266 12910 17278 12962
rect 17330 12910 17342 12962
rect 19170 12910 19182 12962
rect 19234 12910 19246 12962
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 23090 12910 23102 12962
rect 23154 12910 23166 12962
rect 6190 12898 6242 12910
rect 19854 12898 19906 12910
rect 12574 12850 12626 12862
rect 18958 12850 19010 12862
rect 16482 12798 16494 12850
rect 16546 12798 16558 12850
rect 12574 12786 12626 12798
rect 18958 12786 19010 12798
rect 19518 12850 19570 12862
rect 21870 12850 21922 12862
rect 19954 12798 19966 12850
rect 20018 12798 20030 12850
rect 20290 12798 20302 12850
rect 20354 12798 20366 12850
rect 19518 12786 19570 12798
rect 21870 12786 21922 12798
rect 24222 12850 24274 12862
rect 24222 12786 24274 12798
rect 3166 12738 3218 12750
rect 3166 12674 3218 12686
rect 4734 12738 4786 12750
rect 4734 12674 4786 12686
rect 6526 12738 6578 12750
rect 6526 12674 6578 12686
rect 12238 12738 12290 12750
rect 12238 12674 12290 12686
rect 21310 12738 21362 12750
rect 21310 12674 21362 12686
rect 21422 12738 21474 12750
rect 21422 12674 21474 12686
rect 21646 12738 21698 12750
rect 21646 12674 21698 12686
rect 23886 12738 23938 12750
rect 23886 12674 23938 12686
rect 1344 12570 24800 12604
rect 1344 12518 7038 12570
rect 7090 12518 7142 12570
rect 7194 12518 7246 12570
rect 7298 12518 12862 12570
rect 12914 12518 12966 12570
rect 13018 12518 13070 12570
rect 13122 12518 18686 12570
rect 18738 12518 18790 12570
rect 18842 12518 18894 12570
rect 18946 12518 24510 12570
rect 24562 12518 24614 12570
rect 24666 12518 24718 12570
rect 24770 12518 24800 12570
rect 1344 12484 24800 12518
rect 15598 12402 15650 12414
rect 15598 12338 15650 12350
rect 16158 12402 16210 12414
rect 17390 12402 17442 12414
rect 16482 12350 16494 12402
rect 16546 12350 16558 12402
rect 16158 12338 16210 12350
rect 17390 12338 17442 12350
rect 21982 12402 22034 12414
rect 21982 12338 22034 12350
rect 18398 12290 18450 12302
rect 21646 12290 21698 12302
rect 2706 12238 2718 12290
rect 2770 12238 2782 12290
rect 6626 12238 6638 12290
rect 6690 12238 6702 12290
rect 9762 12238 9774 12290
rect 9826 12238 9838 12290
rect 12002 12238 12014 12290
rect 12066 12238 12078 12290
rect 19730 12238 19742 12290
rect 19794 12238 19806 12290
rect 18398 12226 18450 12238
rect 21646 12226 21698 12238
rect 23662 12290 23714 12302
rect 23662 12226 23714 12238
rect 15374 12178 15426 12190
rect 1922 12126 1934 12178
rect 1986 12126 1998 12178
rect 5842 12126 5854 12178
rect 5906 12126 5918 12178
rect 9986 12126 9998 12178
rect 10050 12126 10062 12178
rect 11218 12126 11230 12178
rect 11282 12126 11294 12178
rect 15138 12126 15150 12178
rect 15202 12126 15214 12178
rect 15374 12114 15426 12126
rect 15710 12178 15762 12190
rect 20078 12178 20130 12190
rect 18946 12126 18958 12178
rect 19010 12126 19022 12178
rect 22194 12126 22206 12178
rect 22258 12126 22270 12178
rect 22642 12126 22654 12178
rect 22706 12126 22718 12178
rect 15710 12114 15762 12126
rect 20078 12114 20130 12126
rect 10446 12066 10498 12078
rect 15486 12066 15538 12078
rect 4834 12014 4846 12066
rect 4898 12014 4910 12066
rect 8754 12014 8766 12066
rect 8818 12014 8830 12066
rect 14130 12014 14142 12066
rect 14194 12014 14206 12066
rect 10446 12002 10498 12014
rect 15486 12002 15538 12014
rect 17502 12066 17554 12078
rect 19282 12014 19294 12066
rect 19346 12014 19358 12066
rect 17502 12002 17554 12014
rect 10782 11954 10834 11966
rect 10782 11890 10834 11902
rect 1344 11786 24640 11820
rect 1344 11734 4126 11786
rect 4178 11734 4230 11786
rect 4282 11734 4334 11786
rect 4386 11734 9950 11786
rect 10002 11734 10054 11786
rect 10106 11734 10158 11786
rect 10210 11734 15774 11786
rect 15826 11734 15878 11786
rect 15930 11734 15982 11786
rect 16034 11734 21598 11786
rect 21650 11734 21702 11786
rect 21754 11734 21806 11786
rect 21858 11734 24640 11786
rect 1344 11700 24640 11734
rect 13582 11618 13634 11630
rect 13582 11554 13634 11566
rect 13918 11618 13970 11630
rect 13918 11554 13970 11566
rect 21310 11506 21362 11518
rect 6738 11454 6750 11506
rect 6802 11454 6814 11506
rect 21310 11442 21362 11454
rect 23662 11506 23714 11518
rect 23662 11442 23714 11454
rect 24334 11506 24386 11518
rect 24334 11442 24386 11454
rect 21422 11394 21474 11406
rect 22766 11394 22818 11406
rect 11554 11342 11566 11394
rect 11618 11342 11630 11394
rect 14690 11342 14702 11394
rect 14754 11342 14766 11394
rect 16930 11342 16942 11394
rect 16994 11342 17006 11394
rect 21970 11342 21982 11394
rect 22034 11342 22046 11394
rect 23090 11342 23102 11394
rect 23154 11342 23166 11394
rect 21422 11330 21474 11342
rect 22766 11330 22818 11342
rect 14466 11230 14478 11282
rect 14530 11230 14542 11282
rect 17490 11230 17502 11282
rect 17554 11230 17566 11282
rect 1344 11002 24800 11036
rect 1344 10950 7038 11002
rect 7090 10950 7142 11002
rect 7194 10950 7246 11002
rect 7298 10950 12862 11002
rect 12914 10950 12966 11002
rect 13018 10950 13070 11002
rect 13122 10950 18686 11002
rect 18738 10950 18790 11002
rect 18842 10950 18894 11002
rect 18946 10950 24510 11002
rect 24562 10950 24614 11002
rect 24666 10950 24718 11002
rect 24770 10950 24800 11002
rect 1344 10916 24800 10950
rect 3166 10834 3218 10846
rect 3166 10770 3218 10782
rect 11902 10834 11954 10846
rect 11902 10770 11954 10782
rect 16046 10834 16098 10846
rect 16046 10770 16098 10782
rect 16494 10834 16546 10846
rect 16494 10770 16546 10782
rect 16606 10834 16658 10846
rect 22306 10782 22318 10834
rect 22370 10782 22382 10834
rect 16606 10770 16658 10782
rect 2494 10722 2546 10734
rect 20862 10722 20914 10734
rect 4274 10670 4286 10722
rect 4338 10670 4350 10722
rect 5506 10670 5518 10722
rect 5570 10670 5582 10722
rect 10994 10670 11006 10722
rect 11058 10670 11070 10722
rect 11330 10670 11342 10722
rect 11394 10670 11406 10722
rect 2494 10658 2546 10670
rect 20862 10658 20914 10670
rect 23102 10722 23154 10734
rect 23102 10658 23154 10670
rect 3502 10610 3554 10622
rect 11566 10610 11618 10622
rect 20974 10610 21026 10622
rect 2258 10558 2270 10610
rect 2322 10558 2334 10610
rect 3938 10558 3950 10610
rect 4002 10558 4014 10610
rect 4722 10558 4734 10610
rect 4786 10558 4798 10610
rect 17378 10558 17390 10610
rect 17442 10558 17454 10610
rect 3502 10546 3554 10558
rect 11566 10546 11618 10558
rect 20974 10546 21026 10558
rect 21646 10610 21698 10622
rect 21646 10546 21698 10558
rect 21870 10610 21922 10622
rect 22530 10558 22542 10610
rect 22594 10558 22606 10610
rect 23762 10558 23774 10610
rect 23826 10558 23838 10610
rect 21870 10546 21922 10558
rect 7634 10446 7646 10498
rect 7698 10446 7710 10498
rect 15586 10446 15598 10498
rect 15650 10446 15662 10498
rect 18162 10446 18174 10498
rect 18226 10446 18238 10498
rect 20290 10446 20302 10498
rect 20354 10446 20366 10498
rect 23538 10446 23550 10498
rect 23602 10446 23614 10498
rect 16382 10386 16434 10398
rect 16382 10322 16434 10334
rect 21086 10386 21138 10398
rect 21086 10322 21138 10334
rect 21534 10386 21586 10398
rect 21534 10322 21586 10334
rect 21982 10386 22034 10398
rect 21982 10322 22034 10334
rect 1344 10218 24640 10252
rect 1344 10166 4126 10218
rect 4178 10166 4230 10218
rect 4282 10166 4334 10218
rect 4386 10166 9950 10218
rect 10002 10166 10054 10218
rect 10106 10166 10158 10218
rect 10210 10166 15774 10218
rect 15826 10166 15878 10218
rect 15930 10166 15982 10218
rect 16034 10166 21598 10218
rect 21650 10166 21702 10218
rect 21754 10166 21806 10218
rect 21858 10166 24640 10218
rect 1344 10132 24640 10166
rect 18174 10050 18226 10062
rect 18174 9986 18226 9998
rect 2482 9886 2494 9938
rect 2546 9886 2558 9938
rect 4610 9886 4622 9938
rect 4674 9886 4686 9938
rect 12002 9886 12014 9938
rect 12066 9886 12078 9938
rect 22082 9886 22094 9938
rect 22146 9886 22158 9938
rect 24210 9886 24222 9938
rect 24274 9886 24286 9938
rect 7198 9826 7250 9838
rect 15038 9826 15090 9838
rect 1810 9774 1822 9826
rect 1874 9774 1886 9826
rect 8530 9774 8542 9826
rect 8594 9774 8606 9826
rect 9090 9774 9102 9826
rect 9154 9774 9166 9826
rect 7198 9762 7250 9774
rect 15038 9762 15090 9774
rect 15262 9826 15314 9838
rect 20078 9826 20130 9838
rect 19842 9774 19854 9826
rect 19906 9774 19918 9826
rect 15262 9762 15314 9774
rect 20078 9762 20130 9774
rect 20414 9826 20466 9838
rect 20414 9762 20466 9774
rect 20750 9826 20802 9838
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 20750 9762 20802 9774
rect 14814 9714 14866 9726
rect 9874 9662 9886 9714
rect 9938 9662 9950 9714
rect 14814 9650 14866 9662
rect 18286 9714 18338 9726
rect 18286 9650 18338 9662
rect 18510 9714 18562 9726
rect 18510 9650 18562 9662
rect 19182 9714 19234 9726
rect 19182 9650 19234 9662
rect 20638 9714 20690 9726
rect 20638 9650 20690 9662
rect 6862 9602 6914 9614
rect 6862 9538 6914 9550
rect 8766 9602 8818 9614
rect 8766 9538 8818 9550
rect 14926 9602 14978 9614
rect 14926 9538 14978 9550
rect 1344 9434 24800 9468
rect 1344 9382 7038 9434
rect 7090 9382 7142 9434
rect 7194 9382 7246 9434
rect 7298 9382 12862 9434
rect 12914 9382 12966 9434
rect 13018 9382 13070 9434
rect 13122 9382 18686 9434
rect 18738 9382 18790 9434
rect 18842 9382 18894 9434
rect 18946 9382 24510 9434
rect 24562 9382 24614 9434
rect 24666 9382 24718 9434
rect 24770 9382 24800 9434
rect 1344 9348 24800 9382
rect 4510 9266 4562 9278
rect 4510 9202 4562 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 16270 9266 16322 9278
rect 16270 9202 16322 9214
rect 16606 9266 16658 9278
rect 16606 9202 16658 9214
rect 22094 9266 22146 9278
rect 22094 9202 22146 9214
rect 22878 9154 22930 9166
rect 5394 9102 5406 9154
rect 5458 9102 5470 9154
rect 6850 9102 6862 9154
rect 6914 9102 6926 9154
rect 10658 9102 10670 9154
rect 10722 9102 10734 9154
rect 14914 9102 14926 9154
rect 14978 9102 14990 9154
rect 22878 9090 22930 9102
rect 4846 9042 4898 9054
rect 9998 9042 10050 9054
rect 16494 9042 16546 9054
rect 21086 9042 21138 9054
rect 5618 8990 5630 9042
rect 5682 8990 5694 9042
rect 6066 8990 6078 9042
rect 6130 8990 6142 9042
rect 10434 8990 10446 9042
rect 10498 8990 10510 9042
rect 15698 8990 15710 9042
rect 15762 8990 15774 9042
rect 16034 8990 16046 9042
rect 16098 8990 16110 9042
rect 17378 8990 17390 9042
rect 17442 8990 17454 9042
rect 4846 8978 4898 8990
rect 9998 8978 10050 8990
rect 16494 8978 16546 8990
rect 21086 8978 21138 8990
rect 21310 9042 21362 9054
rect 21310 8978 21362 8990
rect 21422 9042 21474 9054
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 23314 8990 23326 9042
rect 23378 8990 23390 9042
rect 21422 8978 21474 8990
rect 16382 8930 16434 8942
rect 8978 8878 8990 8930
rect 9042 8878 9054 8930
rect 12786 8878 12798 8930
rect 12850 8878 12862 8930
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 23650 8878 23662 8930
rect 23714 8878 23726 8930
rect 16382 8866 16434 8878
rect 1344 8650 24640 8684
rect 1344 8598 4126 8650
rect 4178 8598 4230 8650
rect 4282 8598 4334 8650
rect 4386 8598 9950 8650
rect 10002 8598 10054 8650
rect 10106 8598 10158 8650
rect 10210 8598 15774 8650
rect 15826 8598 15878 8650
rect 15930 8598 15982 8650
rect 16034 8598 21598 8650
rect 21650 8598 21702 8650
rect 21754 8598 21806 8650
rect 21858 8598 24640 8650
rect 1344 8564 24640 8598
rect 18174 8482 18226 8494
rect 18174 8418 18226 8430
rect 6078 8370 6130 8382
rect 4610 8318 4622 8370
rect 4674 8318 4686 8370
rect 6078 8306 6130 8318
rect 12014 8370 12066 8382
rect 12014 8306 12066 8318
rect 15374 8370 15426 8382
rect 15374 8306 15426 8318
rect 15486 8370 15538 8382
rect 15486 8306 15538 8318
rect 15822 8370 15874 8382
rect 15822 8306 15874 8318
rect 18510 8370 18562 8382
rect 24110 8370 24162 8382
rect 22082 8318 22094 8370
rect 22146 8318 22158 8370
rect 18510 8306 18562 8318
rect 24110 8306 24162 8318
rect 20078 8258 20130 8270
rect 1810 8206 1822 8258
rect 1874 8206 1886 8258
rect 6850 8206 6862 8258
rect 6914 8206 6926 8258
rect 11554 8206 11566 8258
rect 11618 8206 11630 8258
rect 13906 8206 13918 8258
rect 13970 8206 13982 8258
rect 19730 8206 19742 8258
rect 19794 8206 19806 8258
rect 23426 8206 23438 8258
rect 23490 8206 23502 8258
rect 23874 8206 23886 8258
rect 23938 8206 23950 8258
rect 20078 8194 20130 8206
rect 9438 8146 9490 8158
rect 13470 8146 13522 8158
rect 2482 8094 2494 8146
rect 2546 8094 2558 8146
rect 6626 8094 6638 8146
rect 6690 8094 6702 8146
rect 11442 8094 11454 8146
rect 11506 8094 11518 8146
rect 9438 8082 9490 8094
rect 13470 8082 13522 8094
rect 20526 8146 20578 8158
rect 20526 8082 20578 8094
rect 20750 8146 20802 8158
rect 20750 8082 20802 8094
rect 21422 8146 21474 8158
rect 21422 8082 21474 8094
rect 21534 8146 21586 8158
rect 21534 8082 21586 8094
rect 21646 8146 21698 8158
rect 21646 8082 21698 8094
rect 5742 8034 5794 8046
rect 5742 7970 5794 7982
rect 9998 8034 10050 8046
rect 9998 7970 10050 7982
rect 12350 8034 12402 8046
rect 12350 7970 12402 7982
rect 15934 8034 15986 8046
rect 15934 7970 15986 7982
rect 18286 8034 18338 8046
rect 20414 8034 20466 8046
rect 19506 7982 19518 8034
rect 19570 7982 19582 8034
rect 18286 7970 18338 7982
rect 20414 7970 20466 7982
rect 22878 8034 22930 8046
rect 22878 7970 22930 7982
rect 1344 7866 24800 7900
rect 1344 7814 7038 7866
rect 7090 7814 7142 7866
rect 7194 7814 7246 7866
rect 7298 7814 12862 7866
rect 12914 7814 12966 7866
rect 13018 7814 13070 7866
rect 13122 7814 18686 7866
rect 18738 7814 18790 7866
rect 18842 7814 18894 7866
rect 18946 7814 24510 7866
rect 24562 7814 24614 7866
rect 24666 7814 24718 7866
rect 24770 7814 24800 7866
rect 1344 7780 24800 7814
rect 2494 7698 2546 7710
rect 2494 7634 2546 7646
rect 19742 7698 19794 7710
rect 19742 7634 19794 7646
rect 22878 7698 22930 7710
rect 22878 7634 22930 7646
rect 23886 7698 23938 7710
rect 23886 7634 23938 7646
rect 7198 7586 7250 7598
rect 22318 7586 22370 7598
rect 4386 7534 4398 7586
rect 4450 7534 4462 7586
rect 6514 7534 6526 7586
rect 6578 7534 6590 7586
rect 8306 7534 8318 7586
rect 8370 7534 8382 7586
rect 11106 7534 11118 7586
rect 11170 7534 11182 7586
rect 12562 7534 12574 7586
rect 12626 7534 12638 7586
rect 16034 7534 16046 7586
rect 16098 7534 16110 7586
rect 7198 7522 7250 7534
rect 22318 7522 22370 7534
rect 23550 7586 23602 7598
rect 23550 7522 23602 7534
rect 24222 7586 24274 7598
rect 24222 7522 24274 7534
rect 3278 7474 3330 7486
rect 2258 7422 2270 7474
rect 2322 7422 2334 7474
rect 2706 7422 2718 7474
rect 2770 7471 2782 7474
rect 3042 7471 3054 7474
rect 2770 7425 3054 7471
rect 2770 7422 2782 7425
rect 3042 7422 3054 7425
rect 3106 7422 3118 7474
rect 3278 7410 3330 7422
rect 3614 7474 3666 7486
rect 5854 7474 5906 7486
rect 7534 7474 7586 7486
rect 10334 7474 10386 7486
rect 12014 7474 12066 7486
rect 18958 7474 19010 7486
rect 4162 7422 4174 7474
rect 4226 7422 4238 7474
rect 6290 7422 6302 7474
rect 6354 7422 6366 7474
rect 8194 7422 8206 7474
rect 8258 7422 8270 7474
rect 10882 7422 10894 7474
rect 10946 7422 10958 7474
rect 12786 7422 12798 7474
rect 12850 7422 12862 7474
rect 16818 7422 16830 7474
rect 16882 7422 16894 7474
rect 18274 7422 18286 7474
rect 18338 7422 18350 7474
rect 3614 7410 3666 7422
rect 5854 7410 5906 7422
rect 7534 7410 7586 7422
rect 10334 7410 10386 7422
rect 12014 7410 12066 7422
rect 18958 7410 19010 7422
rect 19182 7474 19234 7486
rect 19182 7410 19234 7422
rect 19518 7474 19570 7486
rect 19518 7410 19570 7422
rect 21310 7474 21362 7486
rect 21310 7410 21362 7422
rect 21422 7474 21474 7486
rect 21422 7410 21474 7422
rect 21646 7474 21698 7486
rect 22642 7422 22654 7474
rect 22706 7422 22718 7474
rect 23314 7422 23326 7474
rect 23378 7422 23390 7474
rect 21646 7410 21698 7422
rect 19630 7362 19682 7374
rect 13906 7310 13918 7362
rect 13970 7310 13982 7362
rect 19630 7298 19682 7310
rect 5518 7250 5570 7262
rect 5518 7186 5570 7198
rect 9998 7250 10050 7262
rect 9998 7186 10050 7198
rect 11678 7250 11730 7262
rect 11678 7186 11730 7198
rect 21758 7250 21810 7262
rect 21758 7186 21810 7198
rect 1344 7082 24640 7116
rect 1344 7030 4126 7082
rect 4178 7030 4230 7082
rect 4282 7030 4334 7082
rect 4386 7030 9950 7082
rect 10002 7030 10054 7082
rect 10106 7030 10158 7082
rect 10210 7030 15774 7082
rect 15826 7030 15878 7082
rect 15930 7030 15982 7082
rect 16034 7030 21598 7082
rect 21650 7030 21702 7082
rect 21754 7030 21806 7082
rect 21858 7030 24640 7082
rect 1344 6996 24640 7030
rect 9102 6914 9154 6926
rect 9102 6850 9154 6862
rect 18498 6750 18510 6802
rect 18562 6750 18574 6802
rect 20626 6750 20638 6802
rect 20690 6750 20702 6802
rect 24210 6750 24222 6802
rect 24274 6750 24286 6802
rect 4510 6690 4562 6702
rect 9650 6638 9662 6690
rect 9714 6638 9726 6690
rect 11778 6638 11790 6690
rect 11842 6638 11854 6690
rect 17714 6638 17726 6690
rect 17778 6638 17790 6690
rect 21298 6638 21310 6690
rect 21362 6638 21374 6690
rect 22082 6638 22094 6690
rect 22146 6638 22158 6690
rect 4510 6626 4562 6638
rect 8094 6578 8146 6590
rect 8094 6514 8146 6526
rect 8766 6578 8818 6590
rect 9762 6526 9774 6578
rect 9826 6526 9838 6578
rect 8766 6514 8818 6526
rect 4174 6466 4226 6478
rect 4174 6402 4226 6414
rect 7758 6466 7810 6478
rect 7758 6402 7810 6414
rect 12014 6466 12066 6478
rect 12014 6402 12066 6414
rect 1344 6298 24800 6332
rect 1344 6246 7038 6298
rect 7090 6246 7142 6298
rect 7194 6246 7246 6298
rect 7298 6246 12862 6298
rect 12914 6246 12966 6298
rect 13018 6246 13070 6298
rect 13122 6246 18686 6298
rect 18738 6246 18790 6298
rect 18842 6246 18894 6298
rect 18946 6246 24510 6298
rect 24562 6246 24614 6298
rect 24666 6246 24718 6298
rect 24770 6246 24800 6298
rect 1344 6212 24800 6246
rect 20638 6130 20690 6142
rect 20638 6066 20690 6078
rect 22878 6130 22930 6142
rect 22878 6066 22930 6078
rect 3602 5966 3614 6018
rect 3666 5966 3678 6018
rect 6850 5966 6862 6018
rect 6914 5966 6926 6018
rect 13458 5966 13470 6018
rect 13522 5966 13534 6018
rect 20974 5906 21026 5918
rect 2930 5854 2942 5906
rect 2994 5854 3006 5906
rect 6178 5854 6190 5906
rect 6242 5854 6254 5906
rect 14242 5854 14254 5906
rect 14306 5854 14318 5906
rect 20974 5842 21026 5854
rect 23102 5906 23154 5918
rect 23998 5906 24050 5918
rect 23538 5854 23550 5906
rect 23602 5854 23614 5906
rect 23102 5842 23154 5854
rect 23998 5842 24050 5854
rect 5730 5742 5742 5794
rect 5794 5742 5806 5794
rect 8978 5742 8990 5794
rect 9042 5742 9054 5794
rect 11330 5742 11342 5794
rect 11394 5742 11406 5794
rect 1344 5514 24640 5548
rect 1344 5462 4126 5514
rect 4178 5462 4230 5514
rect 4282 5462 4334 5514
rect 4386 5462 9950 5514
rect 10002 5462 10054 5514
rect 10106 5462 10158 5514
rect 10210 5462 15774 5514
rect 15826 5462 15878 5514
rect 15930 5462 15982 5514
rect 16034 5462 21598 5514
rect 21650 5462 21702 5514
rect 21754 5462 21806 5514
rect 21858 5462 24640 5514
rect 1344 5428 24640 5462
rect 23102 5234 23154 5246
rect 23538 5182 23550 5234
rect 23602 5182 23614 5234
rect 23102 5170 23154 5182
rect 23762 5070 23774 5122
rect 23826 5070 23838 5122
rect 1344 4730 24800 4764
rect 1344 4678 7038 4730
rect 7090 4678 7142 4730
rect 7194 4678 7246 4730
rect 7298 4678 12862 4730
rect 12914 4678 12966 4730
rect 13018 4678 13070 4730
rect 13122 4678 18686 4730
rect 18738 4678 18790 4730
rect 18842 4678 18894 4730
rect 18946 4678 24510 4730
rect 24562 4678 24614 4730
rect 24666 4678 24718 4730
rect 24770 4678 24800 4730
rect 1344 4644 24800 4678
rect 23886 4562 23938 4574
rect 23886 4498 23938 4510
rect 24222 4338 24274 4350
rect 24222 4274 24274 4286
rect 23662 4226 23714 4238
rect 23662 4162 23714 4174
rect 1344 3946 24640 3980
rect 1344 3894 4126 3946
rect 4178 3894 4230 3946
rect 4282 3894 4334 3946
rect 4386 3894 9950 3946
rect 10002 3894 10054 3946
rect 10106 3894 10158 3946
rect 10210 3894 15774 3946
rect 15826 3894 15878 3946
rect 15930 3894 15982 3946
rect 16034 3894 21598 3946
rect 21650 3894 21702 3946
rect 21754 3894 21806 3946
rect 21858 3894 24640 3946
rect 1344 3860 24640 3894
rect 23438 3442 23490 3454
rect 23438 3378 23490 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 1344 3162 24800 3196
rect 1344 3110 7038 3162
rect 7090 3110 7142 3162
rect 7194 3110 7246 3162
rect 7298 3110 12862 3162
rect 12914 3110 12966 3162
rect 13018 3110 13070 3162
rect 13122 3110 18686 3162
rect 18738 3110 18790 3162
rect 18842 3110 18894 3162
rect 18946 3110 24510 3162
rect 24562 3110 24614 3162
rect 24666 3110 24718 3162
rect 24770 3110 24800 3162
rect 1344 3076 24800 3110
<< via1 >>
rect 4126 22710 4178 22762
rect 4230 22710 4282 22762
rect 4334 22710 4386 22762
rect 9950 22710 10002 22762
rect 10054 22710 10106 22762
rect 10158 22710 10210 22762
rect 15774 22710 15826 22762
rect 15878 22710 15930 22762
rect 15982 22710 16034 22762
rect 21598 22710 21650 22762
rect 21702 22710 21754 22762
rect 21806 22710 21858 22762
rect 22430 22542 22482 22594
rect 12686 22430 12738 22482
rect 13134 22318 13186 22370
rect 19630 22318 19682 22370
rect 19966 22318 20018 22370
rect 20862 22318 20914 22370
rect 21422 22318 21474 22370
rect 13470 22094 13522 22146
rect 20190 22094 20242 22146
rect 21086 22094 21138 22146
rect 7038 21926 7090 21978
rect 7142 21926 7194 21978
rect 7246 21926 7298 21978
rect 12862 21926 12914 21978
rect 12966 21926 13018 21978
rect 13070 21926 13122 21978
rect 18686 21926 18738 21978
rect 18790 21926 18842 21978
rect 18894 21926 18946 21978
rect 24510 21926 24562 21978
rect 24614 21926 24666 21978
rect 24718 21926 24770 21978
rect 8542 21646 8594 21698
rect 5070 21534 5122 21586
rect 8318 21534 8370 21586
rect 9886 21534 9938 21586
rect 13246 21534 13298 21586
rect 17838 21534 17890 21586
rect 21086 21534 21138 21586
rect 5742 21422 5794 21474
rect 7870 21422 7922 21474
rect 10670 21422 10722 21474
rect 12798 21422 12850 21474
rect 13918 21422 13970 21474
rect 16046 21422 16098 21474
rect 18622 21422 18674 21474
rect 20750 21422 20802 21474
rect 21870 21422 21922 21474
rect 23998 21422 24050 21474
rect 4126 21142 4178 21194
rect 4230 21142 4282 21194
rect 4334 21142 4386 21194
rect 9950 21142 10002 21194
rect 10054 21142 10106 21194
rect 10158 21142 10210 21194
rect 15774 21142 15826 21194
rect 15878 21142 15930 21194
rect 15982 21142 16034 21194
rect 21598 21142 21650 21194
rect 21702 21142 21754 21194
rect 21806 21142 21858 21194
rect 9102 20974 9154 21026
rect 10222 20974 10274 21026
rect 21198 20974 21250 21026
rect 21534 20974 21586 21026
rect 18398 20862 18450 20914
rect 21534 20862 21586 20914
rect 23998 20862 24050 20914
rect 7982 20750 8034 20802
rect 8430 20750 8482 20802
rect 8878 20750 8930 20802
rect 9550 20750 9602 20802
rect 10110 20750 10162 20802
rect 10670 20750 10722 20802
rect 15598 20750 15650 20802
rect 19294 20750 19346 20802
rect 19742 20750 19794 20802
rect 22094 20750 22146 20802
rect 22542 20750 22594 20802
rect 23662 20750 23714 20802
rect 7870 20638 7922 20690
rect 8542 20638 8594 20690
rect 10222 20638 10274 20690
rect 10782 20638 10834 20690
rect 16270 20638 16322 20690
rect 20190 20638 20242 20690
rect 21870 20638 21922 20690
rect 23214 20638 23266 20690
rect 7038 20358 7090 20410
rect 7142 20358 7194 20410
rect 7246 20358 7298 20410
rect 12862 20358 12914 20410
rect 12966 20358 13018 20410
rect 13070 20358 13122 20410
rect 18686 20358 18738 20410
rect 18790 20358 18842 20410
rect 18894 20358 18946 20410
rect 24510 20358 24562 20410
rect 24614 20358 24666 20410
rect 24718 20358 24770 20410
rect 8766 20190 8818 20242
rect 14030 20190 14082 20242
rect 17502 20190 17554 20242
rect 6974 20078 7026 20130
rect 9550 20078 9602 20130
rect 9998 20078 10050 20130
rect 14254 20078 14306 20130
rect 14926 20078 14978 20130
rect 16494 20078 16546 20130
rect 16606 20078 16658 20130
rect 17726 20078 17778 20130
rect 19630 20078 19682 20130
rect 19854 20078 19906 20130
rect 20302 20078 20354 20130
rect 21198 20078 21250 20130
rect 21310 20078 21362 20130
rect 21422 20078 21474 20130
rect 21982 20078 22034 20130
rect 22206 20078 22258 20130
rect 3502 19966 3554 20018
rect 4174 19966 4226 20018
rect 7982 19966 8034 20018
rect 8654 19966 8706 20018
rect 9774 19966 9826 20018
rect 13918 19966 13970 20018
rect 14366 19966 14418 20018
rect 15150 19966 15202 20018
rect 16046 19966 16098 20018
rect 16830 19966 16882 20018
rect 17390 19966 17442 20018
rect 20078 19966 20130 20018
rect 20414 19966 20466 20018
rect 21758 19966 21810 20018
rect 23214 19966 23266 20018
rect 23550 19966 23602 20018
rect 6302 19854 6354 19906
rect 6862 19854 6914 19906
rect 7310 19854 7362 19906
rect 8206 19854 8258 19906
rect 16494 19854 16546 19906
rect 19518 19854 19570 19906
rect 22094 19854 22146 19906
rect 22878 19854 22930 19906
rect 24110 19854 24162 19906
rect 8766 19742 8818 19794
rect 9886 19742 9938 19794
rect 4126 19574 4178 19626
rect 4230 19574 4282 19626
rect 4334 19574 4386 19626
rect 9950 19574 10002 19626
rect 10054 19574 10106 19626
rect 10158 19574 10210 19626
rect 15774 19574 15826 19626
rect 15878 19574 15930 19626
rect 15982 19574 16034 19626
rect 21598 19574 21650 19626
rect 21702 19574 21754 19626
rect 21806 19574 21858 19626
rect 4958 19406 5010 19458
rect 12014 19406 12066 19458
rect 4622 19294 4674 19346
rect 10334 19294 10386 19346
rect 14366 19294 14418 19346
rect 20302 19294 20354 19346
rect 21646 19294 21698 19346
rect 1822 19182 1874 19234
rect 7982 19182 8034 19234
rect 8206 19182 8258 19234
rect 8318 19182 8370 19234
rect 10558 19182 10610 19234
rect 11230 19182 11282 19234
rect 12014 19182 12066 19234
rect 12462 19182 12514 19234
rect 12686 19182 12738 19234
rect 14254 19182 14306 19234
rect 14926 19182 14978 19234
rect 15038 19182 15090 19234
rect 15262 19182 15314 19234
rect 15598 19182 15650 19234
rect 16046 19182 16098 19234
rect 17166 19182 17218 19234
rect 17502 19182 17554 19234
rect 21982 19182 22034 19234
rect 22542 19182 22594 19234
rect 22654 19182 22706 19234
rect 22990 19182 23042 19234
rect 2494 19070 2546 19122
rect 5070 19070 5122 19122
rect 9102 19070 9154 19122
rect 9214 19070 9266 19122
rect 11902 19070 11954 19122
rect 13806 19070 13858 19122
rect 14478 19070 14530 19122
rect 15486 19070 15538 19122
rect 18174 19070 18226 19122
rect 24222 19070 24274 19122
rect 7758 18958 7810 19010
rect 8766 18958 8818 19010
rect 9438 18958 9490 19010
rect 10110 18958 10162 19010
rect 10894 18958 10946 19010
rect 11342 18958 11394 19010
rect 11566 18958 11618 19010
rect 13918 18958 13970 19010
rect 16158 18958 16210 19010
rect 16494 18958 16546 19010
rect 16606 18958 16658 19010
rect 16830 18958 16882 19010
rect 22206 18958 22258 19010
rect 23886 18958 23938 19010
rect 7038 18790 7090 18842
rect 7142 18790 7194 18842
rect 7246 18790 7298 18842
rect 12862 18790 12914 18842
rect 12966 18790 13018 18842
rect 13070 18790 13122 18842
rect 18686 18790 18738 18842
rect 18790 18790 18842 18842
rect 18894 18790 18946 18842
rect 24510 18790 24562 18842
rect 24614 18790 24666 18842
rect 24718 18790 24770 18842
rect 8206 18622 8258 18674
rect 8430 18622 8482 18674
rect 8990 18622 9042 18674
rect 11566 18622 11618 18674
rect 13358 18622 13410 18674
rect 14814 18622 14866 18674
rect 15486 18622 15538 18674
rect 18174 18622 18226 18674
rect 20190 18622 20242 18674
rect 3390 18510 3442 18562
rect 5630 18510 5682 18562
rect 6190 18510 6242 18562
rect 7086 18510 7138 18562
rect 8094 18510 8146 18562
rect 8654 18510 8706 18562
rect 10446 18510 10498 18562
rect 11342 18510 11394 18562
rect 11790 18510 11842 18562
rect 12686 18510 12738 18562
rect 13694 18510 13746 18562
rect 17390 18510 17442 18562
rect 19742 18510 19794 18562
rect 3614 18398 3666 18450
rect 3950 18398 4002 18450
rect 4398 18398 4450 18450
rect 4846 18398 4898 18450
rect 5518 18398 5570 18450
rect 7310 18398 7362 18450
rect 9774 18398 9826 18450
rect 10782 18398 10834 18450
rect 11006 18398 11058 18450
rect 12238 18398 12290 18450
rect 12910 18398 12962 18450
rect 14702 18398 14754 18450
rect 15710 18398 15762 18450
rect 17614 18398 17666 18450
rect 18062 18398 18114 18450
rect 18398 18398 18450 18450
rect 19518 18398 19570 18450
rect 20974 18398 21026 18450
rect 9550 18286 9602 18338
rect 10558 18286 10610 18338
rect 14926 18286 14978 18338
rect 20078 18286 20130 18338
rect 21758 18286 21810 18338
rect 23886 18286 23938 18338
rect 3278 18174 3330 18226
rect 4062 18174 4114 18226
rect 6526 18174 6578 18226
rect 10110 18174 10162 18226
rect 11454 18174 11506 18226
rect 12126 18174 12178 18226
rect 14366 18174 14418 18226
rect 14478 18174 14530 18226
rect 15374 18174 15426 18226
rect 20414 18174 20466 18226
rect 4126 18006 4178 18058
rect 4230 18006 4282 18058
rect 4334 18006 4386 18058
rect 9950 18006 10002 18058
rect 10054 18006 10106 18058
rect 10158 18006 10210 18058
rect 15774 18006 15826 18058
rect 15878 18006 15930 18058
rect 15982 18006 16034 18058
rect 21598 18006 21650 18058
rect 21702 18006 21754 18058
rect 21806 18006 21858 18058
rect 2942 17838 2994 17890
rect 3614 17838 3666 17890
rect 4622 17838 4674 17890
rect 14254 17838 14306 17890
rect 16494 17838 16546 17890
rect 21310 17838 21362 17890
rect 22206 17838 22258 17890
rect 22318 17838 22370 17890
rect 22654 17838 22706 17890
rect 3838 17726 3890 17778
rect 6302 17726 6354 17778
rect 7198 17726 7250 17778
rect 8878 17726 8930 17778
rect 20302 17726 20354 17778
rect 2382 17614 2434 17666
rect 2830 17614 2882 17666
rect 4734 17614 4786 17666
rect 5742 17614 5794 17666
rect 6750 17614 6802 17666
rect 12686 17614 12738 17666
rect 14142 17614 14194 17666
rect 16158 17614 16210 17666
rect 17502 17614 17554 17666
rect 21646 17614 21698 17666
rect 21870 17614 21922 17666
rect 22542 17614 22594 17666
rect 23214 17614 23266 17666
rect 23774 17614 23826 17666
rect 4622 17502 4674 17554
rect 15934 17502 15986 17554
rect 16830 17502 16882 17554
rect 18174 17502 18226 17554
rect 23102 17502 23154 17554
rect 2158 17390 2210 17442
rect 3278 17390 3330 17442
rect 5966 17390 6018 17442
rect 14254 17390 14306 17442
rect 16942 17390 16994 17442
rect 17166 17390 17218 17442
rect 7038 17222 7090 17274
rect 7142 17222 7194 17274
rect 7246 17222 7298 17274
rect 12862 17222 12914 17274
rect 12966 17222 13018 17274
rect 13070 17222 13122 17274
rect 18686 17222 18738 17274
rect 18790 17222 18842 17274
rect 18894 17222 18946 17274
rect 24510 17222 24562 17274
rect 24614 17222 24666 17274
rect 24718 17222 24770 17274
rect 5966 17054 6018 17106
rect 6302 17054 6354 17106
rect 5182 16942 5234 16994
rect 5630 16942 5682 16994
rect 7310 16942 7362 16994
rect 8542 16942 8594 16994
rect 14142 16942 14194 16994
rect 16270 16942 16322 16994
rect 20974 16942 21026 16994
rect 6638 16830 6690 16882
rect 7646 16830 7698 16882
rect 8094 16830 8146 16882
rect 9438 16830 9490 16882
rect 10110 16830 10162 16882
rect 10334 16830 10386 16882
rect 10894 16830 10946 16882
rect 16606 16830 16658 16882
rect 17390 16830 17442 16882
rect 22878 16830 22930 16882
rect 23102 16830 23154 16882
rect 23438 16830 23490 16882
rect 23550 16830 23602 16882
rect 9886 16718 9938 16770
rect 11678 16718 11730 16770
rect 13806 16718 13858 16770
rect 5294 16606 5346 16658
rect 7982 16606 8034 16658
rect 14254 16606 14306 16658
rect 23998 16606 24050 16658
rect 4126 16438 4178 16490
rect 4230 16438 4282 16490
rect 4334 16438 4386 16490
rect 9950 16438 10002 16490
rect 10054 16438 10106 16490
rect 10158 16438 10210 16490
rect 15774 16438 15826 16490
rect 15878 16438 15930 16490
rect 15982 16438 16034 16490
rect 21598 16438 21650 16490
rect 21702 16438 21754 16490
rect 21806 16438 21858 16490
rect 2830 16270 2882 16322
rect 21310 16270 21362 16322
rect 10222 16158 10274 16210
rect 12686 16158 12738 16210
rect 23438 16158 23490 16210
rect 4846 16046 4898 16098
rect 5854 16046 5906 16098
rect 6078 16046 6130 16098
rect 7422 16046 7474 16098
rect 11566 16046 11618 16098
rect 11902 16046 11954 16098
rect 14590 16046 14642 16098
rect 16718 16046 16770 16098
rect 19070 16046 19122 16098
rect 21646 16046 21698 16098
rect 21870 16046 21922 16098
rect 23214 16046 23266 16098
rect 24222 16046 24274 16098
rect 3166 15934 3218 15986
rect 3614 15934 3666 15986
rect 4062 15934 4114 15986
rect 4286 15934 4338 15986
rect 4398 15934 4450 15986
rect 8094 15934 8146 15986
rect 11230 15934 11282 15986
rect 12126 15934 12178 15986
rect 12238 15934 12290 15986
rect 14702 15934 14754 15986
rect 17726 15934 17778 15986
rect 22542 15934 22594 15986
rect 24110 15934 24162 15986
rect 2494 15822 2546 15874
rect 4174 15822 4226 15874
rect 6302 15822 6354 15874
rect 6414 15822 6466 15874
rect 18286 15822 18338 15874
rect 18734 15822 18786 15874
rect 7038 15654 7090 15706
rect 7142 15654 7194 15706
rect 7246 15654 7298 15706
rect 12862 15654 12914 15706
rect 12966 15654 13018 15706
rect 13070 15654 13122 15706
rect 18686 15654 18738 15706
rect 18790 15654 18842 15706
rect 18894 15654 18946 15706
rect 24510 15654 24562 15706
rect 24614 15654 24666 15706
rect 24718 15654 24770 15706
rect 2942 15486 2994 15538
rect 5966 15486 6018 15538
rect 8094 15486 8146 15538
rect 8542 15486 8594 15538
rect 13022 15486 13074 15538
rect 16494 15486 16546 15538
rect 18510 15486 18562 15538
rect 21422 15486 21474 15538
rect 2046 15374 2098 15426
rect 2270 15374 2322 15426
rect 2830 15374 2882 15426
rect 3838 15374 3890 15426
rect 5294 15374 5346 15426
rect 5854 15374 5906 15426
rect 7422 15374 7474 15426
rect 8654 15374 8706 15426
rect 13806 15374 13858 15426
rect 14142 15374 14194 15426
rect 16158 15374 16210 15426
rect 17614 15374 17666 15426
rect 18846 15374 18898 15426
rect 19518 15374 19570 15426
rect 21534 15374 21586 15426
rect 22990 15374 23042 15426
rect 2606 15262 2658 15314
rect 3390 15262 3442 15314
rect 4398 15262 4450 15314
rect 4734 15262 4786 15314
rect 6414 15262 6466 15314
rect 6750 15262 6802 15314
rect 7870 15262 7922 15314
rect 13134 15262 13186 15314
rect 13358 15262 13410 15314
rect 13470 15262 13522 15314
rect 14254 15262 14306 15314
rect 14590 15262 14642 15314
rect 15598 15262 15650 15314
rect 15822 15262 15874 15314
rect 17390 15262 17442 15314
rect 17726 15262 17778 15314
rect 19630 15262 19682 15314
rect 19854 15262 19906 15314
rect 20414 15262 20466 15314
rect 24110 15262 24162 15314
rect 2158 15150 2210 15202
rect 4846 15150 4898 15202
rect 15486 15150 15538 15202
rect 3054 15038 3106 15090
rect 8542 15038 8594 15090
rect 18174 15038 18226 15090
rect 19966 15038 20018 15090
rect 4126 14870 4178 14922
rect 4230 14870 4282 14922
rect 4334 14870 4386 14922
rect 9950 14870 10002 14922
rect 10054 14870 10106 14922
rect 10158 14870 10210 14922
rect 15774 14870 15826 14922
rect 15878 14870 15930 14922
rect 15982 14870 16034 14922
rect 21598 14870 21650 14922
rect 21702 14870 21754 14922
rect 21806 14870 21858 14922
rect 2270 14702 2322 14754
rect 12910 14702 12962 14754
rect 20078 14702 20130 14754
rect 20414 14702 20466 14754
rect 20750 14702 20802 14754
rect 22094 14702 22146 14754
rect 2830 14590 2882 14642
rect 6302 14590 6354 14642
rect 7870 14590 7922 14642
rect 12014 14590 12066 14642
rect 12798 14590 12850 14642
rect 17166 14590 17218 14642
rect 19966 14590 20018 14642
rect 22654 14590 22706 14642
rect 23550 14590 23602 14642
rect 2606 14478 2658 14530
rect 3278 14478 3330 14530
rect 3614 14478 3666 14530
rect 4174 14478 4226 14530
rect 4622 14478 4674 14530
rect 4846 14478 4898 14530
rect 6526 14478 6578 14530
rect 8094 14478 8146 14530
rect 9214 14478 9266 14530
rect 12574 14478 12626 14530
rect 13470 14478 13522 14530
rect 19294 14478 19346 14530
rect 22318 14478 22370 14530
rect 23102 14478 23154 14530
rect 2718 14366 2770 14418
rect 3502 14366 3554 14418
rect 7198 14366 7250 14418
rect 9886 14366 9938 14418
rect 19854 14366 19906 14418
rect 20638 14366 20690 14418
rect 21758 14366 21810 14418
rect 23886 14366 23938 14418
rect 24222 14366 24274 14418
rect 2942 14254 2994 14306
rect 4398 14254 4450 14306
rect 8430 14254 8482 14306
rect 19070 14254 19122 14306
rect 21534 14254 21586 14306
rect 21982 14254 22034 14306
rect 7038 14086 7090 14138
rect 7142 14086 7194 14138
rect 7246 14086 7298 14138
rect 12862 14086 12914 14138
rect 12966 14086 13018 14138
rect 13070 14086 13122 14138
rect 18686 14086 18738 14138
rect 18790 14086 18842 14138
rect 18894 14086 18946 14138
rect 24510 14086 24562 14138
rect 24614 14086 24666 14138
rect 24718 14086 24770 14138
rect 5966 13918 6018 13970
rect 9886 13918 9938 13970
rect 14702 13918 14754 13970
rect 16494 13918 16546 13970
rect 2494 13806 2546 13858
rect 4958 13806 5010 13858
rect 12126 13806 12178 13858
rect 15374 13806 15426 13858
rect 18174 13806 18226 13858
rect 23886 13806 23938 13858
rect 24222 13806 24274 13858
rect 1822 13694 1874 13746
rect 5182 13694 5234 13746
rect 6078 13694 6130 13746
rect 6302 13694 6354 13746
rect 9550 13694 9602 13746
rect 11342 13694 11394 13746
rect 14926 13694 14978 13746
rect 15598 13694 15650 13746
rect 17502 13694 17554 13746
rect 20638 13694 20690 13746
rect 4622 13582 4674 13634
rect 14254 13582 14306 13634
rect 16382 13582 16434 13634
rect 20302 13582 20354 13634
rect 21422 13582 21474 13634
rect 23550 13582 23602 13634
rect 5518 13470 5570 13522
rect 5966 13470 6018 13522
rect 14590 13470 14642 13522
rect 15934 13470 15986 13522
rect 4126 13302 4178 13354
rect 4230 13302 4282 13354
rect 4334 13302 4386 13354
rect 9950 13302 10002 13354
rect 10054 13302 10106 13354
rect 10158 13302 10210 13354
rect 15774 13302 15826 13354
rect 15878 13302 15930 13354
rect 15982 13302 16034 13354
rect 21598 13302 21650 13354
rect 21702 13302 21754 13354
rect 21806 13302 21858 13354
rect 3054 13134 3106 13186
rect 20862 13134 20914 13186
rect 8654 13022 8706 13074
rect 10782 13022 10834 13074
rect 14030 13022 14082 13074
rect 14366 13022 14418 13074
rect 19406 13022 19458 13074
rect 22430 13022 22482 13074
rect 23326 13022 23378 13074
rect 3390 12910 3442 12962
rect 4958 12910 5010 12962
rect 6190 12910 6242 12962
rect 7870 12910 7922 12962
rect 13582 12910 13634 12962
rect 17278 12910 17330 12962
rect 19182 12910 19234 12962
rect 19854 12910 19906 12962
rect 20526 12910 20578 12962
rect 23102 12910 23154 12962
rect 12574 12798 12626 12850
rect 16494 12798 16546 12850
rect 18958 12798 19010 12850
rect 19518 12798 19570 12850
rect 19966 12798 20018 12850
rect 20302 12798 20354 12850
rect 21870 12798 21922 12850
rect 24222 12798 24274 12850
rect 3166 12686 3218 12738
rect 4734 12686 4786 12738
rect 6526 12686 6578 12738
rect 12238 12686 12290 12738
rect 21310 12686 21362 12738
rect 21422 12686 21474 12738
rect 21646 12686 21698 12738
rect 23886 12686 23938 12738
rect 7038 12518 7090 12570
rect 7142 12518 7194 12570
rect 7246 12518 7298 12570
rect 12862 12518 12914 12570
rect 12966 12518 13018 12570
rect 13070 12518 13122 12570
rect 18686 12518 18738 12570
rect 18790 12518 18842 12570
rect 18894 12518 18946 12570
rect 24510 12518 24562 12570
rect 24614 12518 24666 12570
rect 24718 12518 24770 12570
rect 15598 12350 15650 12402
rect 16158 12350 16210 12402
rect 16494 12350 16546 12402
rect 17390 12350 17442 12402
rect 21982 12350 22034 12402
rect 2718 12238 2770 12290
rect 6638 12238 6690 12290
rect 9774 12238 9826 12290
rect 12014 12238 12066 12290
rect 18398 12238 18450 12290
rect 19742 12238 19794 12290
rect 21646 12238 21698 12290
rect 23662 12238 23714 12290
rect 1934 12126 1986 12178
rect 5854 12126 5906 12178
rect 9998 12126 10050 12178
rect 11230 12126 11282 12178
rect 15150 12126 15202 12178
rect 15374 12126 15426 12178
rect 15710 12126 15762 12178
rect 18958 12126 19010 12178
rect 20078 12126 20130 12178
rect 22206 12126 22258 12178
rect 22654 12126 22706 12178
rect 4846 12014 4898 12066
rect 8766 12014 8818 12066
rect 10446 12014 10498 12066
rect 14142 12014 14194 12066
rect 15486 12014 15538 12066
rect 17502 12014 17554 12066
rect 19294 12014 19346 12066
rect 10782 11902 10834 11954
rect 4126 11734 4178 11786
rect 4230 11734 4282 11786
rect 4334 11734 4386 11786
rect 9950 11734 10002 11786
rect 10054 11734 10106 11786
rect 10158 11734 10210 11786
rect 15774 11734 15826 11786
rect 15878 11734 15930 11786
rect 15982 11734 16034 11786
rect 21598 11734 21650 11786
rect 21702 11734 21754 11786
rect 21806 11734 21858 11786
rect 13582 11566 13634 11618
rect 13918 11566 13970 11618
rect 6750 11454 6802 11506
rect 21310 11454 21362 11506
rect 23662 11454 23714 11506
rect 24334 11454 24386 11506
rect 11566 11342 11618 11394
rect 14702 11342 14754 11394
rect 16942 11342 16994 11394
rect 21422 11342 21474 11394
rect 21982 11342 22034 11394
rect 22766 11342 22818 11394
rect 23102 11342 23154 11394
rect 14478 11230 14530 11282
rect 17502 11230 17554 11282
rect 7038 10950 7090 11002
rect 7142 10950 7194 11002
rect 7246 10950 7298 11002
rect 12862 10950 12914 11002
rect 12966 10950 13018 11002
rect 13070 10950 13122 11002
rect 18686 10950 18738 11002
rect 18790 10950 18842 11002
rect 18894 10950 18946 11002
rect 24510 10950 24562 11002
rect 24614 10950 24666 11002
rect 24718 10950 24770 11002
rect 3166 10782 3218 10834
rect 11902 10782 11954 10834
rect 16046 10782 16098 10834
rect 16494 10782 16546 10834
rect 16606 10782 16658 10834
rect 22318 10782 22370 10834
rect 2494 10670 2546 10722
rect 4286 10670 4338 10722
rect 5518 10670 5570 10722
rect 11006 10670 11058 10722
rect 11342 10670 11394 10722
rect 20862 10670 20914 10722
rect 23102 10670 23154 10722
rect 2270 10558 2322 10610
rect 3502 10558 3554 10610
rect 3950 10558 4002 10610
rect 4734 10558 4786 10610
rect 11566 10558 11618 10610
rect 17390 10558 17442 10610
rect 20974 10558 21026 10610
rect 21646 10558 21698 10610
rect 21870 10558 21922 10610
rect 22542 10558 22594 10610
rect 23774 10558 23826 10610
rect 7646 10446 7698 10498
rect 15598 10446 15650 10498
rect 18174 10446 18226 10498
rect 20302 10446 20354 10498
rect 23550 10446 23602 10498
rect 16382 10334 16434 10386
rect 21086 10334 21138 10386
rect 21534 10334 21586 10386
rect 21982 10334 22034 10386
rect 4126 10166 4178 10218
rect 4230 10166 4282 10218
rect 4334 10166 4386 10218
rect 9950 10166 10002 10218
rect 10054 10166 10106 10218
rect 10158 10166 10210 10218
rect 15774 10166 15826 10218
rect 15878 10166 15930 10218
rect 15982 10166 16034 10218
rect 21598 10166 21650 10218
rect 21702 10166 21754 10218
rect 21806 10166 21858 10218
rect 18174 9998 18226 10050
rect 2494 9886 2546 9938
rect 4622 9886 4674 9938
rect 12014 9886 12066 9938
rect 22094 9886 22146 9938
rect 24222 9886 24274 9938
rect 1822 9774 1874 9826
rect 7198 9774 7250 9826
rect 8542 9774 8594 9826
rect 9102 9774 9154 9826
rect 15038 9774 15090 9826
rect 15262 9774 15314 9826
rect 19854 9774 19906 9826
rect 20078 9774 20130 9826
rect 20414 9774 20466 9826
rect 20750 9774 20802 9826
rect 21310 9774 21362 9826
rect 9886 9662 9938 9714
rect 14814 9662 14866 9714
rect 18286 9662 18338 9714
rect 18510 9662 18562 9714
rect 19182 9662 19234 9714
rect 20638 9662 20690 9714
rect 6862 9550 6914 9602
rect 8766 9550 8818 9602
rect 14926 9550 14978 9602
rect 7038 9382 7090 9434
rect 7142 9382 7194 9434
rect 7246 9382 7298 9434
rect 12862 9382 12914 9434
rect 12966 9382 13018 9434
rect 13070 9382 13122 9434
rect 18686 9382 18738 9434
rect 18790 9382 18842 9434
rect 18894 9382 18946 9434
rect 24510 9382 24562 9434
rect 24614 9382 24666 9434
rect 24718 9382 24770 9434
rect 4510 9214 4562 9266
rect 9662 9214 9714 9266
rect 16270 9214 16322 9266
rect 16606 9214 16658 9266
rect 22094 9214 22146 9266
rect 5406 9102 5458 9154
rect 6862 9102 6914 9154
rect 10670 9102 10722 9154
rect 14926 9102 14978 9154
rect 22878 9102 22930 9154
rect 4846 8990 4898 9042
rect 5630 8990 5682 9042
rect 6078 8990 6130 9042
rect 9998 8990 10050 9042
rect 10446 8990 10498 9042
rect 15710 8990 15762 9042
rect 16046 8990 16098 9042
rect 16494 8990 16546 9042
rect 17390 8990 17442 9042
rect 21086 8990 21138 9042
rect 21310 8990 21362 9042
rect 21422 8990 21474 9042
rect 21646 8990 21698 9042
rect 23326 8990 23378 9042
rect 8990 8878 9042 8930
rect 12798 8878 12850 8930
rect 16382 8878 16434 8930
rect 18174 8878 18226 8930
rect 20302 8878 20354 8930
rect 23662 8878 23714 8930
rect 4126 8598 4178 8650
rect 4230 8598 4282 8650
rect 4334 8598 4386 8650
rect 9950 8598 10002 8650
rect 10054 8598 10106 8650
rect 10158 8598 10210 8650
rect 15774 8598 15826 8650
rect 15878 8598 15930 8650
rect 15982 8598 16034 8650
rect 21598 8598 21650 8650
rect 21702 8598 21754 8650
rect 21806 8598 21858 8650
rect 18174 8430 18226 8482
rect 4622 8318 4674 8370
rect 6078 8318 6130 8370
rect 12014 8318 12066 8370
rect 15374 8318 15426 8370
rect 15486 8318 15538 8370
rect 15822 8318 15874 8370
rect 18510 8318 18562 8370
rect 22094 8318 22146 8370
rect 24110 8318 24162 8370
rect 1822 8206 1874 8258
rect 6862 8206 6914 8258
rect 11566 8206 11618 8258
rect 13918 8206 13970 8258
rect 19742 8206 19794 8258
rect 20078 8206 20130 8258
rect 23438 8206 23490 8258
rect 23886 8206 23938 8258
rect 2494 8094 2546 8146
rect 6638 8094 6690 8146
rect 9438 8094 9490 8146
rect 11454 8094 11506 8146
rect 13470 8094 13522 8146
rect 20526 8094 20578 8146
rect 20750 8094 20802 8146
rect 21422 8094 21474 8146
rect 21534 8094 21586 8146
rect 21646 8094 21698 8146
rect 5742 7982 5794 8034
rect 9998 7982 10050 8034
rect 12350 7982 12402 8034
rect 15934 7982 15986 8034
rect 18286 7982 18338 8034
rect 19518 7982 19570 8034
rect 20414 7982 20466 8034
rect 22878 7982 22930 8034
rect 7038 7814 7090 7866
rect 7142 7814 7194 7866
rect 7246 7814 7298 7866
rect 12862 7814 12914 7866
rect 12966 7814 13018 7866
rect 13070 7814 13122 7866
rect 18686 7814 18738 7866
rect 18790 7814 18842 7866
rect 18894 7814 18946 7866
rect 24510 7814 24562 7866
rect 24614 7814 24666 7866
rect 24718 7814 24770 7866
rect 2494 7646 2546 7698
rect 19742 7646 19794 7698
rect 22878 7646 22930 7698
rect 23886 7646 23938 7698
rect 4398 7534 4450 7586
rect 6526 7534 6578 7586
rect 7198 7534 7250 7586
rect 8318 7534 8370 7586
rect 11118 7534 11170 7586
rect 12574 7534 12626 7586
rect 16046 7534 16098 7586
rect 22318 7534 22370 7586
rect 23550 7534 23602 7586
rect 24222 7534 24274 7586
rect 2270 7422 2322 7474
rect 2718 7422 2770 7474
rect 3054 7422 3106 7474
rect 3278 7422 3330 7474
rect 3614 7422 3666 7474
rect 4174 7422 4226 7474
rect 5854 7422 5906 7474
rect 6302 7422 6354 7474
rect 7534 7422 7586 7474
rect 8206 7422 8258 7474
rect 10334 7422 10386 7474
rect 10894 7422 10946 7474
rect 12014 7422 12066 7474
rect 12798 7422 12850 7474
rect 16830 7422 16882 7474
rect 18286 7422 18338 7474
rect 18958 7422 19010 7474
rect 19182 7422 19234 7474
rect 19518 7422 19570 7474
rect 21310 7422 21362 7474
rect 21422 7422 21474 7474
rect 21646 7422 21698 7474
rect 22654 7422 22706 7474
rect 23326 7422 23378 7474
rect 13918 7310 13970 7362
rect 19630 7310 19682 7362
rect 5518 7198 5570 7250
rect 9998 7198 10050 7250
rect 11678 7198 11730 7250
rect 21758 7198 21810 7250
rect 4126 7030 4178 7082
rect 4230 7030 4282 7082
rect 4334 7030 4386 7082
rect 9950 7030 10002 7082
rect 10054 7030 10106 7082
rect 10158 7030 10210 7082
rect 15774 7030 15826 7082
rect 15878 7030 15930 7082
rect 15982 7030 16034 7082
rect 21598 7030 21650 7082
rect 21702 7030 21754 7082
rect 21806 7030 21858 7082
rect 9102 6862 9154 6914
rect 18510 6750 18562 6802
rect 20638 6750 20690 6802
rect 24222 6750 24274 6802
rect 4510 6638 4562 6690
rect 9662 6638 9714 6690
rect 11790 6638 11842 6690
rect 17726 6638 17778 6690
rect 21310 6638 21362 6690
rect 22094 6638 22146 6690
rect 8094 6526 8146 6578
rect 8766 6526 8818 6578
rect 9774 6526 9826 6578
rect 4174 6414 4226 6466
rect 7758 6414 7810 6466
rect 12014 6414 12066 6466
rect 7038 6246 7090 6298
rect 7142 6246 7194 6298
rect 7246 6246 7298 6298
rect 12862 6246 12914 6298
rect 12966 6246 13018 6298
rect 13070 6246 13122 6298
rect 18686 6246 18738 6298
rect 18790 6246 18842 6298
rect 18894 6246 18946 6298
rect 24510 6246 24562 6298
rect 24614 6246 24666 6298
rect 24718 6246 24770 6298
rect 20638 6078 20690 6130
rect 22878 6078 22930 6130
rect 3614 5966 3666 6018
rect 6862 5966 6914 6018
rect 13470 5966 13522 6018
rect 2942 5854 2994 5906
rect 6190 5854 6242 5906
rect 14254 5854 14306 5906
rect 20974 5854 21026 5906
rect 23102 5854 23154 5906
rect 23550 5854 23602 5906
rect 23998 5854 24050 5906
rect 5742 5742 5794 5794
rect 8990 5742 9042 5794
rect 11342 5742 11394 5794
rect 4126 5462 4178 5514
rect 4230 5462 4282 5514
rect 4334 5462 4386 5514
rect 9950 5462 10002 5514
rect 10054 5462 10106 5514
rect 10158 5462 10210 5514
rect 15774 5462 15826 5514
rect 15878 5462 15930 5514
rect 15982 5462 16034 5514
rect 21598 5462 21650 5514
rect 21702 5462 21754 5514
rect 21806 5462 21858 5514
rect 23102 5182 23154 5234
rect 23550 5182 23602 5234
rect 23774 5070 23826 5122
rect 7038 4678 7090 4730
rect 7142 4678 7194 4730
rect 7246 4678 7298 4730
rect 12862 4678 12914 4730
rect 12966 4678 13018 4730
rect 13070 4678 13122 4730
rect 18686 4678 18738 4730
rect 18790 4678 18842 4730
rect 18894 4678 18946 4730
rect 24510 4678 24562 4730
rect 24614 4678 24666 4730
rect 24718 4678 24770 4730
rect 23886 4510 23938 4562
rect 24222 4286 24274 4338
rect 23662 4174 23714 4226
rect 4126 3894 4178 3946
rect 4230 3894 4282 3946
rect 4334 3894 4386 3946
rect 9950 3894 10002 3946
rect 10054 3894 10106 3946
rect 10158 3894 10210 3946
rect 15774 3894 15826 3946
rect 15878 3894 15930 3946
rect 15982 3894 16034 3946
rect 21598 3894 21650 3946
rect 21702 3894 21754 3946
rect 21806 3894 21858 3946
rect 23438 3390 23490 3442
rect 23662 3390 23714 3442
rect 23998 3390 24050 3442
rect 7038 3110 7090 3162
rect 7142 3110 7194 3162
rect 7246 3110 7298 3162
rect 12862 3110 12914 3162
rect 12966 3110 13018 3162
rect 13070 3110 13122 3162
rect 18686 3110 18738 3162
rect 18790 3110 18842 3162
rect 18894 3110 18946 3162
rect 24510 3110 24562 3162
rect 24614 3110 24666 3162
rect 24718 3110 24770 3162
<< metal2 >>
rect 4256 25200 4368 26000
rect 12768 25200 12880 26000
rect 21280 25200 21392 26000
rect 4284 23548 4340 25200
rect 3948 23492 4340 23548
rect 3500 20132 3556 20142
rect 3500 20018 3556 20076
rect 3500 19966 3502 20018
rect 3554 19966 3556 20018
rect 1820 19236 1876 19246
rect 1820 19142 1876 19180
rect 3500 19236 3556 19966
rect 3948 19460 4004 23492
rect 4124 22764 4388 22774
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4124 22698 4388 22708
rect 9948 22764 10212 22774
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 9948 22698 10212 22708
rect 12684 22484 12740 22494
rect 12796 22484 12852 25200
rect 20300 24052 20356 24062
rect 15772 22764 16036 22774
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 15772 22698 16036 22708
rect 12684 22482 13188 22484
rect 12684 22430 12686 22482
rect 12738 22430 13188 22482
rect 12684 22428 13188 22430
rect 12684 22418 12740 22428
rect 13132 22370 13188 22428
rect 13132 22318 13134 22370
rect 13186 22318 13188 22370
rect 13132 22306 13188 22318
rect 17500 22372 17556 22382
rect 13468 22146 13524 22158
rect 13468 22094 13470 22146
rect 13522 22094 13524 22146
rect 7036 21980 7300 21990
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7036 21914 7300 21924
rect 12860 21980 13124 21990
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 12860 21914 13124 21924
rect 8540 21700 8596 21710
rect 8540 21698 8820 21700
rect 8540 21646 8542 21698
rect 8594 21646 8820 21698
rect 8540 21644 8820 21646
rect 8540 21634 8596 21644
rect 5068 21588 5124 21598
rect 4124 21196 4388 21206
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4124 21130 4388 21140
rect 5068 20132 5124 21532
rect 8316 21586 8372 21598
rect 8316 21534 8318 21586
rect 8370 21534 8372 21586
rect 5740 21476 5796 21486
rect 7868 21476 7924 21486
rect 8316 21476 8372 21534
rect 5740 21474 6244 21476
rect 5740 21422 5742 21474
rect 5794 21422 6244 21474
rect 5740 21420 6244 21422
rect 5740 21410 5796 21420
rect 5068 20066 5124 20076
rect 4172 20020 4228 20030
rect 4172 20018 5012 20020
rect 4172 19966 4174 20018
rect 4226 19966 5012 20018
rect 4172 19964 5012 19966
rect 4172 19954 4228 19964
rect 4124 19628 4388 19638
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4124 19562 4388 19572
rect 3948 19404 4564 19460
rect 3500 19170 3556 19180
rect 2492 19124 2548 19134
rect 2492 19122 2996 19124
rect 2492 19070 2494 19122
rect 2546 19070 2996 19122
rect 2492 19068 2996 19070
rect 2492 19058 2548 19068
rect 2940 17892 2996 19068
rect 3388 18562 3444 18574
rect 3388 18510 3390 18562
rect 3442 18510 3444 18562
rect 2716 17890 2996 17892
rect 2716 17838 2942 17890
rect 2994 17838 2996 17890
rect 2716 17836 2996 17838
rect 2380 17668 2436 17678
rect 2380 17574 2436 17612
rect 2156 17442 2212 17454
rect 2156 17390 2158 17442
rect 2210 17390 2212 17442
rect 2156 16324 2212 17390
rect 2212 16268 2324 16324
rect 2156 16258 2212 16268
rect 2268 15540 2324 16268
rect 2716 15988 2772 17836
rect 2940 17826 2996 17836
rect 3276 18226 3332 18238
rect 3276 18174 3278 18226
rect 3330 18174 3332 18226
rect 2828 17668 2884 17678
rect 2828 17574 2884 17612
rect 3276 17668 3332 18174
rect 3276 17602 3332 17612
rect 3388 17556 3444 18510
rect 3612 18450 3668 18462
rect 3948 18452 4004 18462
rect 3612 18398 3614 18450
rect 3666 18398 3668 18450
rect 3612 18340 3668 18398
rect 3612 18274 3668 18284
rect 3724 18396 3948 18452
rect 3612 17892 3668 17902
rect 3724 17892 3780 18396
rect 3948 18358 4004 18396
rect 4396 18452 4452 18462
rect 4396 18358 4452 18396
rect 3612 17890 3780 17892
rect 3612 17838 3614 17890
rect 3666 17838 3780 17890
rect 3612 17836 3780 17838
rect 3836 18228 3892 18238
rect 4060 18228 4116 18238
rect 3612 17826 3668 17836
rect 3836 17778 3892 18172
rect 3836 17726 3838 17778
rect 3890 17726 3892 17778
rect 3836 17714 3892 17726
rect 3948 18226 4116 18228
rect 3948 18174 4062 18226
rect 4114 18174 4116 18226
rect 3948 18172 4116 18174
rect 3388 17490 3444 17500
rect 3276 17442 3332 17454
rect 3276 17390 3278 17442
rect 3330 17390 3332 17442
rect 2828 16324 2884 16334
rect 2828 16230 2884 16268
rect 2044 15426 2100 15438
rect 2044 15374 2046 15426
rect 2098 15374 2100 15426
rect 2044 15316 2100 15374
rect 2268 15426 2324 15484
rect 2268 15374 2270 15426
rect 2322 15374 2324 15426
rect 2268 15362 2324 15374
rect 2492 15874 2548 15886
rect 2492 15822 2494 15874
rect 2546 15822 2548 15874
rect 2044 15250 2100 15260
rect 2156 15202 2212 15214
rect 2156 15150 2158 15202
rect 2210 15150 2212 15202
rect 2156 14756 2212 15150
rect 2492 14868 2548 15822
rect 2604 15316 2660 15326
rect 2604 15222 2660 15260
rect 2716 15204 2772 15932
rect 3164 16100 3220 16110
rect 3164 15986 3220 16044
rect 3164 15934 3166 15986
rect 3218 15934 3220 15986
rect 3164 15922 3220 15934
rect 3276 15988 3332 17390
rect 3948 16324 4004 18172
rect 4060 18162 4116 18172
rect 4124 18060 4388 18070
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4124 17994 4388 18004
rect 4124 16492 4388 16502
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4124 16426 4388 16436
rect 3948 16268 4452 16324
rect 3612 15988 3668 15998
rect 3276 15986 3892 15988
rect 3276 15934 3614 15986
rect 3666 15934 3892 15986
rect 3276 15932 3892 15934
rect 3612 15922 3668 15932
rect 3388 15764 3444 15774
rect 2940 15540 2996 15550
rect 2940 15538 3332 15540
rect 2940 15486 2942 15538
rect 2994 15486 3332 15538
rect 2940 15484 3332 15486
rect 2940 15474 2996 15484
rect 2828 15428 2884 15438
rect 2828 15334 2884 15372
rect 2716 15148 3108 15204
rect 3052 15090 3108 15148
rect 3052 15038 3054 15090
rect 3106 15038 3108 15090
rect 3052 15026 3108 15038
rect 2492 14812 3220 14868
rect 2268 14756 2324 14766
rect 2156 14754 2324 14756
rect 2156 14702 2270 14754
rect 2322 14702 2324 14754
rect 2156 14700 2324 14702
rect 2268 14690 2324 14700
rect 2380 14700 2884 14756
rect 2380 13860 2436 14700
rect 2828 14642 2884 14700
rect 2828 14590 2830 14642
rect 2882 14590 2884 14642
rect 2828 14578 2884 14590
rect 2604 14532 2660 14542
rect 2604 14438 2660 14476
rect 2716 14420 2772 14430
rect 2716 14326 2772 14364
rect 2940 14308 2996 14318
rect 3164 14308 3220 14812
rect 3276 14756 3332 15484
rect 3388 15314 3444 15708
rect 3388 15262 3390 15314
rect 3442 15262 3444 15314
rect 3388 15250 3444 15262
rect 3500 15428 3556 15438
rect 3276 14700 3444 14756
rect 3276 14532 3332 14542
rect 3276 14438 3332 14476
rect 3388 14308 3444 14700
rect 3500 14418 3556 15372
rect 3836 15426 3892 15932
rect 3836 15374 3838 15426
rect 3890 15374 3892 15426
rect 3836 15362 3892 15374
rect 3948 15204 4004 16268
rect 4060 15988 4116 15998
rect 4060 15894 4116 15932
rect 4284 15988 4340 15998
rect 4284 15894 4340 15932
rect 4396 15986 4452 16268
rect 4396 15934 4398 15986
rect 4450 15934 4452 15986
rect 4396 15922 4452 15934
rect 3836 15148 4004 15204
rect 4172 15874 4228 15886
rect 4172 15822 4174 15874
rect 4226 15822 4228 15874
rect 3836 15092 3892 15148
rect 4172 15092 4228 15822
rect 4396 15764 4452 15774
rect 4396 15314 4452 15708
rect 4396 15262 4398 15314
rect 4450 15262 4452 15314
rect 4396 15250 4452 15262
rect 3612 15036 3892 15092
rect 3948 15036 4228 15092
rect 3612 14530 3668 15036
rect 3612 14478 3614 14530
rect 3666 14478 3668 14530
rect 3612 14466 3668 14478
rect 3948 14532 4004 15036
rect 4124 14924 4388 14934
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4124 14858 4388 14868
rect 4172 14532 4228 14542
rect 3948 14530 4228 14532
rect 3948 14478 4174 14530
rect 4226 14478 4228 14530
rect 3948 14476 4228 14478
rect 4172 14466 4228 14476
rect 3500 14366 3502 14418
rect 3554 14366 3556 14418
rect 3500 14354 3556 14366
rect 2940 14306 3220 14308
rect 2940 14254 2942 14306
rect 2994 14254 3220 14306
rect 2940 14252 3220 14254
rect 3276 14252 3444 14308
rect 4396 14306 4452 14318
rect 4396 14254 4398 14306
rect 4450 14254 4452 14306
rect 2940 14242 2996 14252
rect 3276 14196 3332 14252
rect 3052 14140 3332 14196
rect 2492 13860 2548 13870
rect 2380 13858 2548 13860
rect 2380 13806 2494 13858
rect 2546 13806 2548 13858
rect 2380 13804 2548 13806
rect 2492 13794 2548 13804
rect 1820 13746 1876 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 12180 1876 13694
rect 3052 13186 3108 14140
rect 4396 13636 4452 14254
rect 4508 14308 4564 19404
rect 4956 19458 5012 19964
rect 4956 19406 4958 19458
rect 5010 19406 5012 19458
rect 4620 19348 4676 19358
rect 4620 19254 4676 19292
rect 4844 18450 4900 18462
rect 4844 18398 4846 18450
rect 4898 18398 4900 18450
rect 4844 18340 4900 18398
rect 4844 18274 4900 18284
rect 4620 17892 4676 17902
rect 4620 17798 4676 17836
rect 4732 17668 4788 17678
rect 4732 17574 4788 17612
rect 4620 17556 4676 17566
rect 4620 17462 4676 17500
rect 4844 16100 4900 16110
rect 4620 15876 4676 15886
rect 4620 15428 4676 15820
rect 4844 15764 4900 16044
rect 4844 15698 4900 15708
rect 4956 15988 5012 19406
rect 5068 19122 5124 19134
rect 5068 19070 5070 19122
rect 5122 19070 5124 19122
rect 5068 17892 5124 19070
rect 6188 18788 6244 21420
rect 7868 21474 8372 21476
rect 7868 21422 7870 21474
rect 7922 21422 8372 21474
rect 7868 21420 8372 21422
rect 7868 21410 7924 21420
rect 8316 21252 8372 21420
rect 8316 21196 8596 21252
rect 7980 20804 8036 20814
rect 7980 20710 8036 20748
rect 8428 20804 8484 20842
rect 8428 20738 8484 20748
rect 7868 20690 7924 20702
rect 7868 20638 7870 20690
rect 7922 20638 7924 20690
rect 7036 20412 7300 20422
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7036 20346 7300 20356
rect 6972 20244 7028 20254
rect 6972 20130 7028 20188
rect 6972 20078 6974 20130
rect 7026 20078 7028 20130
rect 6972 20066 7028 20078
rect 6300 19908 6356 19918
rect 6860 19908 6916 19918
rect 6300 19906 6916 19908
rect 6300 19854 6302 19906
rect 6354 19854 6862 19906
rect 6914 19854 6916 19906
rect 6300 19852 6916 19854
rect 6300 19842 6356 19852
rect 6748 19348 6804 19358
rect 6188 18732 6468 18788
rect 5628 18564 5684 18574
rect 6188 18564 6244 18574
rect 5628 18562 6244 18564
rect 5628 18510 5630 18562
rect 5682 18510 6190 18562
rect 6242 18510 6244 18562
rect 5628 18508 6244 18510
rect 5516 18450 5572 18462
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 5516 18340 5572 18398
rect 5516 18274 5572 18284
rect 5068 17826 5124 17836
rect 5628 17668 5684 18508
rect 6188 18498 6244 18508
rect 6300 18452 6356 18462
rect 5628 17602 5684 17612
rect 5740 17892 5796 17902
rect 5740 17666 5796 17836
rect 6300 17778 6356 18396
rect 6300 17726 6302 17778
rect 6354 17726 6356 17778
rect 6300 17714 6356 17726
rect 5740 17614 5742 17666
rect 5794 17614 5796 17666
rect 5740 17602 5796 17614
rect 5964 17444 6020 17454
rect 5516 17442 6020 17444
rect 5516 17390 5966 17442
rect 6018 17390 6020 17442
rect 5516 17388 6020 17390
rect 5180 17108 5236 17118
rect 5180 16994 5236 17052
rect 5180 16942 5182 16994
rect 5234 16942 5236 16994
rect 5180 16930 5236 16942
rect 5292 16660 5348 16670
rect 5292 16566 5348 16604
rect 4956 15540 5012 15932
rect 4620 14530 4676 15372
rect 4732 15484 5012 15540
rect 5292 15876 5348 15886
rect 4732 15314 4788 15484
rect 5292 15426 5348 15820
rect 5516 15764 5572 17388
rect 5964 17378 6020 17388
rect 5964 17108 6020 17118
rect 5964 17014 6020 17052
rect 6300 17108 6356 17118
rect 6412 17108 6468 18732
rect 6524 18228 6580 18238
rect 6524 18134 6580 18172
rect 6748 17666 6804 19292
rect 6860 19236 6916 19852
rect 7308 19908 7364 19918
rect 7868 19908 7924 20638
rect 8540 20690 8596 21196
rect 8540 20638 8542 20690
rect 8594 20638 8596 20690
rect 8540 20626 8596 20638
rect 7980 20244 8036 20254
rect 7980 20018 8036 20188
rect 8764 20242 8820 21644
rect 9100 21588 9156 21598
rect 8988 21532 9100 21588
rect 8764 20190 8766 20242
rect 8818 20190 8820 20242
rect 7980 19966 7982 20018
rect 8034 19966 8036 20018
rect 7980 19954 8036 19966
rect 8092 20132 8148 20142
rect 7308 19906 7476 19908
rect 7308 19854 7310 19906
rect 7362 19854 7476 19906
rect 7308 19852 7476 19854
rect 7308 19842 7364 19852
rect 6860 18676 6916 19180
rect 7036 18844 7300 18854
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7036 18778 7300 18788
rect 6860 18620 7140 18676
rect 7084 18562 7140 18620
rect 7084 18510 7086 18562
rect 7138 18510 7140 18562
rect 7084 18498 7140 18510
rect 7308 18452 7364 18490
rect 7196 18396 7308 18452
rect 7196 17778 7252 18396
rect 7308 18386 7364 18396
rect 7308 18228 7364 18238
rect 7420 18228 7476 19852
rect 7868 19842 7924 19852
rect 7980 19236 8036 19246
rect 8092 19236 8148 20076
rect 8764 20132 8820 20190
rect 8876 20802 8932 20814
rect 8876 20750 8878 20802
rect 8930 20750 8932 20802
rect 8876 20244 8932 20750
rect 8876 20178 8932 20188
rect 8764 20066 8820 20076
rect 8652 20020 8708 20030
rect 8652 19926 8708 19964
rect 8204 19908 8260 19918
rect 8204 19906 8596 19908
rect 8204 19854 8206 19906
rect 8258 19854 8596 19906
rect 8204 19852 8596 19854
rect 8204 19842 8260 19852
rect 8540 19796 8596 19852
rect 8764 19796 8820 19806
rect 8540 19740 8764 19796
rect 8764 19702 8820 19740
rect 8316 19684 8372 19694
rect 8316 19348 8372 19628
rect 8204 19236 8260 19246
rect 8092 19234 8260 19236
rect 8092 19182 8206 19234
rect 8258 19182 8260 19234
rect 8092 19180 8260 19182
rect 7980 19142 8036 19180
rect 8204 19170 8260 19180
rect 8316 19234 8372 19292
rect 8316 19182 8318 19234
rect 8370 19182 8372 19234
rect 8316 19170 8372 19182
rect 8428 19124 8484 19134
rect 7364 18172 7476 18228
rect 7756 19010 7812 19022
rect 7756 18958 7758 19010
rect 7810 18958 7812 19010
rect 7756 18452 7812 18958
rect 8204 18788 8260 18798
rect 8204 18674 8260 18732
rect 8204 18622 8206 18674
rect 8258 18622 8260 18674
rect 8204 18610 8260 18622
rect 8428 18674 8484 19068
rect 8428 18622 8430 18674
rect 8482 18622 8484 18674
rect 8428 18610 8484 18622
rect 8764 19010 8820 19022
rect 8988 19012 9044 21532
rect 9100 21522 9156 21532
rect 9884 21588 9940 21598
rect 9884 21494 9940 21532
rect 13244 21588 13300 21598
rect 13244 21494 13300 21532
rect 10668 21476 10724 21486
rect 12796 21476 12852 21486
rect 10668 21474 10948 21476
rect 10668 21422 10670 21474
rect 10722 21422 10948 21474
rect 10668 21420 10948 21422
rect 10668 21410 10724 21420
rect 9948 21196 10212 21206
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 9948 21130 10212 21140
rect 9100 21028 9156 21038
rect 10220 21028 10276 21038
rect 9100 21026 9268 21028
rect 9100 20974 9102 21026
rect 9154 20974 9268 21026
rect 9100 20972 9268 20974
rect 9100 20962 9156 20972
rect 9100 19124 9156 19134
rect 9100 19030 9156 19068
rect 9212 19122 9268 20972
rect 9996 21026 10276 21028
rect 9996 20974 10222 21026
rect 10274 20974 10276 21026
rect 9996 20972 10276 20974
rect 9548 20802 9604 20814
rect 9548 20750 9550 20802
rect 9602 20750 9604 20802
rect 9548 20356 9604 20750
rect 9212 19070 9214 19122
rect 9266 19070 9268 19122
rect 8764 18958 8766 19010
rect 8818 18958 8820 19010
rect 8092 18564 8148 18574
rect 8092 18470 8148 18508
rect 8652 18562 8708 18574
rect 8652 18510 8654 18562
rect 8706 18510 8708 18562
rect 7308 18162 7364 18172
rect 7196 17726 7198 17778
rect 7250 17726 7252 17778
rect 7196 17714 7252 17726
rect 6748 17614 6750 17666
rect 6802 17614 6804 17666
rect 6748 17602 6804 17614
rect 7036 17276 7300 17286
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7036 17210 7300 17220
rect 6300 17106 6580 17108
rect 6300 17054 6302 17106
rect 6354 17054 6580 17106
rect 6300 17052 6580 17054
rect 6300 17042 6356 17052
rect 5628 16994 5684 17006
rect 5628 16942 5630 16994
rect 5682 16942 5684 16994
rect 5628 16100 5684 16942
rect 5628 16034 5684 16044
rect 5852 16098 5908 16110
rect 5852 16046 5854 16098
rect 5906 16046 5908 16098
rect 5516 15698 5572 15708
rect 5292 15374 5294 15426
rect 5346 15374 5348 15426
rect 5292 15362 5348 15374
rect 5852 15540 5908 16046
rect 6076 16100 6132 16110
rect 6524 16100 6580 17052
rect 7308 16994 7364 17006
rect 7308 16942 7310 16994
rect 7362 16942 7364 16994
rect 6076 16006 6132 16044
rect 6188 16044 6580 16100
rect 6636 16882 6692 16894
rect 6636 16830 6638 16882
rect 6690 16830 6692 16882
rect 6636 16660 6692 16830
rect 6076 15764 6132 15774
rect 5852 15426 5908 15484
rect 5852 15374 5854 15426
rect 5906 15374 5908 15426
rect 5852 15362 5908 15374
rect 5964 15538 6020 15550
rect 5964 15486 5966 15538
rect 6018 15486 6020 15538
rect 4732 15262 4734 15314
rect 4786 15262 4788 15314
rect 4732 15250 4788 15262
rect 4620 14478 4622 14530
rect 4674 14478 4676 14530
rect 4620 14466 4676 14478
rect 4844 15202 4900 15214
rect 4844 15150 4846 15202
rect 4898 15150 4900 15202
rect 4844 14532 4900 15150
rect 4844 14530 5012 14532
rect 4844 14478 4846 14530
rect 4898 14478 5012 14530
rect 4844 14476 5012 14478
rect 4844 14466 4900 14476
rect 4508 14242 4564 14252
rect 4956 13858 5012 14476
rect 4956 13806 4958 13858
rect 5010 13806 5012 13858
rect 4956 13794 5012 13806
rect 5068 14196 5124 14206
rect 4396 13570 4452 13580
rect 4620 13634 4676 13646
rect 5068 13636 5124 14140
rect 5964 14196 6020 15486
rect 5964 14130 6020 14140
rect 5964 13972 6020 13982
rect 5180 13970 6020 13972
rect 5180 13918 5966 13970
rect 6018 13918 6020 13970
rect 5180 13916 6020 13918
rect 5180 13746 5236 13916
rect 5964 13906 6020 13916
rect 5180 13694 5182 13746
rect 5234 13694 5236 13746
rect 5180 13682 5236 13694
rect 6076 13746 6132 15708
rect 6076 13694 6078 13746
rect 6130 13694 6132 13746
rect 6076 13682 6132 13694
rect 6188 15428 6244 16044
rect 6300 15874 6356 15886
rect 6300 15822 6302 15874
rect 6354 15822 6356 15874
rect 6300 15764 6356 15822
rect 6300 15698 6356 15708
rect 6412 15874 6468 15886
rect 6412 15822 6414 15874
rect 6466 15822 6468 15874
rect 6412 15540 6468 15822
rect 4620 13582 4622 13634
rect 4674 13582 4676 13634
rect 4620 13524 4676 13582
rect 4620 13458 4676 13468
rect 4956 13580 5124 13636
rect 4124 13356 4388 13366
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4124 13290 4388 13300
rect 3052 13134 3054 13186
rect 3106 13134 3108 13186
rect 3052 13122 3108 13134
rect 3388 12962 3444 12974
rect 3388 12910 3390 12962
rect 3442 12910 3444 12962
rect 3164 12738 3220 12750
rect 3164 12686 3166 12738
rect 3218 12686 3220 12738
rect 3164 12404 3220 12686
rect 2716 12348 3220 12404
rect 2716 12290 2772 12348
rect 2716 12238 2718 12290
rect 2770 12238 2772 12290
rect 2716 12226 2772 12238
rect 1932 12180 1988 12190
rect 1820 12178 1988 12180
rect 1820 12126 1934 12178
rect 1986 12126 1988 12178
rect 1820 12124 1988 12126
rect 1820 10612 1876 12124
rect 1932 12114 1988 12124
rect 3388 11620 3444 12910
rect 4956 12962 5012 13580
rect 5404 13524 5460 13534
rect 5404 13300 5460 13468
rect 5516 13524 5572 13534
rect 5964 13524 6020 13534
rect 6188 13524 6244 15372
rect 6300 15484 6468 15540
rect 6300 14642 6356 15484
rect 6412 15316 6468 15354
rect 6412 15250 6468 15260
rect 6636 15316 6692 16604
rect 7308 15876 7364 16942
rect 7756 16996 7812 18396
rect 8652 18452 8708 18510
rect 8764 18564 8820 18958
rect 8764 18498 8820 18508
rect 8876 18956 9044 19012
rect 7756 16930 7812 16940
rect 8204 18228 8260 18238
rect 7644 16884 7700 16894
rect 7644 16790 7700 16828
rect 8092 16884 8148 16894
rect 8092 16790 8148 16828
rect 7980 16660 8036 16670
rect 7868 16658 8036 16660
rect 7868 16606 7982 16658
rect 8034 16606 8036 16658
rect 7868 16604 8036 16606
rect 7420 16100 7476 16110
rect 7420 16006 7476 16044
rect 7308 15810 7364 15820
rect 6636 15250 6692 15260
rect 6748 15764 6804 15774
rect 6748 15428 6804 15708
rect 7036 15708 7300 15718
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7036 15642 7300 15652
rect 6748 15314 6804 15372
rect 7420 15428 7476 15438
rect 7868 15428 7924 16604
rect 7980 16594 8036 16604
rect 8204 16436 8260 18172
rect 8652 18116 8708 18396
rect 8652 18050 8708 18060
rect 8876 17780 8932 18956
rect 9212 18900 9268 19070
rect 8988 18844 9268 18900
rect 9324 20300 9604 20356
rect 8988 18674 9044 18844
rect 9324 18788 9380 20300
rect 9548 20130 9604 20142
rect 9548 20078 9550 20130
rect 9602 20078 9604 20130
rect 9548 19796 9604 20078
rect 9996 20130 10052 20972
rect 10220 20962 10276 20972
rect 10108 20804 10164 20814
rect 10668 20804 10724 20814
rect 10108 20710 10164 20748
rect 10220 20802 10724 20804
rect 10220 20750 10670 20802
rect 10722 20750 10724 20802
rect 10220 20748 10724 20750
rect 10220 20690 10276 20748
rect 10668 20738 10724 20748
rect 10220 20638 10222 20690
rect 10274 20638 10276 20690
rect 10220 20626 10276 20638
rect 10780 20690 10836 20702
rect 10780 20638 10782 20690
rect 10834 20638 10836 20690
rect 9996 20078 9998 20130
rect 10050 20078 10052 20130
rect 9996 20066 10052 20078
rect 10332 20132 10388 20142
rect 9548 19730 9604 19740
rect 9772 20018 9828 20030
rect 9772 19966 9774 20018
rect 9826 19966 9828 20018
rect 9772 19124 9828 19966
rect 9884 19796 9940 19834
rect 9884 19730 9940 19740
rect 9948 19628 10212 19638
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 9948 19562 10212 19572
rect 10332 19346 10388 20076
rect 10780 20132 10836 20638
rect 10780 20066 10836 20076
rect 10892 19460 10948 21420
rect 12684 21474 12852 21476
rect 12684 21422 12798 21474
rect 12850 21422 12852 21474
rect 12684 21420 12852 21422
rect 10892 19394 10948 19404
rect 11228 19796 11284 19806
rect 10332 19294 10334 19346
rect 10386 19294 10388 19346
rect 10332 19282 10388 19294
rect 10556 19234 10612 19246
rect 10556 19182 10558 19234
rect 10610 19182 10612 19234
rect 9772 19068 9940 19124
rect 9324 18722 9380 18732
rect 9436 19010 9492 19022
rect 9436 18958 9438 19010
rect 9490 18958 9492 19010
rect 8988 18622 8990 18674
rect 9042 18622 9044 18674
rect 8988 18610 9044 18622
rect 9436 18676 9492 18958
rect 9436 18620 9828 18676
rect 9772 18450 9828 18620
rect 9772 18398 9774 18450
rect 9826 18398 9828 18450
rect 9772 18386 9828 18398
rect 9884 18452 9940 19068
rect 10108 19012 10164 19022
rect 10108 19010 10276 19012
rect 10108 18958 10110 19010
rect 10162 18958 10276 19010
rect 10108 18956 10276 18958
rect 10108 18946 10164 18956
rect 9884 18386 9940 18396
rect 9548 18338 9604 18350
rect 9548 18286 9550 18338
rect 9602 18286 9604 18338
rect 9548 18228 9604 18286
rect 10108 18228 10164 18238
rect 8876 17686 8932 17724
rect 9212 17780 9268 17790
rect 8540 16996 8596 17006
rect 8540 16902 8596 16940
rect 7420 15426 7924 15428
rect 7420 15374 7422 15426
rect 7474 15374 7924 15426
rect 7420 15372 7924 15374
rect 7420 15362 7476 15372
rect 6748 15262 6750 15314
rect 6802 15262 6804 15314
rect 6748 15250 6804 15262
rect 7868 15314 7924 15372
rect 7868 15262 7870 15314
rect 7922 15262 7924 15314
rect 7868 15250 7924 15262
rect 7980 16380 8260 16436
rect 6300 14590 6302 14642
rect 6354 14590 6356 14642
rect 6300 14578 6356 14590
rect 6524 14980 6580 14990
rect 6524 14530 6580 14924
rect 7868 14644 7924 14654
rect 7980 14644 8036 16380
rect 9212 16100 9268 17724
rect 9548 16996 9604 18172
rect 9548 16930 9604 16940
rect 9772 18226 10164 18228
rect 9772 18174 10110 18226
rect 10162 18174 10164 18226
rect 9772 18172 10164 18174
rect 9436 16884 9492 16894
rect 9436 16790 9492 16828
rect 9772 16772 9828 18172
rect 10108 18162 10164 18172
rect 10220 18228 10276 18956
rect 10444 18564 10500 18574
rect 10556 18564 10612 19182
rect 11228 19234 11284 19740
rect 12012 19460 12068 19470
rect 12684 19460 12740 21420
rect 12796 21410 12852 21420
rect 12860 20412 13124 20422
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 12860 20346 13124 20356
rect 13468 20244 13524 22094
rect 15596 21588 15652 21598
rect 13916 21476 13972 21486
rect 15148 21476 15204 21486
rect 13916 21474 14084 21476
rect 13916 21422 13918 21474
rect 13970 21422 14084 21474
rect 13916 21420 14084 21422
rect 13916 21410 13972 21420
rect 13356 20188 13524 20244
rect 14028 20242 14084 21420
rect 14028 20190 14030 20242
rect 14082 20190 14084 20242
rect 12796 19460 12852 19470
rect 12684 19404 12796 19460
rect 12012 19366 12068 19404
rect 12796 19394 12852 19404
rect 11228 19182 11230 19234
rect 11282 19182 11284 19234
rect 11228 19170 11284 19182
rect 12012 19234 12068 19246
rect 12012 19182 12014 19234
rect 12066 19182 12068 19234
rect 11900 19124 11956 19134
rect 11900 19030 11956 19068
rect 10892 19010 10948 19022
rect 11340 19012 11396 19022
rect 11564 19012 11620 19022
rect 10892 18958 10894 19010
rect 10946 18958 10948 19010
rect 10892 18676 10948 18958
rect 11116 18956 11340 19012
rect 10892 18610 10948 18620
rect 11004 18788 11060 18798
rect 10780 18564 10836 18574
rect 10556 18508 10780 18564
rect 10444 18470 10500 18508
rect 10780 18450 10836 18508
rect 10780 18398 10782 18450
rect 10834 18398 10836 18450
rect 10780 18386 10836 18398
rect 11004 18450 11060 18732
rect 11116 18564 11172 18956
rect 11340 18918 11396 18956
rect 11452 19010 11620 19012
rect 11452 18958 11566 19010
rect 11618 18958 11620 19010
rect 11452 18956 11620 18958
rect 11452 18676 11508 18956
rect 11564 18946 11620 18956
rect 12012 19012 12068 19182
rect 12460 19234 12516 19246
rect 12460 19182 12462 19234
rect 12514 19182 12516 19234
rect 12012 18946 12068 18956
rect 12348 19124 12404 19134
rect 11340 18620 11508 18676
rect 11564 18676 11620 18686
rect 11228 18564 11284 18574
rect 11116 18508 11228 18564
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 10220 18162 10276 18172
rect 10556 18338 10612 18350
rect 10556 18286 10558 18338
rect 10610 18286 10612 18338
rect 9948 18060 10212 18070
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 9948 17994 10212 18004
rect 10556 17444 10612 18286
rect 10108 17388 10612 17444
rect 10892 17780 10948 17790
rect 10108 16882 10164 17388
rect 10108 16830 10110 16882
rect 10162 16830 10164 16882
rect 10108 16818 10164 16830
rect 10332 16996 10388 17006
rect 10332 16882 10388 16940
rect 10332 16830 10334 16882
rect 10386 16830 10388 16882
rect 10332 16818 10388 16830
rect 10892 16882 10948 17724
rect 10892 16830 10894 16882
rect 10946 16830 10948 16882
rect 10892 16818 10948 16830
rect 9884 16772 9940 16782
rect 9772 16770 9940 16772
rect 9772 16718 9886 16770
rect 9938 16718 9940 16770
rect 9772 16716 9940 16718
rect 9884 16706 9940 16716
rect 9948 16492 10212 16502
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 9948 16426 10212 16436
rect 10220 16212 10276 16222
rect 11004 16212 11060 18398
rect 10220 16210 11060 16212
rect 10220 16158 10222 16210
rect 10274 16158 11060 16210
rect 10220 16156 11060 16158
rect 10220 16146 10276 16156
rect 8092 15986 8148 15998
rect 8092 15934 8094 15986
rect 8146 15934 8148 15986
rect 8092 15540 8148 15934
rect 8540 15540 8596 15550
rect 8092 15538 8596 15540
rect 8092 15486 8094 15538
rect 8146 15486 8542 15538
rect 8594 15486 8596 15538
rect 8092 15484 8596 15486
rect 8092 14980 8148 15484
rect 8540 15474 8596 15484
rect 8652 15428 8708 15438
rect 8652 15334 8708 15372
rect 8092 14914 8148 14924
rect 8540 15090 8596 15102
rect 8540 15038 8542 15090
rect 8594 15038 8596 15090
rect 7868 14642 8036 14644
rect 7868 14590 7870 14642
rect 7922 14590 8036 14642
rect 7868 14588 8036 14590
rect 7868 14578 7924 14588
rect 6524 14478 6526 14530
rect 6578 14478 6580 14530
rect 6300 13748 6356 13758
rect 6524 13748 6580 14478
rect 8092 14532 8148 14542
rect 8540 14532 8596 15038
rect 8092 14530 8596 14532
rect 8092 14478 8094 14530
rect 8146 14478 8596 14530
rect 8092 14476 8596 14478
rect 9212 14530 9268 16044
rect 11228 15986 11284 18508
rect 11340 18562 11396 18620
rect 11564 18582 11620 18620
rect 11340 18510 11342 18562
rect 11394 18510 11396 18562
rect 11340 18498 11396 18510
rect 11788 18562 11844 18574
rect 11788 18510 11790 18562
rect 11842 18510 11844 18562
rect 11788 18452 11844 18510
rect 12236 18452 12292 18462
rect 11788 18396 12236 18452
rect 12236 18358 12292 18396
rect 11452 18226 11508 18238
rect 11452 18174 11454 18226
rect 11506 18174 11508 18226
rect 11452 17108 11508 18174
rect 11452 17042 11508 17052
rect 12124 18226 12180 18238
rect 12124 18174 12126 18226
rect 12178 18174 12180 18226
rect 12124 16996 12180 18174
rect 12012 16940 12124 16996
rect 11564 16884 11620 16894
rect 11564 16324 11620 16828
rect 11676 16772 11732 16782
rect 11676 16770 11956 16772
rect 11676 16718 11678 16770
rect 11730 16718 11956 16770
rect 11676 16716 11956 16718
rect 11676 16706 11732 16716
rect 11564 16098 11620 16268
rect 11564 16046 11566 16098
rect 11618 16046 11620 16098
rect 11564 16034 11620 16046
rect 11900 16098 11956 16716
rect 11900 16046 11902 16098
rect 11954 16046 11956 16098
rect 11900 16034 11956 16046
rect 11228 15934 11230 15986
rect 11282 15934 11284 15986
rect 11228 15922 11284 15934
rect 12012 15092 12068 16940
rect 12124 16930 12180 16940
rect 12348 16772 12404 19068
rect 12460 18676 12516 19182
rect 12684 19236 12740 19246
rect 12684 19142 12740 19180
rect 12860 18844 13124 18854
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 12860 18778 13124 18788
rect 12460 18610 12516 18620
rect 13356 18674 13412 20188
rect 14028 20178 14084 20190
rect 14252 20188 14532 20244
rect 14252 20130 14308 20188
rect 14252 20078 14254 20130
rect 14306 20078 14308 20130
rect 14252 20066 14308 20078
rect 14476 20132 14532 20188
rect 14924 20132 14980 20142
rect 14476 20130 14980 20132
rect 14476 20078 14926 20130
rect 14978 20078 14980 20130
rect 14476 20076 14980 20078
rect 13916 20020 13972 20030
rect 13916 20018 14196 20020
rect 13916 19966 13918 20018
rect 13970 19966 14196 20018
rect 13916 19964 14196 19966
rect 13916 19954 13972 19964
rect 14140 19236 14196 19964
rect 14364 20018 14420 20030
rect 14364 19966 14366 20018
rect 14418 19966 14420 20018
rect 14364 19346 14420 19966
rect 14364 19294 14366 19346
rect 14418 19294 14420 19346
rect 14364 19282 14420 19294
rect 14252 19236 14308 19246
rect 14140 19234 14308 19236
rect 14140 19182 14254 19234
rect 14306 19182 14308 19234
rect 14140 19180 14308 19182
rect 13804 19124 13860 19134
rect 13804 19030 13860 19068
rect 13916 19012 13972 19022
rect 14252 19012 14308 19180
rect 14476 19124 14532 20076
rect 14924 20066 14980 20076
rect 15148 20018 15204 21420
rect 15596 20804 15652 21532
rect 16044 21476 16100 21486
rect 16044 21382 16100 21420
rect 15772 21196 16036 21206
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 15772 21130 16036 21140
rect 15596 20710 15652 20748
rect 16268 20692 16324 20702
rect 16268 20690 16436 20692
rect 16268 20638 16270 20690
rect 16322 20638 16436 20690
rect 16268 20636 16436 20638
rect 16268 20626 16324 20636
rect 15148 19966 15150 20018
rect 15202 19966 15204 20018
rect 14476 19030 14532 19068
rect 14924 19234 14980 19246
rect 14924 19182 14926 19234
rect 14978 19182 14980 19234
rect 13916 19010 14196 19012
rect 13916 18958 13918 19010
rect 13970 18958 14196 19010
rect 13916 18956 14196 18958
rect 13916 18946 13972 18956
rect 13356 18622 13358 18674
rect 13410 18622 13412 18674
rect 12684 18562 12740 18574
rect 12684 18510 12686 18562
rect 12738 18510 12740 18562
rect 12684 18340 12740 18510
rect 12684 18274 12740 18284
rect 12908 18450 12964 18462
rect 12908 18398 12910 18450
rect 12962 18398 12964 18450
rect 12908 18228 12964 18398
rect 13356 18452 13412 18622
rect 14140 18676 14196 18956
rect 14252 18946 14308 18956
rect 14924 18900 14980 19182
rect 15036 19234 15092 19246
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 15036 19012 15092 19182
rect 15036 18946 15092 18956
rect 14812 18676 14868 18686
rect 14140 18620 14756 18676
rect 13356 18386 13412 18396
rect 13692 18562 13748 18574
rect 13692 18510 13694 18562
rect 13746 18510 13748 18562
rect 12684 17666 12740 17678
rect 12684 17614 12686 17666
rect 12738 17614 12740 17666
rect 12684 16884 12740 17614
rect 12908 17556 12964 18172
rect 13692 18228 13748 18510
rect 14700 18450 14756 18620
rect 14812 18582 14868 18620
rect 14924 18564 14980 18844
rect 14924 18498 14980 18508
rect 14700 18398 14702 18450
rect 14754 18398 14756 18450
rect 14700 18386 14756 18398
rect 14924 18340 14980 18350
rect 14924 18246 14980 18284
rect 13692 18162 13748 18172
rect 14364 18228 14420 18238
rect 14252 17892 14308 17902
rect 14364 17892 14420 18172
rect 14476 18228 14532 18238
rect 14476 18226 14868 18228
rect 14476 18174 14478 18226
rect 14530 18174 14868 18226
rect 14476 18172 14868 18174
rect 14476 18162 14532 18172
rect 14252 17890 14420 17892
rect 14252 17838 14254 17890
rect 14306 17838 14420 17890
rect 14252 17836 14420 17838
rect 14252 17826 14308 17836
rect 14140 17668 14196 17678
rect 14140 17666 14756 17668
rect 14140 17614 14142 17666
rect 14194 17614 14756 17666
rect 14140 17612 14756 17614
rect 14140 17602 14196 17612
rect 12908 17490 12964 17500
rect 14252 17442 14308 17454
rect 14252 17390 14254 17442
rect 14306 17390 14308 17442
rect 12860 17276 13124 17286
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 12860 17210 13124 17220
rect 14140 16996 14196 17006
rect 14252 16996 14308 17390
rect 12684 16818 12740 16828
rect 13804 16994 14308 16996
rect 13804 16942 14142 16994
rect 14194 16942 14308 16994
rect 13804 16940 14308 16942
rect 12124 16716 12404 16772
rect 13804 16770 13860 16940
rect 14140 16930 14196 16940
rect 13804 16718 13806 16770
rect 13858 16718 13860 16770
rect 12124 15986 12180 16716
rect 13804 16706 13860 16718
rect 14252 16660 14308 16670
rect 14252 16658 14644 16660
rect 14252 16606 14254 16658
rect 14306 16606 14644 16658
rect 14252 16604 14644 16606
rect 14252 16594 14308 16604
rect 13804 16548 13860 16558
rect 12684 16324 12740 16334
rect 12684 16210 12740 16268
rect 12684 16158 12686 16210
rect 12738 16158 12740 16210
rect 12684 16146 12740 16158
rect 12124 15934 12126 15986
rect 12178 15934 12180 15986
rect 12124 15922 12180 15934
rect 12236 15988 12292 15998
rect 12236 15894 12292 15932
rect 12860 15708 13124 15718
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 12860 15642 13124 15652
rect 13020 15540 13076 15550
rect 12012 15026 12068 15036
rect 12124 15538 13076 15540
rect 12124 15486 13022 15538
rect 13074 15486 13076 15538
rect 12124 15484 13076 15486
rect 9948 14924 10212 14934
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 9948 14858 10212 14868
rect 12012 14644 12068 14654
rect 9212 14478 9214 14530
rect 9266 14478 9268 14530
rect 7196 14420 7252 14430
rect 8092 14420 8148 14476
rect 7196 14418 7476 14420
rect 7196 14366 7198 14418
rect 7250 14366 7476 14418
rect 7196 14364 7476 14366
rect 7196 14354 7252 14364
rect 7036 14140 7300 14150
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7036 14074 7300 14084
rect 6300 13746 6580 13748
rect 6300 13694 6302 13746
rect 6354 13694 6580 13746
rect 6300 13692 6580 13694
rect 6300 13682 6356 13692
rect 5516 13522 5908 13524
rect 5516 13470 5518 13522
rect 5570 13470 5908 13522
rect 5516 13468 5908 13470
rect 5516 13458 5572 13468
rect 5404 13244 5796 13300
rect 4956 12910 4958 12962
rect 5010 12910 5012 12962
rect 4956 12898 5012 12910
rect 4732 12738 4788 12750
rect 4732 12686 4734 12738
rect 4786 12686 4788 12738
rect 4124 11788 4388 11798
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4124 11722 4388 11732
rect 4732 11732 4788 12686
rect 4732 11666 4788 11676
rect 4844 12066 4900 12078
rect 4844 12014 4846 12066
rect 4898 12014 4900 12066
rect 3388 11554 3444 11564
rect 1820 9826 1876 10556
rect 2268 10892 3220 10948
rect 2268 10610 2324 10892
rect 3164 10834 3220 10892
rect 3164 10782 3166 10834
rect 3218 10782 3220 10834
rect 3164 10770 3220 10782
rect 2268 10558 2270 10610
rect 2322 10558 2324 10610
rect 2268 10546 2324 10558
rect 2492 10722 2548 10734
rect 2492 10670 2494 10722
rect 2546 10670 2548 10722
rect 2492 9938 2548 10670
rect 3500 10724 3556 10734
rect 3500 10610 3556 10668
rect 4284 10724 4340 10734
rect 4620 10724 4676 10734
rect 4284 10722 4564 10724
rect 4284 10670 4286 10722
rect 4338 10670 4564 10722
rect 4284 10668 4564 10670
rect 4284 10658 4340 10668
rect 3500 10558 3502 10610
rect 3554 10558 3556 10610
rect 3500 10546 3556 10558
rect 3948 10610 4004 10622
rect 3948 10558 3950 10610
rect 4002 10558 4004 10610
rect 2492 9886 2494 9938
rect 2546 9886 2548 9938
rect 2492 9874 2548 9886
rect 1820 9774 1822 9826
rect 1874 9774 1876 9826
rect 1820 8428 1876 9774
rect 3612 8484 3668 8494
rect 1820 8372 2996 8428
rect 1820 8258 1876 8372
rect 1820 8206 1822 8258
rect 1874 8206 1876 8258
rect 1820 8194 1876 8206
rect 2492 8146 2548 8158
rect 2492 8094 2494 8146
rect 2546 8094 2548 8146
rect 2492 7698 2548 8094
rect 2492 7646 2494 7698
rect 2546 7646 2548 7698
rect 2492 7634 2548 7646
rect 2268 7476 2324 7486
rect 2716 7476 2772 7486
rect 2268 7474 2772 7476
rect 2268 7422 2270 7474
rect 2322 7422 2718 7474
rect 2770 7422 2772 7474
rect 2268 7420 2772 7422
rect 2268 7410 2324 7420
rect 2716 7410 2772 7420
rect 2940 5906 2996 8372
rect 3052 7476 3108 7486
rect 3276 7476 3332 7486
rect 3052 7474 3332 7476
rect 3052 7422 3054 7474
rect 3106 7422 3278 7474
rect 3330 7422 3332 7474
rect 3052 7420 3332 7422
rect 3052 7410 3108 7420
rect 3276 7410 3332 7420
rect 3612 7474 3668 8428
rect 3948 8428 4004 10558
rect 4124 10220 4388 10230
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4124 10154 4388 10164
rect 4508 9266 4564 10668
rect 4620 9938 4676 10668
rect 4732 10612 4788 10622
rect 4732 10518 4788 10556
rect 4620 9886 4622 9938
rect 4674 9886 4676 9938
rect 4620 9874 4676 9886
rect 4508 9214 4510 9266
rect 4562 9214 4564 9266
rect 4508 9202 4564 9214
rect 4620 9156 4676 9166
rect 4124 8652 4388 8662
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4124 8586 4388 8596
rect 4620 8484 4676 9100
rect 4844 9042 4900 12014
rect 5516 11732 5572 11742
rect 5516 10722 5572 11676
rect 5516 10670 5518 10722
rect 5570 10670 5572 10722
rect 5516 10658 5572 10670
rect 5404 9156 5460 9166
rect 5404 9062 5460 9100
rect 4844 8990 4846 9042
rect 4898 8990 4900 9042
rect 4844 8978 4900 8990
rect 5628 9042 5684 9054
rect 5628 8990 5630 9042
rect 5682 8990 5684 9042
rect 3948 8372 4228 8428
rect 3612 7422 3614 7474
rect 3666 7422 3668 7474
rect 3612 7410 3668 7422
rect 4172 7476 4228 8372
rect 4620 8370 4676 8428
rect 4620 8318 4622 8370
rect 4674 8318 4676 8370
rect 4620 8306 4676 8318
rect 5628 8260 5684 8990
rect 5740 8428 5796 13244
rect 5852 13188 5908 13468
rect 5964 13522 6244 13524
rect 5964 13470 5966 13522
rect 6018 13470 6244 13522
rect 5964 13468 6244 13470
rect 5964 13458 6020 13468
rect 5852 13132 6244 13188
rect 6188 12962 6244 13132
rect 6188 12910 6190 12962
rect 6242 12910 6244 12962
rect 6188 12898 6244 12910
rect 6524 12740 6580 12750
rect 6524 12738 6692 12740
rect 6524 12686 6526 12738
rect 6578 12686 6692 12738
rect 6524 12684 6692 12686
rect 6524 12674 6580 12684
rect 6636 12290 6692 12684
rect 7036 12572 7300 12582
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7036 12506 7300 12516
rect 6636 12238 6638 12290
rect 6690 12238 6692 12290
rect 6636 12226 6692 12238
rect 5852 12178 5908 12190
rect 5852 12126 5854 12178
rect 5906 12126 5908 12178
rect 5852 11508 5908 12126
rect 5852 10612 5908 11452
rect 6748 11508 6804 11518
rect 6748 11414 6804 11452
rect 7036 11004 7300 11014
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7036 10938 7300 10948
rect 5908 10556 6132 10612
rect 5852 10546 5908 10556
rect 6076 9044 6132 10556
rect 7196 9828 7252 9838
rect 7420 9828 7476 14364
rect 8092 14354 8148 14364
rect 8428 14306 8484 14318
rect 8428 14254 8430 14306
rect 8482 14254 8484 14306
rect 8428 13860 8484 14254
rect 8428 13794 8484 13804
rect 9212 13748 9268 14478
rect 11788 14642 12068 14644
rect 11788 14590 12014 14642
rect 12066 14590 12068 14642
rect 11788 14588 12068 14590
rect 9884 14418 9940 14430
rect 9884 14366 9886 14418
rect 9938 14366 9940 14418
rect 9884 13970 9940 14366
rect 9884 13918 9886 13970
rect 9938 13918 9940 13970
rect 9884 13906 9940 13918
rect 9436 13860 9492 13870
rect 9492 13804 9604 13860
rect 9436 13794 9492 13804
rect 9212 13682 9268 13692
rect 9548 13746 9604 13804
rect 9548 13694 9550 13746
rect 9602 13694 9604 13746
rect 9548 13682 9604 13694
rect 11340 13748 11396 13758
rect 11340 13654 11396 13692
rect 8652 13636 8708 13646
rect 8652 13074 8708 13580
rect 9948 13356 10212 13366
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 9948 13290 10212 13300
rect 8652 13022 8654 13074
rect 8706 13022 8708 13074
rect 8652 13010 8708 13022
rect 10780 13076 10836 13086
rect 10780 13074 11508 13076
rect 10780 13022 10782 13074
rect 10834 13022 11508 13074
rect 10780 13020 11508 13022
rect 10780 13010 10836 13020
rect 7868 12962 7924 12974
rect 7868 12910 7870 12962
rect 7922 12910 7924 12962
rect 7868 11508 7924 12910
rect 11340 12852 11396 12862
rect 9772 12290 9828 12302
rect 9772 12238 9774 12290
rect 9826 12238 9828 12290
rect 8764 12068 8820 12078
rect 8764 11974 8820 12012
rect 7868 11442 7924 11452
rect 9100 11956 9156 11966
rect 9100 11508 9156 11900
rect 7196 9826 7476 9828
rect 7196 9774 7198 9826
rect 7250 9774 7476 9826
rect 7196 9772 7476 9774
rect 7644 10498 7700 10510
rect 7644 10446 7646 10498
rect 7698 10446 7700 10498
rect 7196 9762 7252 9772
rect 6860 9602 6916 9614
rect 6860 9550 6862 9602
rect 6914 9550 6916 9602
rect 6860 9154 6916 9550
rect 7036 9436 7300 9446
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7036 9370 7300 9380
rect 6860 9102 6862 9154
rect 6914 9102 6916 9154
rect 6860 9090 6916 9102
rect 6076 9042 6244 9044
rect 6076 8990 6078 9042
rect 6130 8990 6244 9042
rect 6076 8988 6244 8990
rect 6076 8978 6132 8988
rect 5740 8372 6132 8428
rect 6076 8370 6132 8372
rect 6076 8318 6078 8370
rect 6130 8318 6132 8370
rect 6076 8306 6132 8318
rect 5628 8194 5684 8204
rect 5852 8148 5908 8158
rect 4396 8036 4452 8046
rect 4396 7586 4452 7980
rect 5740 8036 5796 8046
rect 5740 7942 5796 7980
rect 4396 7534 4398 7586
rect 4450 7534 4452 7586
rect 4396 7522 4452 7534
rect 5852 7476 5908 8092
rect 4172 7382 4228 7420
rect 5740 7474 5908 7476
rect 5740 7422 5854 7474
rect 5906 7422 5908 7474
rect 5740 7420 5908 7422
rect 4508 7252 4564 7262
rect 4124 7084 4388 7094
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4124 7018 4388 7028
rect 4508 6690 4564 7196
rect 5516 7252 5572 7262
rect 5516 7158 5572 7196
rect 4508 6638 4510 6690
rect 4562 6638 4564 6690
rect 4508 6626 4564 6638
rect 4172 6468 4228 6478
rect 3612 6466 4228 6468
rect 3612 6414 4174 6466
rect 4226 6414 4228 6466
rect 3612 6412 4228 6414
rect 3612 6018 3668 6412
rect 4172 6402 4228 6412
rect 3612 5966 3614 6018
rect 3666 5966 3668 6018
rect 3612 5954 3668 5966
rect 2940 5854 2942 5906
rect 2994 5854 2996 5906
rect 2940 5842 2996 5854
rect 5740 5794 5796 7420
rect 5852 7410 5908 7420
rect 6188 5906 6244 8988
rect 7644 8428 7700 10446
rect 8540 9828 8596 9838
rect 8540 9826 8708 9828
rect 8540 9774 8542 9826
rect 8594 9774 8708 9826
rect 8540 9772 8708 9774
rect 8540 9762 8596 9772
rect 8652 9380 8708 9772
rect 9100 9826 9156 11452
rect 9772 10724 9828 12238
rect 9996 12292 10052 12302
rect 9996 12178 10052 12236
rect 11340 12292 11396 12796
rect 9996 12126 9998 12178
rect 10050 12126 10052 12178
rect 9996 12114 10052 12126
rect 11228 12178 11284 12190
rect 11228 12126 11230 12178
rect 11282 12126 11284 12178
rect 10444 12068 10500 12078
rect 10444 11974 10500 12012
rect 10780 11956 10836 11966
rect 10668 11954 10836 11956
rect 10668 11902 10782 11954
rect 10834 11902 10836 11954
rect 10668 11900 10836 11902
rect 9948 11788 10212 11798
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 9948 11722 10212 11732
rect 9772 10658 9828 10668
rect 9948 10220 10212 10230
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 9948 10154 10212 10164
rect 9100 9774 9102 9826
rect 9154 9774 9156 9826
rect 9100 9762 9156 9774
rect 9884 9714 9940 9726
rect 9884 9662 9886 9714
rect 9938 9662 9940 9714
rect 8764 9604 8820 9614
rect 9884 9604 9940 9662
rect 8764 9602 9940 9604
rect 8764 9550 8766 9602
rect 8818 9550 9940 9602
rect 8764 9548 9940 9550
rect 8764 9538 8820 9548
rect 8652 9324 9716 9380
rect 9660 9266 9716 9324
rect 9660 9214 9662 9266
rect 9714 9214 9716 9266
rect 9660 9202 9716 9214
rect 10668 9154 10724 11900
rect 10780 11890 10836 11900
rect 11228 11956 11284 12126
rect 11228 11890 11284 11900
rect 10668 9102 10670 9154
rect 10722 9102 10724 9154
rect 10668 9090 10724 9102
rect 11004 10722 11060 10734
rect 11004 10670 11006 10722
rect 11058 10670 11060 10722
rect 11004 9940 11060 10670
rect 11340 10722 11396 12236
rect 11340 10670 11342 10722
rect 11394 10670 11396 10722
rect 11340 10658 11396 10670
rect 11452 10612 11508 13020
rect 11564 11396 11620 11406
rect 11564 11302 11620 11340
rect 11564 10612 11620 10622
rect 11452 10610 11620 10612
rect 11452 10558 11566 10610
rect 11618 10558 11620 10610
rect 11452 10556 11620 10558
rect 11564 10546 11620 10556
rect 9996 9044 10052 9054
rect 9996 8950 10052 8988
rect 10444 9042 10500 9054
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 7532 8372 7700 8428
rect 8988 8930 9044 8942
rect 8988 8878 8990 8930
rect 9042 8878 9044 8930
rect 6860 8260 6916 8270
rect 6636 8148 6692 8158
rect 6636 8054 6692 8092
rect 6300 8036 6356 8046
rect 6300 7476 6356 7980
rect 6860 7700 6916 8204
rect 7036 7868 7300 7878
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7036 7802 7300 7812
rect 6860 7634 6916 7644
rect 6524 7588 6580 7598
rect 6524 7494 6580 7532
rect 7196 7588 7252 7598
rect 7196 7494 7252 7532
rect 6300 7382 6356 7420
rect 7532 7474 7588 8372
rect 7532 7422 7534 7474
rect 7586 7422 7588 7474
rect 7532 7410 7588 7422
rect 8204 7700 8260 7710
rect 8204 7474 8260 7644
rect 8316 7588 8372 7598
rect 8316 7494 8372 7532
rect 8204 7422 8206 7474
rect 8258 7422 8260 7474
rect 8204 7410 8260 7422
rect 8988 7476 9044 8878
rect 9948 8652 10212 8662
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 9948 8586 10212 8596
rect 9436 8146 9492 8158
rect 9436 8094 9438 8146
rect 9490 8094 9492 8146
rect 9436 8036 9492 8094
rect 9436 7970 9492 7980
rect 9996 8034 10052 8046
rect 9996 7982 9998 8034
rect 10050 7982 10052 8034
rect 9996 7812 10052 7982
rect 10444 8036 10500 8990
rect 11004 9044 11060 9884
rect 11004 8978 11060 8988
rect 11788 8428 11844 14588
rect 12012 14578 12068 14588
rect 12124 13858 12180 15484
rect 13020 15474 13076 15484
rect 13804 15426 13860 16492
rect 14588 16098 14644 16604
rect 14588 16046 14590 16098
rect 14642 16046 14644 16098
rect 13804 15374 13806 15426
rect 13858 15374 13860 15426
rect 13804 15362 13860 15374
rect 14140 15988 14196 15998
rect 14140 15426 14196 15932
rect 14140 15374 14142 15426
rect 14194 15374 14196 15426
rect 14140 15362 14196 15374
rect 13132 15316 13188 15326
rect 13132 15222 13188 15260
rect 13356 15316 13412 15326
rect 13356 15222 13412 15260
rect 13468 15314 13524 15326
rect 13468 15262 13470 15314
rect 13522 15262 13524 15314
rect 13468 15092 13524 15262
rect 14252 15316 14308 15326
rect 14252 15222 14308 15260
rect 14588 15314 14644 16046
rect 14700 15988 14756 17612
rect 14812 16548 14868 18172
rect 15148 17332 15204 19966
rect 16044 20018 16100 20030
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 16044 19796 16100 19966
rect 16380 19908 16436 20636
rect 17500 20242 17556 22316
rect 18396 22372 18452 22382
rect 17500 20190 17502 20242
rect 17554 20190 17556 20242
rect 17500 20178 17556 20190
rect 17836 21586 17892 21598
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 17836 20804 17892 21534
rect 18396 20914 18452 22316
rect 19628 22372 19684 22382
rect 19964 22372 20020 22382
rect 20300 22372 20356 23996
rect 21308 22596 21364 25200
rect 21596 22764 21860 22774
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21596 22698 21860 22708
rect 21308 22530 21364 22540
rect 22428 22596 22484 22606
rect 22428 22502 22484 22540
rect 19628 22370 20356 22372
rect 19628 22318 19630 22370
rect 19682 22318 19966 22370
rect 20018 22318 20356 22370
rect 19628 22316 20356 22318
rect 20860 22370 20916 22382
rect 20860 22318 20862 22370
rect 20914 22318 20916 22370
rect 19628 22306 19684 22316
rect 19964 22306 20020 22316
rect 20860 22260 20916 22318
rect 21420 22372 21476 22382
rect 21420 22278 21476 22316
rect 21308 22260 21364 22270
rect 20860 22194 20916 22204
rect 21196 22204 21308 22260
rect 20188 22148 20244 22158
rect 20188 22054 20244 22092
rect 21084 22146 21140 22158
rect 21084 22094 21086 22146
rect 21138 22094 21140 22146
rect 18684 21980 18948 21990
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18684 21914 18948 21924
rect 21084 21924 21140 22094
rect 21084 21858 21140 21868
rect 21084 21586 21140 21598
rect 21084 21534 21086 21586
rect 21138 21534 21140 21586
rect 18620 21476 18676 21486
rect 18620 21474 19460 21476
rect 18620 21422 18622 21474
rect 18674 21422 19460 21474
rect 18620 21420 19460 21422
rect 18620 21410 18676 21420
rect 18396 20862 18398 20914
rect 18450 20862 18452 20914
rect 18396 20850 18452 20862
rect 16492 20132 16548 20170
rect 16492 20066 16548 20076
rect 16604 20130 16660 20142
rect 16604 20078 16606 20130
rect 16658 20078 16660 20130
rect 16492 19908 16548 19918
rect 16380 19906 16548 19908
rect 16380 19854 16494 19906
rect 16546 19854 16548 19906
rect 16380 19852 16548 19854
rect 16492 19842 16548 19852
rect 16044 19730 16100 19740
rect 15772 19628 16036 19638
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 15772 19562 16036 19572
rect 15596 19460 15652 19470
rect 15260 19236 15316 19246
rect 15260 19142 15316 19180
rect 15596 19236 15652 19404
rect 16044 19236 16100 19246
rect 16604 19236 16660 20078
rect 17724 20132 17780 20142
rect 17724 20038 17780 20076
rect 16828 20020 16884 20030
rect 17388 20020 17444 20030
rect 15596 19234 16100 19236
rect 15596 19182 15598 19234
rect 15650 19182 16046 19234
rect 16098 19182 16100 19234
rect 15596 19180 16100 19182
rect 15596 19170 15652 19180
rect 16044 19170 16100 19180
rect 16380 19180 16660 19236
rect 16716 20018 17444 20020
rect 16716 19966 16830 20018
rect 16882 19966 17390 20018
rect 17442 19966 17444 20018
rect 16716 19964 17444 19966
rect 15484 19124 15540 19134
rect 15484 19030 15540 19068
rect 15372 19012 15428 19022
rect 15372 18676 15428 18956
rect 16156 19010 16212 19022
rect 16156 18958 16158 19010
rect 16210 18958 16212 19010
rect 15484 18676 15540 18686
rect 15372 18674 15540 18676
rect 15372 18622 15486 18674
rect 15538 18622 15540 18674
rect 15372 18620 15540 18622
rect 15484 18610 15540 18620
rect 15708 18452 15764 18462
rect 15596 18450 15764 18452
rect 15596 18398 15710 18450
rect 15762 18398 15764 18450
rect 15596 18396 15764 18398
rect 15372 18228 15428 18238
rect 15372 18134 15428 18172
rect 15596 17556 15652 18396
rect 15708 18386 15764 18396
rect 16156 18340 16212 18958
rect 15772 18060 16036 18070
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 15772 17994 16036 18004
rect 16156 17892 16212 18284
rect 16156 17826 16212 17836
rect 16156 17666 16212 17678
rect 16156 17614 16158 17666
rect 16210 17614 16212 17666
rect 15932 17556 15988 17566
rect 15596 17500 15932 17556
rect 15932 17462 15988 17500
rect 15260 17332 15316 17342
rect 15148 17276 15260 17332
rect 15260 17266 15316 17276
rect 14812 16482 14868 16492
rect 15772 16492 16036 16502
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 15772 16426 16036 16436
rect 16156 16324 16212 17614
rect 15260 16268 16212 16324
rect 16268 17556 16324 17566
rect 16268 16994 16324 17500
rect 16268 16942 16270 16994
rect 16322 16942 16324 16994
rect 14700 15986 14980 15988
rect 14700 15934 14702 15986
rect 14754 15934 14980 15986
rect 14700 15932 14980 15934
rect 14700 15922 14756 15932
rect 14588 15262 14590 15314
rect 14642 15262 14644 15314
rect 14588 15250 14644 15262
rect 12908 15036 13524 15092
rect 14700 15204 14756 15214
rect 12908 14754 12964 15036
rect 12908 14702 12910 14754
rect 12962 14702 12964 14754
rect 12908 14690 12964 14702
rect 12796 14644 12852 14654
rect 12796 14550 12852 14588
rect 12572 14532 12628 14542
rect 12572 14438 12628 14476
rect 13468 14532 13524 14542
rect 13468 14438 13524 14476
rect 12860 14140 13124 14150
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 12860 14074 13124 14084
rect 14700 13970 14756 15148
rect 14700 13918 14702 13970
rect 14754 13918 14756 13970
rect 14700 13906 14756 13918
rect 14924 14644 14980 15932
rect 12124 13806 12126 13858
rect 12178 13806 12180 13858
rect 12124 13794 12180 13806
rect 14924 13746 14980 14588
rect 14924 13694 14926 13746
rect 14978 13694 14980 13746
rect 14252 13636 14308 13646
rect 14252 13542 14308 13580
rect 14924 13636 14980 13694
rect 14924 13570 14980 13580
rect 13692 13524 13748 13534
rect 13580 12964 13636 12974
rect 13692 12964 13748 13468
rect 14588 13524 14644 13534
rect 14588 13430 14644 13468
rect 14028 13076 14084 13086
rect 14028 12982 14084 13020
rect 14364 13074 14420 13086
rect 14364 13022 14366 13074
rect 14418 13022 14420 13074
rect 13580 12962 13748 12964
rect 13580 12910 13582 12962
rect 13634 12910 13748 12962
rect 13580 12908 13748 12910
rect 13580 12898 13636 12908
rect 12572 12850 12628 12862
rect 12572 12798 12574 12850
rect 12626 12798 12628 12850
rect 12236 12740 12292 12750
rect 12012 12738 12292 12740
rect 12012 12686 12238 12738
rect 12290 12686 12292 12738
rect 12012 12684 12292 12686
rect 12012 12290 12068 12684
rect 12236 12674 12292 12684
rect 12012 12238 12014 12290
rect 12066 12238 12068 12290
rect 12012 12226 12068 12238
rect 12572 11620 12628 12798
rect 12860 12572 13124 12582
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 12860 12506 13124 12516
rect 12572 11554 12628 11564
rect 13580 11620 13636 11630
rect 13580 11526 13636 11564
rect 11900 11284 11956 11294
rect 11900 10834 11956 11228
rect 12860 11004 13124 11014
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 12860 10938 13124 10948
rect 11900 10782 11902 10834
rect 11954 10782 11956 10834
rect 11900 10770 11956 10782
rect 12012 9940 12068 9950
rect 12012 9846 12068 9884
rect 12860 9436 13124 9446
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 12860 9370 13124 9380
rect 12796 9044 12852 9054
rect 12796 8930 12852 8988
rect 12796 8878 12798 8930
rect 12850 8878 12852 8930
rect 12796 8866 12852 8878
rect 11788 8372 12068 8428
rect 12012 8370 12068 8372
rect 12012 8318 12014 8370
rect 12066 8318 12068 8370
rect 12012 8306 12068 8318
rect 11564 8260 11620 8270
rect 11564 8166 11620 8204
rect 13692 8260 13748 12908
rect 14364 12404 14420 13022
rect 15260 13076 15316 16268
rect 16268 16212 16324 16942
rect 15820 16156 16324 16212
rect 15708 15428 15764 15438
rect 15596 15316 15652 15326
rect 15484 15204 15540 15242
rect 15596 15222 15652 15260
rect 15708 15148 15764 15372
rect 15820 15314 15876 16156
rect 15820 15262 15822 15314
rect 15874 15262 15876 15314
rect 15820 15250 15876 15262
rect 16156 15426 16212 15438
rect 16156 15374 16158 15426
rect 16210 15374 16212 15426
rect 15484 15138 15540 15148
rect 15372 15092 15428 15102
rect 15372 13858 15428 15036
rect 15372 13806 15374 13858
rect 15426 13806 15428 13858
rect 15372 13794 15428 13806
rect 15596 15092 15764 15148
rect 15596 13746 15652 15092
rect 15772 14924 16036 14934
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 15772 14858 16036 14868
rect 16156 13860 16212 15374
rect 16380 13972 16436 19180
rect 16492 19010 16548 19022
rect 16492 18958 16494 19010
rect 16546 18958 16548 19010
rect 16492 18452 16548 18958
rect 16604 19010 16660 19022
rect 16604 18958 16606 19010
rect 16658 18958 16660 19010
rect 16604 18900 16660 18958
rect 16604 18834 16660 18844
rect 16492 18386 16548 18396
rect 16492 17892 16548 17902
rect 16716 17892 16772 19964
rect 16828 19954 16884 19964
rect 17388 19954 17444 19964
rect 17388 19796 17444 19806
rect 17164 19236 17220 19246
rect 17164 19142 17220 19180
rect 16828 19012 16884 19022
rect 16828 19010 17108 19012
rect 16828 18958 16830 19010
rect 16882 18958 17108 19010
rect 16828 18956 17108 18958
rect 16828 18946 16884 18956
rect 16492 17890 16772 17892
rect 16492 17838 16494 17890
rect 16546 17838 16772 17890
rect 16492 17836 16772 17838
rect 16492 17826 16548 17836
rect 16828 17556 16884 17566
rect 16828 17462 16884 17500
rect 16940 17444 16996 17454
rect 16940 17350 16996 17388
rect 16828 17332 16884 17342
rect 16604 16882 16660 16894
rect 16604 16830 16606 16882
rect 16658 16830 16660 16882
rect 16492 15876 16548 15886
rect 16492 15538 16548 15820
rect 16492 15486 16494 15538
rect 16546 15486 16548 15538
rect 16492 15474 16548 15486
rect 16604 15428 16660 16830
rect 16716 16100 16772 16110
rect 16828 16100 16884 17276
rect 16716 16098 16884 16100
rect 16716 16046 16718 16098
rect 16770 16046 16884 16098
rect 16716 16044 16884 16046
rect 17052 16660 17108 18956
rect 17388 18564 17444 19740
rect 17500 19236 17556 19246
rect 17836 19236 17892 20748
rect 19292 20802 19348 20814
rect 19292 20750 19294 20802
rect 19346 20750 19348 20802
rect 18684 20412 18948 20422
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18684 20346 18948 20356
rect 17500 19234 17892 19236
rect 17500 19182 17502 19234
rect 17554 19182 17892 19234
rect 17500 19180 17892 19182
rect 17500 19170 17556 19180
rect 17388 18116 17444 18508
rect 17612 18900 17668 18910
rect 17612 18450 17668 18844
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18386 17668 18398
rect 17388 18060 17668 18116
rect 17500 17668 17556 17678
rect 17164 17444 17220 17454
rect 17164 17350 17220 17388
rect 16716 16034 16772 16044
rect 17052 15540 17108 16604
rect 17052 15474 17108 15484
rect 17164 16884 17220 16894
rect 17164 16772 17220 16828
rect 17388 16882 17444 16894
rect 17388 16830 17390 16882
rect 17442 16830 17444 16882
rect 17388 16772 17444 16830
rect 17164 16716 17444 16772
rect 16604 15362 16660 15372
rect 17164 14644 17220 16716
rect 17500 16660 17556 17612
rect 16940 14642 17220 14644
rect 16940 14590 17166 14642
rect 17218 14590 17220 14642
rect 16940 14588 17220 14590
rect 16492 13972 16548 13982
rect 16380 13970 16548 13972
rect 16380 13918 16494 13970
rect 16546 13918 16548 13970
rect 16380 13916 16548 13918
rect 16492 13906 16548 13916
rect 16156 13794 16212 13804
rect 15596 13694 15598 13746
rect 15650 13694 15652 13746
rect 15596 13682 15652 13694
rect 16380 13634 16436 13646
rect 16380 13582 16382 13634
rect 16434 13582 16436 13634
rect 15932 13524 15988 13534
rect 15932 13522 16212 13524
rect 15932 13470 15934 13522
rect 15986 13470 16212 13522
rect 15932 13468 16212 13470
rect 15932 13458 15988 13468
rect 15772 13356 16036 13366
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 15772 13290 16036 13300
rect 15260 13010 15316 13020
rect 14364 12338 14420 12348
rect 15596 12740 15652 12750
rect 15596 12402 15652 12684
rect 15596 12350 15598 12402
rect 15650 12350 15652 12402
rect 15596 12338 15652 12350
rect 15708 12404 15764 12414
rect 14140 12180 14196 12190
rect 14140 12068 14196 12124
rect 15148 12180 15204 12190
rect 15148 12086 15204 12124
rect 15372 12178 15428 12190
rect 15708 12180 15764 12348
rect 15372 12126 15374 12178
rect 15426 12126 15428 12178
rect 13916 12066 14196 12068
rect 13916 12014 14142 12066
rect 14194 12014 14196 12066
rect 13916 12012 14196 12014
rect 13916 11618 13972 12012
rect 14140 12002 14196 12012
rect 15372 11788 15428 12126
rect 15596 12178 15764 12180
rect 15596 12126 15710 12178
rect 15762 12126 15764 12178
rect 15596 12124 15764 12126
rect 15484 12068 15540 12078
rect 15484 11974 15540 12012
rect 13916 11566 13918 11618
rect 13970 11566 13972 11618
rect 13916 11554 13972 11566
rect 15260 11732 15428 11788
rect 14700 11508 14756 11518
rect 14700 11394 14756 11452
rect 14700 11342 14702 11394
rect 14754 11342 14756 11394
rect 14476 11284 14532 11294
rect 14476 11190 14532 11228
rect 14700 9716 14756 11342
rect 15260 10836 15316 11732
rect 15596 11508 15652 12124
rect 15708 12114 15764 12124
rect 16156 12402 16212 13468
rect 16380 12740 16436 13582
rect 16604 13076 16660 13086
rect 16492 12852 16548 12862
rect 16492 12758 16548 12796
rect 16380 12674 16436 12684
rect 16156 12350 16158 12402
rect 16210 12350 16212 12402
rect 15772 11788 16036 11798
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 15772 11722 16036 11732
rect 15596 11442 15652 11452
rect 15036 9826 15092 9838
rect 15036 9774 15038 9826
rect 15090 9774 15092 9826
rect 14812 9716 14868 9726
rect 14700 9714 14868 9716
rect 14700 9662 14814 9714
rect 14866 9662 14868 9714
rect 14700 9660 14868 9662
rect 14812 9268 14868 9660
rect 14812 9202 14868 9212
rect 14924 9602 14980 9614
rect 14924 9550 14926 9602
rect 14978 9550 14980 9602
rect 14924 9154 14980 9550
rect 14924 9102 14926 9154
rect 14978 9102 14980 9154
rect 14924 9090 14980 9102
rect 15036 8428 15092 9774
rect 15260 9826 15316 10780
rect 16044 10836 16100 10846
rect 16156 10836 16212 12350
rect 16492 12404 16548 12414
rect 16492 12310 16548 12348
rect 16044 10834 16212 10836
rect 16044 10782 16046 10834
rect 16098 10782 16212 10834
rect 16044 10780 16212 10782
rect 16492 10836 16548 10846
rect 16044 10770 16100 10780
rect 15260 9774 15262 9826
rect 15314 9774 15316 9826
rect 15260 9762 15316 9774
rect 15596 10498 15652 10510
rect 15596 10446 15598 10498
rect 15650 10446 15652 10498
rect 15596 10388 15652 10446
rect 16380 10388 16436 10398
rect 15596 10386 16436 10388
rect 15596 10334 16382 10386
rect 16434 10334 16436 10386
rect 15596 10332 16436 10334
rect 15484 9044 15540 9054
rect 15036 8372 15316 8428
rect 15372 8372 15428 8382
rect 15260 8370 15428 8372
rect 15260 8318 15374 8370
rect 15426 8318 15428 8370
rect 15260 8316 15428 8318
rect 15372 8306 15428 8316
rect 15484 8370 15540 8988
rect 15484 8318 15486 8370
rect 15538 8318 15540 8370
rect 15484 8306 15540 8318
rect 13916 8260 13972 8270
rect 13748 8258 13972 8260
rect 13748 8206 13918 8258
rect 13970 8206 13972 8258
rect 13748 8204 13972 8206
rect 13692 8194 13748 8204
rect 13916 8194 13972 8204
rect 10444 7970 10500 7980
rect 10892 8148 10948 8158
rect 9660 7756 9996 7812
rect 8988 7410 9044 7420
rect 9100 7588 9156 7598
rect 9100 6916 9156 7532
rect 8988 6914 9156 6916
rect 8988 6862 9102 6914
rect 9154 6862 9156 6914
rect 8988 6860 9156 6862
rect 8092 6580 8148 6590
rect 8092 6486 8148 6524
rect 8764 6580 8820 6590
rect 8764 6486 8820 6524
rect 7756 6468 7812 6478
rect 6860 6466 7812 6468
rect 6860 6414 7758 6466
rect 7810 6414 7812 6466
rect 6860 6412 7812 6414
rect 6860 6018 6916 6412
rect 7756 6402 7812 6412
rect 7036 6300 7300 6310
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7036 6234 7300 6244
rect 6860 5966 6862 6018
rect 6914 5966 6916 6018
rect 6860 5954 6916 5966
rect 6188 5854 6190 5906
rect 6242 5854 6244 5906
rect 6188 5842 6244 5854
rect 5740 5742 5742 5794
rect 5794 5742 5796 5794
rect 5740 5730 5796 5742
rect 8988 5794 9044 6860
rect 9100 6850 9156 6860
rect 9660 6690 9716 7756
rect 9996 7746 10052 7756
rect 10892 7700 10948 8092
rect 10332 7476 10388 7486
rect 10332 7382 10388 7420
rect 10892 7474 10948 7644
rect 11452 8146 11508 8158
rect 11452 8094 11454 8146
rect 11506 8094 11508 8146
rect 11116 7588 11172 7598
rect 11172 7532 11396 7588
rect 11116 7494 11172 7532
rect 10892 7422 10894 7474
rect 10946 7422 10948 7474
rect 10892 7410 10948 7422
rect 9996 7252 10052 7262
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9660 6626 9716 6638
rect 9772 7250 10052 7252
rect 9772 7198 9998 7250
rect 10050 7198 10052 7250
rect 9772 7196 10052 7198
rect 9772 6578 9828 7196
rect 9996 7186 10052 7196
rect 9948 7084 10212 7094
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 9948 7018 10212 7028
rect 9772 6526 9774 6578
rect 9826 6526 9828 6578
rect 9772 6514 9828 6526
rect 8988 5742 8990 5794
rect 9042 5742 9044 5794
rect 8988 5730 9044 5742
rect 11340 5794 11396 7532
rect 11452 7364 11508 8094
rect 13468 8148 13524 8158
rect 13468 8054 13524 8092
rect 12348 8036 12404 8046
rect 12348 8034 12628 8036
rect 12348 7982 12350 8034
rect 12402 7982 12628 8034
rect 12348 7980 12628 7982
rect 12348 7970 12404 7980
rect 12012 7588 12068 7598
rect 12012 7474 12068 7532
rect 12572 7586 12628 7980
rect 12860 7868 13124 7878
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 12860 7802 13124 7812
rect 12572 7534 12574 7586
rect 12626 7534 12628 7586
rect 12572 7522 12628 7534
rect 12796 7588 12852 7598
rect 12012 7422 12014 7474
rect 12066 7422 12068 7474
rect 12012 7410 12068 7422
rect 12796 7474 12852 7532
rect 15484 7588 15540 7598
rect 15596 7588 15652 10332
rect 16380 10322 16436 10332
rect 15772 10220 16036 10230
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 16492 10164 16548 10780
rect 16604 10834 16660 13020
rect 16940 11396 16996 14588
rect 17164 14578 17220 14588
rect 17276 16604 17556 16660
rect 17276 13748 17332 16604
rect 17612 16548 17668 18060
rect 17388 16492 17668 16548
rect 17724 17892 17780 17902
rect 17388 15314 17444 16492
rect 17724 15986 17780 17836
rect 17836 17668 17892 19180
rect 19292 19908 19348 20750
rect 19404 19908 19460 21420
rect 20748 21474 20804 21486
rect 20748 21422 20750 21474
rect 20802 21422 20804 21474
rect 19740 20804 19796 20814
rect 19740 20710 19796 20748
rect 20748 20804 20804 21422
rect 20188 20692 20244 20702
rect 20076 20690 20244 20692
rect 20076 20638 20190 20690
rect 20242 20638 20244 20690
rect 20076 20636 20244 20638
rect 20076 20244 20132 20636
rect 20188 20626 20244 20636
rect 19852 20188 20132 20244
rect 20748 20244 20804 20748
rect 19628 20130 19684 20142
rect 19628 20078 19630 20130
rect 19682 20078 19684 20130
rect 19516 19908 19572 19918
rect 19404 19906 19572 19908
rect 19404 19854 19518 19906
rect 19570 19854 19572 19906
rect 19404 19852 19572 19854
rect 19292 19236 19348 19852
rect 19516 19842 19572 19852
rect 19292 19170 19348 19180
rect 18172 19122 18228 19134
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 18674 18228 19070
rect 18684 18844 18948 18854
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18684 18778 18948 18788
rect 18172 18622 18174 18674
rect 18226 18622 18228 18674
rect 18172 18610 18228 18622
rect 19628 18564 19684 20078
rect 19852 20130 19908 20188
rect 20748 20178 20804 20188
rect 19852 20078 19854 20130
rect 19906 20078 19908 20130
rect 19852 20066 19908 20078
rect 20300 20130 20356 20142
rect 20300 20078 20302 20130
rect 20354 20078 20356 20130
rect 20076 20018 20132 20030
rect 20076 19966 20078 20018
rect 20130 19966 20132 20018
rect 20076 19908 20132 19966
rect 20076 19842 20132 19852
rect 20300 19460 20356 20078
rect 20300 19346 20356 19404
rect 20300 19294 20302 19346
rect 20354 19294 20356 19346
rect 20188 18676 20244 18686
rect 20300 18676 20356 19294
rect 20188 18674 20356 18676
rect 20188 18622 20190 18674
rect 20242 18622 20356 18674
rect 20188 18620 20356 18622
rect 20412 20018 20468 20030
rect 20412 19966 20414 20018
rect 20466 19966 20468 20018
rect 20188 18610 20244 18620
rect 19740 18564 19796 18574
rect 19628 18508 19740 18564
rect 19740 18470 19796 18508
rect 18060 18452 18116 18462
rect 18060 18358 18116 18396
rect 18396 18450 18452 18462
rect 19516 18452 19572 18462
rect 18396 18398 18398 18450
rect 18450 18398 18452 18450
rect 18396 18340 18452 18398
rect 18396 18274 18452 18284
rect 19068 18396 19516 18452
rect 17836 17602 17892 17612
rect 17724 15934 17726 15986
rect 17778 15934 17780 15986
rect 17724 15922 17780 15934
rect 18172 17554 18228 17566
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 17612 15540 17668 15550
rect 17612 15426 17668 15484
rect 18172 15540 18228 17502
rect 19068 17444 19124 18396
rect 19516 18358 19572 18396
rect 20076 18340 20132 18350
rect 20076 18246 20132 18284
rect 20412 18226 20468 19966
rect 20972 18452 21028 18462
rect 21084 18452 21140 21534
rect 21196 21026 21252 22204
rect 21308 22194 21364 22204
rect 23660 22148 23716 22158
rect 23548 21924 23604 21934
rect 21868 21476 21924 21486
rect 21196 20974 21198 21026
rect 21250 20974 21252 21026
rect 21196 20962 21252 20974
rect 21308 21474 21924 21476
rect 21308 21422 21870 21474
rect 21922 21422 21924 21474
rect 21308 21420 21924 21422
rect 20972 18450 21140 18452
rect 20972 18398 20974 18450
rect 21026 18398 21140 18450
rect 20972 18396 21140 18398
rect 21196 20130 21252 20142
rect 21196 20078 21198 20130
rect 21250 20078 21252 20130
rect 21196 18564 21252 20078
rect 21308 20130 21364 21420
rect 21868 21410 21924 21420
rect 21596 21196 21860 21206
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21596 21130 21860 21140
rect 21532 21026 21588 21038
rect 21532 20974 21534 21026
rect 21586 20974 21588 21026
rect 21532 20914 21588 20974
rect 21532 20862 21534 20914
rect 21586 20862 21588 20914
rect 21532 20850 21588 20862
rect 22540 20916 22596 20926
rect 22092 20802 22148 20814
rect 22092 20750 22094 20802
rect 22146 20750 22148 20802
rect 21868 20692 21924 20702
rect 21644 20690 21924 20692
rect 21644 20638 21870 20690
rect 21922 20638 21924 20690
rect 21644 20636 21924 20638
rect 21308 20078 21310 20130
rect 21362 20078 21364 20130
rect 21308 20066 21364 20078
rect 21420 20132 21476 20142
rect 21644 20132 21700 20636
rect 21868 20626 21924 20636
rect 21420 20130 21700 20132
rect 21420 20078 21422 20130
rect 21474 20078 21700 20130
rect 21420 20076 21700 20078
rect 21980 20244 22036 20254
rect 21980 20130 22036 20188
rect 21980 20078 21982 20130
rect 22034 20078 22036 20130
rect 21420 20066 21476 20076
rect 21980 20066 22036 20078
rect 21756 20018 21812 20030
rect 21756 19966 21758 20018
rect 21810 19966 21812 20018
rect 21756 19796 21812 19966
rect 20636 18228 20692 18238
rect 20412 18174 20414 18226
rect 20466 18174 20468 18226
rect 20412 17892 20468 18174
rect 20412 17826 20468 17836
rect 20524 18172 20636 18228
rect 18684 17276 18948 17286
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18684 17210 18948 17220
rect 19068 16100 19124 17388
rect 20300 17778 20356 17790
rect 20300 17726 20302 17778
rect 20354 17726 20356 17778
rect 19068 16098 19684 16100
rect 19068 16046 19070 16098
rect 19122 16046 19684 16098
rect 19068 16044 19684 16046
rect 19068 16034 19124 16044
rect 18284 15876 18340 15886
rect 18284 15782 18340 15820
rect 18732 15876 18788 15886
rect 18732 15874 19124 15876
rect 18732 15822 18734 15874
rect 18786 15822 19124 15874
rect 18732 15820 19124 15822
rect 18732 15810 18788 15820
rect 19068 15764 19124 15820
rect 18684 15708 18948 15718
rect 19068 15708 19236 15764
rect 18172 15474 18228 15484
rect 18508 15652 18564 15662
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18684 15642 18948 15652
rect 18508 15538 18564 15596
rect 18508 15486 18510 15538
rect 18562 15486 18564 15538
rect 18508 15474 18564 15486
rect 17612 15374 17614 15426
rect 17666 15374 17668 15426
rect 17612 15362 17668 15374
rect 18844 15428 18900 15438
rect 18844 15334 18900 15372
rect 17388 15262 17390 15314
rect 17442 15262 17444 15314
rect 17388 15250 17444 15262
rect 17724 15314 17780 15326
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 17500 13748 17556 13758
rect 17276 13692 17500 13748
rect 17276 12962 17332 13692
rect 17500 13654 17556 13692
rect 17724 13524 17780 15262
rect 18172 15090 18228 15102
rect 18172 15038 18174 15090
rect 18226 15038 18228 15090
rect 18172 14532 18228 15038
rect 18172 14466 18228 14476
rect 18172 14308 18228 14318
rect 18172 13858 18228 14252
rect 19068 14308 19124 14318
rect 19068 14214 19124 14252
rect 18684 14140 18948 14150
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18684 14074 18948 14084
rect 18172 13806 18174 13858
rect 18226 13806 18228 13858
rect 18172 13794 18228 13806
rect 17724 13458 17780 13468
rect 18396 13524 18452 13534
rect 18452 13468 18564 13524
rect 18396 13458 18452 13468
rect 17276 12910 17278 12962
rect 17330 12910 17332 12962
rect 17276 12898 17332 12910
rect 17388 12852 17444 12862
rect 17388 12402 17444 12796
rect 17388 12350 17390 12402
rect 17442 12350 17444 12402
rect 17388 12338 17444 12350
rect 18396 12292 18452 12302
rect 18508 12292 18564 13468
rect 19180 12964 19236 15708
rect 19516 15540 19572 15550
rect 19516 15426 19572 15484
rect 19516 15374 19518 15426
rect 19570 15374 19572 15426
rect 19516 15362 19572 15374
rect 19628 15314 19684 16044
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19628 15250 19684 15262
rect 19852 15316 19908 15326
rect 19852 15222 19908 15260
rect 20300 15148 20356 17726
rect 20524 17220 20580 18172
rect 20636 18162 20692 18172
rect 20972 17668 21028 18396
rect 20412 17164 20580 17220
rect 20636 17220 20692 17230
rect 20412 15314 20468 17164
rect 20412 15262 20414 15314
rect 20466 15262 20468 15314
rect 20412 15250 20468 15262
rect 20524 15988 20580 15998
rect 20524 15316 20580 15932
rect 19964 15090 20020 15102
rect 19964 15038 19966 15090
rect 20018 15038 20020 15090
rect 19964 14642 20020 15038
rect 20076 15092 20132 15102
rect 20076 14754 20132 15036
rect 20076 14702 20078 14754
rect 20130 14702 20132 14754
rect 20076 14690 20132 14702
rect 20188 15092 20356 15148
rect 19964 14590 19966 14642
rect 20018 14590 20020 14642
rect 19964 14578 20020 14590
rect 20188 14644 20244 15092
rect 20412 14756 20468 14766
rect 20524 14756 20580 15260
rect 20412 14754 20580 14756
rect 20412 14702 20414 14754
rect 20466 14702 20580 14754
rect 20412 14700 20580 14702
rect 20412 14690 20468 14700
rect 19292 14532 19348 14542
rect 20188 14532 20244 14588
rect 19292 14438 19348 14476
rect 20076 14476 20244 14532
rect 19852 14420 19908 14430
rect 20076 14420 20132 14476
rect 19852 14418 20132 14420
rect 19852 14366 19854 14418
rect 19906 14366 20132 14418
rect 19852 14364 20132 14366
rect 20636 14418 20692 17164
rect 20972 16994 21028 17612
rect 20972 16942 20974 16994
rect 21026 16942 21028 16994
rect 20972 16930 21028 16942
rect 20748 16212 20804 16222
rect 20748 14754 20804 16156
rect 20748 14702 20750 14754
rect 20802 14702 20804 14754
rect 20748 14690 20804 14702
rect 20860 15092 20916 15102
rect 20636 14366 20638 14418
rect 20690 14366 20692 14418
rect 19852 14354 19908 14364
rect 20636 14354 20692 14366
rect 20636 13748 20692 13758
rect 20636 13654 20692 13692
rect 19404 13636 19460 13646
rect 20300 13636 20356 13646
rect 19404 13074 19460 13580
rect 19404 13022 19406 13074
rect 19458 13022 19460 13074
rect 19404 13010 19460 13022
rect 20188 13634 20356 13636
rect 20188 13582 20302 13634
rect 20354 13582 20356 13634
rect 20188 13580 20356 13582
rect 19068 12962 19236 12964
rect 19068 12910 19182 12962
rect 19234 12910 19236 12962
rect 19068 12908 19236 12910
rect 18956 12852 19012 12862
rect 18956 12758 19012 12796
rect 18684 12572 18948 12582
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18684 12506 18948 12516
rect 18396 12290 18564 12292
rect 18396 12238 18398 12290
rect 18450 12238 18564 12290
rect 18396 12236 18564 12238
rect 18956 12292 19012 12302
rect 18396 12226 18452 12236
rect 18956 12178 19012 12236
rect 18956 12126 18958 12178
rect 19010 12126 19012 12178
rect 18956 12114 19012 12126
rect 17500 12068 17556 12078
rect 17500 11974 17556 12012
rect 16940 11302 16996 11340
rect 17500 11284 17556 11294
rect 16604 10782 16606 10834
rect 16658 10782 16660 10834
rect 16604 10770 16660 10782
rect 17388 11282 17556 11284
rect 17388 11230 17502 11282
rect 17554 11230 17556 11282
rect 17388 11228 17556 11230
rect 15772 10154 16036 10164
rect 16268 10108 16548 10164
rect 17388 10610 17444 11228
rect 17500 11218 17556 11228
rect 18684 11004 18948 11014
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18684 10938 18948 10948
rect 17388 10558 17390 10610
rect 17442 10558 17444 10610
rect 17388 10164 17444 10558
rect 16268 9266 16324 10108
rect 16268 9214 16270 9266
rect 16322 9214 16324 9266
rect 16268 9202 16324 9214
rect 16604 9268 16660 9278
rect 16604 9174 16660 9212
rect 15708 9042 15764 9054
rect 15708 8990 15710 9042
rect 15762 8990 15764 9042
rect 15708 8820 15764 8990
rect 16044 9044 16100 9054
rect 16044 8950 16100 8988
rect 16492 9042 16548 9054
rect 16492 8990 16494 9042
rect 16546 8990 16548 9042
rect 15708 8754 15764 8764
rect 16380 8930 16436 8942
rect 16380 8878 16382 8930
rect 16434 8878 16436 8930
rect 15772 8652 16036 8662
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 16380 8596 16436 8878
rect 15772 8586 16036 8596
rect 16156 8540 16436 8596
rect 16156 8484 16212 8540
rect 15820 8428 16212 8484
rect 15820 8370 15876 8428
rect 15820 8318 15822 8370
rect 15874 8318 15876 8370
rect 15820 8306 15876 8318
rect 15932 8036 15988 8046
rect 15932 8034 16100 8036
rect 15932 7982 15934 8034
rect 15986 7982 16100 8034
rect 15932 7980 16100 7982
rect 15932 7970 15988 7980
rect 15540 7532 15652 7588
rect 16044 7586 16100 7980
rect 16044 7534 16046 7586
rect 16098 7534 16100 7586
rect 15484 7522 15540 7532
rect 16044 7522 16100 7534
rect 12796 7422 12798 7474
rect 12850 7422 12852 7474
rect 12796 7410 12852 7422
rect 11452 7298 11508 7308
rect 13916 7364 13972 7374
rect 13916 7270 13972 7308
rect 16492 7364 16548 8990
rect 17388 9042 17444 10108
rect 18172 10498 18228 10510
rect 18172 10446 18174 10498
rect 18226 10446 18228 10498
rect 18172 10050 18228 10446
rect 18172 9998 18174 10050
rect 18226 9998 18228 10050
rect 18172 9986 18228 9998
rect 18284 10052 18340 10062
rect 18284 9716 18340 9996
rect 19068 10052 19124 12908
rect 19180 12898 19236 12908
rect 19852 12962 19908 12974
rect 19852 12910 19854 12962
rect 19906 12910 19908 12962
rect 19516 12850 19572 12862
rect 19516 12798 19518 12850
rect 19570 12798 19572 12850
rect 19292 12066 19348 12078
rect 19292 12014 19294 12066
rect 19346 12014 19348 12066
rect 19292 11732 19348 12014
rect 19292 11666 19348 11676
rect 19516 11508 19572 12798
rect 19740 12292 19796 12302
rect 19852 12292 19908 12910
rect 19796 12236 19908 12292
rect 19964 12850 20020 12862
rect 19964 12798 19966 12850
rect 20018 12798 20020 12850
rect 19964 12740 20020 12798
rect 19740 12198 19796 12236
rect 19516 11442 19572 11452
rect 19068 9986 19124 9996
rect 19964 11396 20020 12684
rect 20076 12180 20132 12190
rect 20188 12180 20244 13580
rect 20300 13570 20356 13580
rect 20860 13186 20916 15036
rect 20860 13134 20862 13186
rect 20914 13134 20916 13186
rect 20860 13122 20916 13134
rect 20300 13076 20356 13086
rect 20300 12850 20356 13020
rect 20300 12798 20302 12850
rect 20354 12798 20356 12850
rect 20300 12786 20356 12798
rect 20524 12962 20580 12974
rect 20524 12910 20526 12962
rect 20578 12910 20580 12962
rect 20132 12124 20244 12180
rect 20076 12086 20132 12124
rect 19964 10388 20020 11340
rect 20524 10836 20580 12910
rect 20524 10770 20580 10780
rect 20636 12292 20692 12302
rect 20300 10498 20356 10510
rect 20300 10446 20302 10498
rect 20354 10446 20356 10498
rect 20300 10388 20356 10446
rect 19964 10332 20356 10388
rect 19852 9828 19908 9838
rect 19964 9828 20020 10332
rect 19852 9826 20020 9828
rect 19852 9774 19854 9826
rect 19906 9774 20020 9826
rect 19852 9772 20020 9774
rect 20076 9828 20132 9838
rect 20412 9828 20468 9838
rect 20076 9826 20468 9828
rect 20076 9774 20078 9826
rect 20130 9774 20414 9826
rect 20466 9774 20468 9826
rect 20076 9772 20468 9774
rect 19852 9762 19908 9772
rect 20076 9762 20132 9772
rect 20412 9762 20468 9772
rect 18508 9716 18564 9726
rect 19180 9716 19236 9726
rect 18284 9714 18452 9716
rect 18284 9662 18286 9714
rect 18338 9662 18452 9714
rect 18284 9660 18452 9662
rect 18284 9650 18340 9660
rect 17388 8990 17390 9042
rect 17442 8990 17444 9042
rect 16492 7298 16548 7308
rect 16828 8820 16884 8830
rect 16828 7474 16884 8764
rect 17388 8820 17444 8990
rect 17388 8754 17444 8764
rect 18172 8930 18228 8942
rect 18172 8878 18174 8930
rect 18226 8878 18228 8930
rect 18172 8482 18228 8878
rect 18172 8430 18174 8482
rect 18226 8430 18228 8482
rect 18172 8418 18228 8430
rect 18396 8428 18452 9660
rect 18508 9714 19236 9716
rect 18508 9662 18510 9714
rect 18562 9662 19182 9714
rect 19234 9662 19236 9714
rect 18508 9660 19236 9662
rect 18508 9650 18564 9660
rect 19180 9650 19236 9660
rect 20636 9714 20692 12236
rect 21196 10948 21252 18508
rect 21420 19740 21812 19796
rect 21868 20020 21924 20030
rect 21868 19796 21924 19964
rect 22092 19906 22148 20750
rect 22540 20802 22596 20860
rect 22540 20750 22542 20802
rect 22594 20750 22596 20802
rect 22540 20738 22596 20750
rect 23212 20692 23268 20702
rect 23212 20598 23268 20636
rect 23212 20244 23268 20254
rect 22092 19854 22094 19906
rect 22146 19854 22148 19906
rect 22092 19842 22148 19854
rect 22204 20130 22260 20142
rect 22204 20078 22206 20130
rect 22258 20078 22260 20130
rect 21868 19740 22036 19796
rect 21308 17892 21364 17902
rect 21420 17892 21476 19740
rect 21596 19628 21860 19638
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21596 19562 21860 19572
rect 21644 19348 21700 19358
rect 21980 19348 22036 19740
rect 22204 19460 22260 20078
rect 23212 20018 23268 20188
rect 23212 19966 23214 20018
rect 23266 19966 23268 20018
rect 23212 19954 23268 19966
rect 23548 20018 23604 21868
rect 23660 20802 23716 22092
rect 24508 21980 24772 21990
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24508 21914 24772 21924
rect 23996 21474 24052 21486
rect 23996 21422 23998 21474
rect 24050 21422 24052 21474
rect 23996 20916 24052 21422
rect 23996 20822 24052 20860
rect 23660 20750 23662 20802
rect 23714 20750 23716 20802
rect 23660 20738 23716 20750
rect 24508 20412 24772 20422
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24508 20346 24772 20356
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 23548 19954 23604 19966
rect 22876 19908 22932 19918
rect 22876 19814 22932 19852
rect 24108 19906 24164 19918
rect 24108 19854 24110 19906
rect 24162 19854 24164 19906
rect 22260 19404 22708 19460
rect 22204 19366 22260 19404
rect 21644 19346 22036 19348
rect 21644 19294 21646 19346
rect 21698 19294 22036 19346
rect 21644 19292 22036 19294
rect 21644 19282 21700 19292
rect 21980 19234 22036 19292
rect 22540 19236 22596 19246
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21980 19170 22036 19182
rect 22092 19234 22596 19236
rect 22092 19182 22542 19234
rect 22594 19182 22596 19234
rect 22092 19180 22596 19182
rect 21756 18340 21812 18350
rect 21756 18338 22036 18340
rect 21756 18286 21758 18338
rect 21810 18286 22036 18338
rect 21756 18284 22036 18286
rect 21756 18274 21812 18284
rect 21596 18060 21860 18070
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21596 17994 21860 18004
rect 21364 17836 21476 17892
rect 21980 17892 22036 18284
rect 22092 18228 22148 19180
rect 22540 19170 22596 19180
rect 22652 19234 22708 19404
rect 22652 19182 22654 19234
rect 22706 19182 22708 19234
rect 22652 19170 22708 19182
rect 22988 19234 23044 19246
rect 22988 19182 22990 19234
rect 23042 19182 23044 19234
rect 22204 19010 22260 19022
rect 22988 19012 23044 19182
rect 23884 19012 23940 19022
rect 22204 18958 22206 19010
rect 22258 18958 22260 19010
rect 22204 18900 22260 18958
rect 22764 18956 23044 19012
rect 23772 19010 23940 19012
rect 23772 18958 23886 19010
rect 23938 18958 23940 19010
rect 23772 18956 23940 18958
rect 22764 18900 22820 18956
rect 22204 18844 22820 18900
rect 22092 18162 22148 18172
rect 22316 18452 22372 18462
rect 22204 17892 22260 17902
rect 21980 17890 22260 17892
rect 21980 17838 22206 17890
rect 22258 17838 22260 17890
rect 21980 17836 22260 17838
rect 21308 17798 21364 17836
rect 22204 17826 22260 17836
rect 22316 17890 22372 18396
rect 22316 17838 22318 17890
rect 22370 17838 22372 17890
rect 22316 17826 22372 17838
rect 22652 17892 22708 17902
rect 22652 17798 22708 17836
rect 21644 17668 21700 17678
rect 21420 17666 21700 17668
rect 21420 17614 21646 17666
rect 21698 17614 21700 17666
rect 21420 17612 21700 17614
rect 21420 16884 21476 17612
rect 21644 17602 21700 17612
rect 21868 17666 21924 17678
rect 22540 17668 22596 17678
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21868 17220 21924 17614
rect 21868 17154 21924 17164
rect 22428 17666 22596 17668
rect 22428 17614 22542 17666
rect 22594 17614 22596 17666
rect 22428 17612 22596 17614
rect 21308 16828 21476 16884
rect 21980 16884 22036 16894
rect 21308 16322 21364 16828
rect 21308 16270 21310 16322
rect 21362 16270 21364 16322
rect 21308 15988 21364 16270
rect 21308 15922 21364 15932
rect 21420 16660 21476 16670
rect 21420 15538 21476 16604
rect 21596 16492 21860 16502
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21596 16426 21860 16436
rect 21420 15486 21422 15538
rect 21474 15486 21476 15538
rect 21420 14756 21476 15486
rect 21644 16098 21700 16110
rect 21644 16046 21646 16098
rect 21698 16046 21700 16098
rect 21532 15426 21588 15438
rect 21532 15374 21534 15426
rect 21586 15374 21588 15426
rect 21532 15092 21588 15374
rect 21644 15204 21700 16046
rect 21868 16100 21924 16110
rect 21868 16006 21924 16044
rect 21644 15138 21700 15148
rect 21532 15026 21588 15036
rect 21596 14924 21860 14934
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21596 14858 21860 14868
rect 21420 14700 21812 14756
rect 21756 14418 21812 14700
rect 21756 14366 21758 14418
rect 21810 14366 21812 14418
rect 21756 14354 21812 14366
rect 21532 14308 21588 14318
rect 21532 14214 21588 14252
rect 21980 14306 22036 16828
rect 22428 16212 22484 17612
rect 22540 17602 22596 17612
rect 23212 17666 23268 17678
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 23100 17556 23156 17566
rect 22764 17554 23156 17556
rect 22764 17502 23102 17554
rect 23154 17502 23156 17554
rect 22764 17500 23156 17502
rect 22764 16772 22820 17500
rect 23100 17490 23156 17500
rect 23212 17220 23268 17614
rect 23772 17666 23828 18956
rect 23884 18946 23940 18956
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23772 17602 23828 17614
rect 23884 18338 23940 18350
rect 23884 18286 23886 18338
rect 23938 18286 23940 18338
rect 23212 17154 23268 17164
rect 23884 17220 23940 18286
rect 23884 17154 23940 17164
rect 22428 16146 22484 16156
rect 22540 16716 22820 16772
rect 22876 16882 22932 16894
rect 22876 16830 22878 16882
rect 22930 16830 22932 16882
rect 22540 15986 22596 16716
rect 22876 16660 22932 16830
rect 23100 16884 23156 16894
rect 23100 16790 23156 16828
rect 23436 16882 23492 16894
rect 23436 16830 23438 16882
rect 23490 16830 23492 16882
rect 22876 16594 22932 16604
rect 23436 16324 23492 16830
rect 22540 15934 22542 15986
rect 22594 15934 22596 15986
rect 22540 15922 22596 15934
rect 22652 16268 23492 16324
rect 22652 15764 22708 16268
rect 23436 16210 23492 16268
rect 23436 16158 23438 16210
rect 23490 16158 23492 16210
rect 23436 16146 23492 16158
rect 23548 16882 23604 16894
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 22316 15708 22708 15764
rect 23212 16098 23268 16110
rect 23212 16046 23214 16098
rect 23266 16046 23268 16098
rect 22092 15428 22148 15438
rect 22092 14754 22148 15372
rect 22092 14702 22094 14754
rect 22146 14702 22148 14754
rect 22092 14690 22148 14702
rect 22316 14530 22372 15708
rect 22988 15428 23044 15438
rect 22988 15334 23044 15372
rect 22316 14478 22318 14530
rect 22370 14478 22372 14530
rect 22316 14466 22372 14478
rect 22428 15092 22484 15102
rect 21980 14254 21982 14306
rect 22034 14254 22036 14306
rect 21420 13636 21476 13646
rect 21420 13542 21476 13580
rect 21596 13356 21860 13366
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21596 13290 21860 13300
rect 21868 12850 21924 12862
rect 21868 12798 21870 12850
rect 21922 12798 21924 12850
rect 21308 12738 21364 12750
rect 21308 12686 21310 12738
rect 21362 12686 21364 12738
rect 21308 12068 21364 12686
rect 21420 12738 21476 12750
rect 21420 12686 21422 12738
rect 21474 12686 21476 12738
rect 21420 12292 21476 12686
rect 21644 12740 21700 12750
rect 21644 12646 21700 12684
rect 21420 12226 21476 12236
rect 21644 12292 21700 12302
rect 21644 12198 21700 12236
rect 21308 12012 21476 12068
rect 21308 11508 21364 11518
rect 21308 11414 21364 11452
rect 21420 11394 21476 12012
rect 21868 11956 21924 12798
rect 21980 12402 22036 14254
rect 21980 12350 21982 12402
rect 22034 12350 22036 12402
rect 21980 12338 22036 12350
rect 22092 13076 22148 13086
rect 22092 12180 22148 13020
rect 22428 13074 22484 15036
rect 22652 14644 22708 14654
rect 22652 14550 22708 14588
rect 23100 14530 23156 14542
rect 23100 14478 23102 14530
rect 23154 14478 23156 14530
rect 23100 14420 23156 14478
rect 23100 14354 23156 14364
rect 22428 13022 22430 13074
rect 22482 13022 22484 13074
rect 22428 13010 22484 13022
rect 23100 13860 23156 13870
rect 23100 12962 23156 13804
rect 23100 12910 23102 12962
rect 23154 12910 23156 12962
rect 23100 12898 23156 12910
rect 23100 12740 23156 12750
rect 21868 11890 21924 11900
rect 21980 12124 22148 12180
rect 22204 12404 22260 12414
rect 22204 12178 22260 12348
rect 22204 12126 22206 12178
rect 22258 12126 22260 12178
rect 21596 11788 21860 11798
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21596 11722 21860 11732
rect 21420 11342 21422 11394
rect 21474 11342 21476 11394
rect 21420 11330 21476 11342
rect 21980 11394 22036 12124
rect 22204 12114 22260 12126
rect 22540 12292 22596 12302
rect 22092 11956 22148 11966
rect 22148 11900 22372 11956
rect 22092 11890 22148 11900
rect 21980 11342 21982 11394
rect 22034 11342 22036 11394
rect 21980 11330 22036 11342
rect 21196 10892 21924 10948
rect 20860 10722 20916 10734
rect 20860 10670 20862 10722
rect 20914 10670 20916 10722
rect 20748 10612 20804 10622
rect 20748 9826 20804 10556
rect 20748 9774 20750 9826
rect 20802 9774 20804 9826
rect 20748 9762 20804 9774
rect 20636 9662 20638 9714
rect 20690 9662 20692 9714
rect 20636 9650 20692 9662
rect 20860 9492 20916 10670
rect 20972 10612 21028 10622
rect 21644 10612 21700 10622
rect 20972 10610 21700 10612
rect 20972 10558 20974 10610
rect 21026 10558 21646 10610
rect 21698 10558 21700 10610
rect 20972 10556 21700 10558
rect 20972 10546 21028 10556
rect 21644 10546 21700 10556
rect 21756 10612 21812 10622
rect 21084 10388 21140 10398
rect 18684 9436 18948 9446
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 20860 9426 20916 9436
rect 20972 10386 21140 10388
rect 20972 10334 21086 10386
rect 21138 10334 21140 10386
rect 20972 10332 21140 10334
rect 18684 9370 18948 9380
rect 19740 9044 19796 9054
rect 18508 8484 18564 8504
rect 18396 8372 18564 8428
rect 18508 8370 18564 8372
rect 18508 8318 18510 8370
rect 18562 8318 18564 8370
rect 18508 8306 18564 8318
rect 19628 8484 19684 8494
rect 16828 7422 16830 7474
rect 16882 7422 16884 7474
rect 11676 7250 11732 7262
rect 11676 7198 11678 7250
rect 11730 7198 11732 7250
rect 11676 6692 11732 7198
rect 15772 7084 16036 7094
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 15772 7018 16036 7028
rect 11788 6692 11844 6702
rect 11676 6690 11844 6692
rect 11676 6638 11790 6690
rect 11842 6638 11844 6690
rect 11676 6636 11844 6638
rect 11788 6626 11844 6636
rect 16828 6692 16884 7422
rect 18284 8036 18340 8046
rect 18284 7474 18340 7980
rect 19516 8034 19572 8046
rect 19516 7982 19518 8034
rect 19570 7982 19572 8034
rect 19516 7924 19572 7982
rect 18684 7868 18948 7878
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 19516 7858 19572 7868
rect 18684 7802 18948 7812
rect 19628 7700 19684 8428
rect 19740 8258 19796 8988
rect 20300 9044 20356 9054
rect 20300 8930 20356 8988
rect 20300 8878 20302 8930
rect 20354 8878 20356 8930
rect 20300 8866 20356 8878
rect 20972 8372 21028 10332
rect 21084 10322 21140 10332
rect 21532 10388 21588 10398
rect 21756 10388 21812 10556
rect 21532 10386 21812 10388
rect 21532 10334 21534 10386
rect 21586 10334 21812 10386
rect 21532 10332 21812 10334
rect 21868 10610 21924 10892
rect 22092 10836 22148 10846
rect 22148 10780 22260 10836
rect 22092 10770 22148 10780
rect 21868 10558 21870 10610
rect 21922 10558 21924 10610
rect 21868 10388 21924 10558
rect 21532 10322 21588 10332
rect 21868 10322 21924 10332
rect 21980 10388 22036 10398
rect 21980 10386 22148 10388
rect 21980 10334 21982 10386
rect 22034 10334 22148 10386
rect 21980 10332 22148 10334
rect 21980 10322 22036 10332
rect 21596 10220 21860 10230
rect 21308 10164 21364 10174
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21596 10154 21860 10164
rect 21980 10164 22036 10174
rect 21308 9826 21364 10108
rect 21308 9774 21310 9826
rect 21362 9774 21364 9826
rect 21308 9762 21364 9774
rect 21644 9492 21700 9502
rect 21084 9044 21140 9054
rect 21084 8950 21140 8988
rect 21308 9042 21364 9054
rect 21308 8990 21310 9042
rect 21362 8990 21364 9042
rect 21308 8484 21364 8990
rect 21420 9042 21476 9054
rect 21420 8990 21422 9042
rect 21474 8990 21476 9042
rect 21420 8596 21476 8990
rect 21644 9042 21700 9436
rect 21644 8990 21646 9042
rect 21698 8990 21700 9042
rect 21644 8978 21700 8990
rect 21596 8652 21860 8662
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21596 8586 21860 8596
rect 21420 8530 21476 8540
rect 19740 8206 19742 8258
rect 19794 8206 19796 8258
rect 19740 8194 19796 8206
rect 20076 8258 20132 8270
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 20076 8148 20132 8206
rect 19740 7700 19796 7710
rect 19628 7698 19796 7700
rect 19628 7646 19742 7698
rect 19794 7646 19796 7698
rect 19628 7644 19796 7646
rect 19740 7634 19796 7644
rect 18284 7422 18286 7474
rect 18338 7422 18340 7474
rect 18284 7410 18340 7422
rect 18956 7476 19012 7486
rect 18956 7382 19012 7420
rect 19180 7476 19236 7486
rect 19516 7476 19572 7486
rect 19180 7474 19572 7476
rect 19180 7422 19182 7474
rect 19234 7422 19518 7474
rect 19570 7422 19572 7474
rect 19180 7420 19572 7422
rect 19180 7410 19236 7420
rect 19516 7410 19572 7420
rect 20076 7476 20132 8092
rect 20524 8146 20580 8158
rect 20524 8094 20526 8146
rect 20578 8094 20580 8146
rect 20412 8036 20468 8046
rect 20412 7942 20468 7980
rect 20524 7924 20580 8094
rect 20524 7858 20580 7868
rect 20748 8146 20804 8158
rect 20748 8094 20750 8146
rect 20802 8094 20804 8146
rect 20748 7812 20804 8094
rect 20748 7746 20804 7756
rect 20076 7410 20132 7420
rect 20524 7476 20580 7486
rect 19628 7362 19684 7374
rect 19628 7310 19630 7362
rect 19682 7310 19684 7362
rect 19628 6916 19684 7310
rect 18508 6860 19684 6916
rect 18508 6802 18564 6860
rect 18508 6750 18510 6802
rect 18562 6750 18564 6802
rect 18508 6738 18564 6750
rect 12012 6468 12068 6478
rect 12012 6374 12068 6412
rect 13468 6468 13524 6478
rect 12860 6300 13124 6310
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 12860 6234 13124 6244
rect 13468 6018 13524 6412
rect 13468 5966 13470 6018
rect 13522 5966 13524 6018
rect 13468 5954 13524 5966
rect 14252 5908 14308 5918
rect 14252 5814 14308 5852
rect 16828 5908 16884 6636
rect 17724 6692 17780 6702
rect 17724 6598 17780 6636
rect 18684 6300 18948 6310
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18684 6234 18948 6244
rect 20524 6132 20580 7420
rect 20972 7476 21028 8316
rect 21084 8428 21364 8484
rect 21644 8484 21700 8494
rect 21980 8484 22036 10108
rect 22092 9938 22148 10332
rect 22092 9886 22094 9938
rect 22146 9886 22148 9938
rect 22092 9874 22148 9886
rect 22092 9268 22148 9278
rect 22204 9268 22260 10780
rect 22316 10834 22372 11900
rect 22540 11060 22596 12236
rect 22652 12180 22708 12190
rect 22652 12178 22932 12180
rect 22652 12126 22654 12178
rect 22706 12126 22932 12178
rect 22652 12124 22932 12126
rect 22652 12114 22708 12124
rect 22764 11396 22820 11406
rect 22764 11302 22820 11340
rect 22540 11004 22820 11060
rect 22316 10782 22318 10834
rect 22370 10782 22372 10834
rect 22316 10612 22372 10782
rect 22316 10546 22372 10556
rect 22540 10836 22596 10846
rect 22540 10610 22596 10780
rect 22540 10558 22542 10610
rect 22594 10558 22596 10610
rect 22540 10546 22596 10558
rect 22092 9266 22260 9268
rect 22092 9214 22094 9266
rect 22146 9214 22260 9266
rect 22092 9212 22260 9214
rect 22092 9202 22148 9212
rect 21084 8148 21140 8428
rect 21084 8082 21140 8092
rect 21420 8146 21476 8158
rect 21420 8094 21422 8146
rect 21474 8094 21476 8146
rect 20972 7410 21028 7420
rect 21308 8036 21364 8046
rect 21308 7474 21364 7980
rect 21420 7924 21476 8094
rect 21532 8148 21588 8158
rect 21532 8054 21588 8092
rect 21644 8146 21700 8428
rect 21644 8094 21646 8146
rect 21698 8094 21700 8146
rect 21420 7858 21476 7868
rect 21644 7812 21700 8094
rect 21644 7746 21700 7756
rect 21756 8428 22036 8484
rect 21308 7422 21310 7474
rect 21362 7422 21364 7474
rect 21308 7410 21364 7422
rect 21420 7476 21476 7486
rect 21420 7382 21476 7420
rect 21644 7476 21700 7486
rect 21756 7476 21812 8428
rect 22092 8372 22148 8382
rect 22092 8278 22148 8316
rect 22652 7700 22708 7710
rect 22316 7588 22372 7598
rect 22652 7588 22708 7644
rect 22316 7586 22708 7588
rect 22316 7534 22318 7586
rect 22370 7534 22708 7586
rect 22316 7532 22708 7534
rect 22316 7522 22372 7532
rect 21644 7474 21812 7476
rect 21644 7422 21646 7474
rect 21698 7422 21812 7474
rect 21644 7420 21812 7422
rect 22652 7474 22708 7532
rect 22652 7422 22654 7474
rect 22706 7422 22708 7474
rect 21644 7410 21700 7420
rect 22652 7410 22708 7422
rect 21756 7252 21812 7262
rect 21756 7250 22036 7252
rect 21756 7198 21758 7250
rect 21810 7198 22036 7250
rect 21756 7196 22036 7198
rect 21756 7186 21812 7196
rect 21596 7084 21860 7094
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21596 7018 21860 7028
rect 20636 6804 20692 6814
rect 20636 6802 20804 6804
rect 20636 6750 20638 6802
rect 20690 6750 20804 6802
rect 20636 6748 20804 6750
rect 20636 6738 20692 6748
rect 20636 6132 20692 6142
rect 20524 6130 20692 6132
rect 20524 6078 20638 6130
rect 20690 6078 20692 6130
rect 20524 6076 20692 6078
rect 20636 6066 20692 6076
rect 20748 5908 20804 6748
rect 21308 6692 21364 6702
rect 21980 6692 22036 7196
rect 22092 6692 22148 6702
rect 21980 6690 22148 6692
rect 21980 6638 22094 6690
rect 22146 6638 22148 6690
rect 21980 6636 22148 6638
rect 21308 6598 21364 6636
rect 22092 6626 22148 6636
rect 20972 5908 21028 5918
rect 20748 5906 21028 5908
rect 20748 5854 20974 5906
rect 21026 5854 21028 5906
rect 20748 5852 21028 5854
rect 16828 5842 16884 5852
rect 11340 5742 11342 5794
rect 11394 5742 11396 5794
rect 11340 5730 11396 5742
rect 4124 5516 4388 5526
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4124 5450 4388 5460
rect 9948 5516 10212 5526
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 9948 5450 10212 5460
rect 15772 5516 16036 5526
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 15772 5450 16036 5460
rect 20972 5236 21028 5852
rect 22764 5684 22820 11004
rect 22876 9154 22932 12124
rect 23100 11394 23156 12684
rect 23100 11342 23102 11394
rect 23154 11342 23156 11394
rect 23100 11330 23156 11342
rect 23100 10724 23156 10734
rect 23212 10724 23268 16046
rect 23324 16100 23380 16110
rect 23324 14644 23380 16044
rect 23548 15876 23604 16830
rect 23996 16658 24052 16670
rect 23996 16606 23998 16658
rect 24050 16606 24052 16658
rect 23996 16324 24052 16606
rect 23996 16258 24052 16268
rect 24108 15986 24164 19854
rect 24220 19908 24276 19918
rect 24220 19122 24276 19852
rect 24220 19070 24222 19122
rect 24274 19070 24276 19122
rect 24220 18004 24276 19070
rect 24508 18844 24772 18854
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24508 18778 24772 18788
rect 24220 17938 24276 17948
rect 24508 17276 24772 17286
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24508 17210 24772 17220
rect 24108 15934 24110 15986
rect 24162 15934 24164 15986
rect 24108 15922 24164 15934
rect 24220 16098 24276 16110
rect 24220 16046 24222 16098
rect 24274 16046 24276 16098
rect 23548 15810 23604 15820
rect 24108 15314 24164 15326
rect 24108 15262 24110 15314
rect 24162 15262 24164 15314
rect 24108 15148 24164 15262
rect 23324 14578 23380 14588
rect 23548 15092 24164 15148
rect 23548 14642 23604 15092
rect 24220 14644 24276 16046
rect 23548 14590 23550 14642
rect 23602 14590 23604 14642
rect 23548 14578 23604 14590
rect 24108 14588 24276 14644
rect 24332 15988 24388 15998
rect 23884 14420 23940 14430
rect 23884 14326 23940 14364
rect 23884 13860 23940 13870
rect 23884 13766 23940 13804
rect 23548 13634 23604 13646
rect 23548 13582 23550 13634
rect 23602 13582 23604 13634
rect 23324 13076 23380 13086
rect 23548 13076 23604 13582
rect 23380 13020 23604 13076
rect 23324 12982 23380 13020
rect 23884 12740 23940 12750
rect 23884 12646 23940 12684
rect 23660 12290 23716 12302
rect 23660 12238 23662 12290
rect 23714 12238 23716 12290
rect 23100 10722 23268 10724
rect 23100 10670 23102 10722
rect 23154 10670 23268 10722
rect 23100 10668 23268 10670
rect 23548 12180 23604 12190
rect 23100 10658 23156 10668
rect 23548 10498 23604 12124
rect 23660 11506 23716 12238
rect 23660 11454 23662 11506
rect 23714 11454 23716 11506
rect 23660 11442 23716 11454
rect 23548 10446 23550 10498
rect 23602 10446 23604 10498
rect 23548 10434 23604 10446
rect 23772 10610 23828 10622
rect 23772 10558 23774 10610
rect 23826 10558 23828 10610
rect 22876 9102 22878 9154
rect 22930 9102 22932 9154
rect 22876 9090 22932 9102
rect 23324 9044 23380 9054
rect 23324 8950 23380 8988
rect 23660 8930 23716 8942
rect 23660 8878 23662 8930
rect 23714 8878 23716 8930
rect 23436 8260 23492 8270
rect 22988 8258 23492 8260
rect 22988 8206 23438 8258
rect 23490 8206 23492 8258
rect 22988 8204 23492 8206
rect 22876 8036 22932 8046
rect 22876 7942 22932 7980
rect 22876 7700 22932 7710
rect 22988 7700 23044 8204
rect 23436 8194 23492 8204
rect 22876 7698 23044 7700
rect 22876 7646 22878 7698
rect 22930 7646 23044 7698
rect 22876 7644 23044 7646
rect 23324 8036 23380 8046
rect 22876 7634 22932 7644
rect 22876 7476 22932 7486
rect 22876 6130 22932 7420
rect 22876 6078 22878 6130
rect 22930 6078 22932 6130
rect 22876 6066 22932 6078
rect 23324 7474 23380 7980
rect 23324 7422 23326 7474
rect 23378 7422 23380 7474
rect 22988 6020 23044 6030
rect 23044 5964 23156 6020
rect 22988 5954 23044 5964
rect 23100 5906 23156 5964
rect 23100 5854 23102 5906
rect 23154 5854 23156 5906
rect 23100 5842 23156 5854
rect 23324 5908 23380 7422
rect 23324 5842 23380 5852
rect 23548 7586 23604 7598
rect 23548 7534 23550 7586
rect 23602 7534 23604 7586
rect 23548 5906 23604 7534
rect 23548 5854 23550 5906
rect 23602 5854 23604 5906
rect 23548 5842 23604 5854
rect 22764 5628 23156 5684
rect 21596 5516 21860 5526
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21596 5450 21860 5460
rect 20972 5170 21028 5180
rect 23100 5234 23156 5628
rect 23100 5182 23102 5234
rect 23154 5182 23156 5234
rect 23100 5170 23156 5182
rect 23548 5236 23604 5246
rect 23548 5142 23604 5180
rect 23660 4900 23716 8878
rect 23772 7700 23828 10558
rect 23884 9492 23940 9502
rect 23884 8258 23940 9436
rect 24108 8370 24164 14588
rect 24220 14420 24276 14430
rect 24332 14420 24388 15932
rect 24508 15708 24772 15718
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24508 15642 24772 15652
rect 24220 14418 24388 14420
rect 24220 14366 24222 14418
rect 24274 14366 24388 14418
rect 24220 14364 24388 14366
rect 24220 14308 24276 14364
rect 24220 14242 24276 14252
rect 24508 14140 24772 14150
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24508 14074 24772 14084
rect 24220 13972 24276 13982
rect 24220 13860 24276 13916
rect 24220 13858 24388 13860
rect 24220 13806 24222 13858
rect 24274 13806 24388 13858
rect 24220 13804 24388 13806
rect 24220 13794 24276 13804
rect 24220 12852 24276 12862
rect 24220 11956 24276 12796
rect 24220 11890 24276 11900
rect 24332 11506 24388 13804
rect 24508 12572 24772 12582
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24508 12506 24772 12516
rect 24332 11454 24334 11506
rect 24386 11454 24388 11506
rect 24332 11442 24388 11454
rect 24508 11004 24772 11014
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24508 10938 24772 10948
rect 24220 9938 24276 9950
rect 24220 9886 24222 9938
rect 24274 9886 24276 9938
rect 24220 9492 24276 9886
rect 24220 9426 24276 9436
rect 24332 9940 24388 9950
rect 24108 8318 24110 8370
rect 24162 8318 24164 8370
rect 24108 8306 24164 8318
rect 23884 8206 23886 8258
rect 23938 8206 23940 8258
rect 23884 8194 23940 8206
rect 24108 7812 24164 7822
rect 23884 7700 23940 7710
rect 23772 7698 23940 7700
rect 23772 7646 23886 7698
rect 23938 7646 23940 7698
rect 23772 7644 23940 7646
rect 23884 7634 23940 7644
rect 24108 6804 24164 7756
rect 24220 7588 24276 7598
rect 24332 7588 24388 9884
rect 24508 9436 24772 9446
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24508 9370 24772 9380
rect 24508 7868 24772 7878
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24508 7802 24772 7812
rect 24220 7586 24388 7588
rect 24220 7534 24222 7586
rect 24274 7534 24388 7586
rect 24220 7532 24388 7534
rect 24220 7476 24276 7532
rect 24220 7410 24276 7420
rect 24220 6804 24276 6814
rect 24108 6802 24276 6804
rect 24108 6750 24222 6802
rect 24274 6750 24276 6802
rect 24108 6748 24276 6750
rect 23996 5908 24052 5918
rect 24220 5908 24276 6748
rect 24508 6300 24772 6310
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24508 6234 24772 6244
rect 23996 5906 24276 5908
rect 23996 5854 23998 5906
rect 24050 5854 24276 5906
rect 23996 5852 24276 5854
rect 23996 5842 24052 5852
rect 23772 5124 23828 5134
rect 23772 5122 23940 5124
rect 23772 5070 23774 5122
rect 23826 5070 23940 5122
rect 23772 5068 23940 5070
rect 23772 5058 23828 5068
rect 23548 4844 23716 4900
rect 7036 4732 7300 4742
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7036 4666 7300 4676
rect 12860 4732 13124 4742
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 12860 4666 13124 4676
rect 18684 4732 18948 4742
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18684 4666 18948 4676
rect 4124 3948 4388 3958
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4124 3882 4388 3892
rect 9948 3948 10212 3958
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 9948 3882 10212 3892
rect 15772 3948 16036 3958
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 15772 3882 16036 3892
rect 21596 3948 21860 3958
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21596 3882 21860 3892
rect 23436 3444 23492 3482
rect 23548 3444 23604 4844
rect 23884 4562 23940 5068
rect 24508 4732 24772 4742
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24508 4666 24772 4676
rect 23884 4510 23886 4562
rect 23938 4510 23940 4562
rect 23884 4498 23940 4510
rect 24220 4338 24276 4350
rect 24220 4286 24222 4338
rect 24274 4286 24276 4338
rect 23660 4228 23716 4238
rect 24220 4228 24276 4286
rect 23660 4226 24276 4228
rect 23660 4174 23662 4226
rect 23714 4174 24276 4226
rect 23660 4172 24276 4174
rect 23660 4162 23716 4172
rect 24220 3892 24276 4172
rect 24220 3826 24276 3836
rect 23660 3444 23716 3454
rect 23548 3442 23716 3444
rect 23548 3390 23662 3442
rect 23714 3390 23716 3442
rect 23548 3388 23716 3390
rect 23436 3378 23492 3388
rect 23660 3378 23716 3388
rect 23884 3444 23940 3454
rect 23996 3444 24052 3482
rect 23940 3442 24052 3444
rect 23940 3390 23998 3442
rect 24050 3390 24052 3442
rect 23940 3388 24052 3390
rect 23884 3378 23940 3388
rect 7036 3164 7300 3174
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7036 3098 7300 3108
rect 12860 3164 13124 3174
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 12860 3098 13124 3108
rect 18684 3164 18948 3174
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18684 3098 18948 3108
rect 23996 1876 24052 3388
rect 24508 3164 24772 3174
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24508 3098 24772 3108
rect 23996 1810 24052 1820
<< via2 >>
rect 3500 20076 3556 20132
rect 1820 19234 1876 19236
rect 1820 19182 1822 19234
rect 1822 19182 1874 19234
rect 1874 19182 1876 19234
rect 1820 19180 1876 19182
rect 4124 22762 4180 22764
rect 4124 22710 4126 22762
rect 4126 22710 4178 22762
rect 4178 22710 4180 22762
rect 4124 22708 4180 22710
rect 4228 22762 4284 22764
rect 4228 22710 4230 22762
rect 4230 22710 4282 22762
rect 4282 22710 4284 22762
rect 4228 22708 4284 22710
rect 4332 22762 4388 22764
rect 4332 22710 4334 22762
rect 4334 22710 4386 22762
rect 4386 22710 4388 22762
rect 4332 22708 4388 22710
rect 9948 22762 10004 22764
rect 9948 22710 9950 22762
rect 9950 22710 10002 22762
rect 10002 22710 10004 22762
rect 9948 22708 10004 22710
rect 10052 22762 10108 22764
rect 10052 22710 10054 22762
rect 10054 22710 10106 22762
rect 10106 22710 10108 22762
rect 10052 22708 10108 22710
rect 10156 22762 10212 22764
rect 10156 22710 10158 22762
rect 10158 22710 10210 22762
rect 10210 22710 10212 22762
rect 10156 22708 10212 22710
rect 20300 23996 20356 24052
rect 15772 22762 15828 22764
rect 15772 22710 15774 22762
rect 15774 22710 15826 22762
rect 15826 22710 15828 22762
rect 15772 22708 15828 22710
rect 15876 22762 15932 22764
rect 15876 22710 15878 22762
rect 15878 22710 15930 22762
rect 15930 22710 15932 22762
rect 15876 22708 15932 22710
rect 15980 22762 16036 22764
rect 15980 22710 15982 22762
rect 15982 22710 16034 22762
rect 16034 22710 16036 22762
rect 15980 22708 16036 22710
rect 17500 22316 17556 22372
rect 7036 21978 7092 21980
rect 7036 21926 7038 21978
rect 7038 21926 7090 21978
rect 7090 21926 7092 21978
rect 7036 21924 7092 21926
rect 7140 21978 7196 21980
rect 7140 21926 7142 21978
rect 7142 21926 7194 21978
rect 7194 21926 7196 21978
rect 7140 21924 7196 21926
rect 7244 21978 7300 21980
rect 7244 21926 7246 21978
rect 7246 21926 7298 21978
rect 7298 21926 7300 21978
rect 7244 21924 7300 21926
rect 12860 21978 12916 21980
rect 12860 21926 12862 21978
rect 12862 21926 12914 21978
rect 12914 21926 12916 21978
rect 12860 21924 12916 21926
rect 12964 21978 13020 21980
rect 12964 21926 12966 21978
rect 12966 21926 13018 21978
rect 13018 21926 13020 21978
rect 12964 21924 13020 21926
rect 13068 21978 13124 21980
rect 13068 21926 13070 21978
rect 13070 21926 13122 21978
rect 13122 21926 13124 21978
rect 13068 21924 13124 21926
rect 5068 21586 5124 21588
rect 5068 21534 5070 21586
rect 5070 21534 5122 21586
rect 5122 21534 5124 21586
rect 5068 21532 5124 21534
rect 4124 21194 4180 21196
rect 4124 21142 4126 21194
rect 4126 21142 4178 21194
rect 4178 21142 4180 21194
rect 4124 21140 4180 21142
rect 4228 21194 4284 21196
rect 4228 21142 4230 21194
rect 4230 21142 4282 21194
rect 4282 21142 4284 21194
rect 4228 21140 4284 21142
rect 4332 21194 4388 21196
rect 4332 21142 4334 21194
rect 4334 21142 4386 21194
rect 4386 21142 4388 21194
rect 4332 21140 4388 21142
rect 5068 20076 5124 20132
rect 4124 19626 4180 19628
rect 4124 19574 4126 19626
rect 4126 19574 4178 19626
rect 4178 19574 4180 19626
rect 4124 19572 4180 19574
rect 4228 19626 4284 19628
rect 4228 19574 4230 19626
rect 4230 19574 4282 19626
rect 4282 19574 4284 19626
rect 4228 19572 4284 19574
rect 4332 19626 4388 19628
rect 4332 19574 4334 19626
rect 4334 19574 4386 19626
rect 4386 19574 4388 19626
rect 4332 19572 4388 19574
rect 3500 19180 3556 19236
rect 2380 17666 2436 17668
rect 2380 17614 2382 17666
rect 2382 17614 2434 17666
rect 2434 17614 2436 17666
rect 2380 17612 2436 17614
rect 2156 16268 2212 16324
rect 2828 17666 2884 17668
rect 2828 17614 2830 17666
rect 2830 17614 2882 17666
rect 2882 17614 2884 17666
rect 2828 17612 2884 17614
rect 3276 17612 3332 17668
rect 3612 18284 3668 18340
rect 3948 18450 4004 18452
rect 3948 18398 3950 18450
rect 3950 18398 4002 18450
rect 4002 18398 4004 18450
rect 3948 18396 4004 18398
rect 4396 18450 4452 18452
rect 4396 18398 4398 18450
rect 4398 18398 4450 18450
rect 4450 18398 4452 18450
rect 4396 18396 4452 18398
rect 3836 18172 3892 18228
rect 3388 17500 3444 17556
rect 2828 16322 2884 16324
rect 2828 16270 2830 16322
rect 2830 16270 2882 16322
rect 2882 16270 2884 16322
rect 2828 16268 2884 16270
rect 2716 15932 2772 15988
rect 2268 15484 2324 15540
rect 2044 15260 2100 15316
rect 2604 15314 2660 15316
rect 2604 15262 2606 15314
rect 2606 15262 2658 15314
rect 2658 15262 2660 15314
rect 2604 15260 2660 15262
rect 3164 16044 3220 16100
rect 4124 18058 4180 18060
rect 4124 18006 4126 18058
rect 4126 18006 4178 18058
rect 4178 18006 4180 18058
rect 4124 18004 4180 18006
rect 4228 18058 4284 18060
rect 4228 18006 4230 18058
rect 4230 18006 4282 18058
rect 4282 18006 4284 18058
rect 4228 18004 4284 18006
rect 4332 18058 4388 18060
rect 4332 18006 4334 18058
rect 4334 18006 4386 18058
rect 4386 18006 4388 18058
rect 4332 18004 4388 18006
rect 4124 16490 4180 16492
rect 4124 16438 4126 16490
rect 4126 16438 4178 16490
rect 4178 16438 4180 16490
rect 4124 16436 4180 16438
rect 4228 16490 4284 16492
rect 4228 16438 4230 16490
rect 4230 16438 4282 16490
rect 4282 16438 4284 16490
rect 4228 16436 4284 16438
rect 4332 16490 4388 16492
rect 4332 16438 4334 16490
rect 4334 16438 4386 16490
rect 4386 16438 4388 16490
rect 4332 16436 4388 16438
rect 3388 15708 3444 15764
rect 2828 15426 2884 15428
rect 2828 15374 2830 15426
rect 2830 15374 2882 15426
rect 2882 15374 2884 15426
rect 2828 15372 2884 15374
rect 2604 14530 2660 14532
rect 2604 14478 2606 14530
rect 2606 14478 2658 14530
rect 2658 14478 2660 14530
rect 2604 14476 2660 14478
rect 2716 14418 2772 14420
rect 2716 14366 2718 14418
rect 2718 14366 2770 14418
rect 2770 14366 2772 14418
rect 2716 14364 2772 14366
rect 3500 15372 3556 15428
rect 3276 14530 3332 14532
rect 3276 14478 3278 14530
rect 3278 14478 3330 14530
rect 3330 14478 3332 14530
rect 3276 14476 3332 14478
rect 4060 15986 4116 15988
rect 4060 15934 4062 15986
rect 4062 15934 4114 15986
rect 4114 15934 4116 15986
rect 4060 15932 4116 15934
rect 4284 15986 4340 15988
rect 4284 15934 4286 15986
rect 4286 15934 4338 15986
rect 4338 15934 4340 15986
rect 4284 15932 4340 15934
rect 4396 15708 4452 15764
rect 4124 14922 4180 14924
rect 4124 14870 4126 14922
rect 4126 14870 4178 14922
rect 4178 14870 4180 14922
rect 4124 14868 4180 14870
rect 4228 14922 4284 14924
rect 4228 14870 4230 14922
rect 4230 14870 4282 14922
rect 4282 14870 4284 14922
rect 4228 14868 4284 14870
rect 4332 14922 4388 14924
rect 4332 14870 4334 14922
rect 4334 14870 4386 14922
rect 4386 14870 4388 14922
rect 4332 14868 4388 14870
rect 4620 19346 4676 19348
rect 4620 19294 4622 19346
rect 4622 19294 4674 19346
rect 4674 19294 4676 19346
rect 4620 19292 4676 19294
rect 4844 18284 4900 18340
rect 4620 17890 4676 17892
rect 4620 17838 4622 17890
rect 4622 17838 4674 17890
rect 4674 17838 4676 17890
rect 4620 17836 4676 17838
rect 4732 17666 4788 17668
rect 4732 17614 4734 17666
rect 4734 17614 4786 17666
rect 4786 17614 4788 17666
rect 4732 17612 4788 17614
rect 4620 17554 4676 17556
rect 4620 17502 4622 17554
rect 4622 17502 4674 17554
rect 4674 17502 4676 17554
rect 4620 17500 4676 17502
rect 4844 16098 4900 16100
rect 4844 16046 4846 16098
rect 4846 16046 4898 16098
rect 4898 16046 4900 16098
rect 4844 16044 4900 16046
rect 4620 15820 4676 15876
rect 4844 15708 4900 15764
rect 7980 20802 8036 20804
rect 7980 20750 7982 20802
rect 7982 20750 8034 20802
rect 8034 20750 8036 20802
rect 7980 20748 8036 20750
rect 8428 20802 8484 20804
rect 8428 20750 8430 20802
rect 8430 20750 8482 20802
rect 8482 20750 8484 20802
rect 8428 20748 8484 20750
rect 7036 20410 7092 20412
rect 7036 20358 7038 20410
rect 7038 20358 7090 20410
rect 7090 20358 7092 20410
rect 7036 20356 7092 20358
rect 7140 20410 7196 20412
rect 7140 20358 7142 20410
rect 7142 20358 7194 20410
rect 7194 20358 7196 20410
rect 7140 20356 7196 20358
rect 7244 20410 7300 20412
rect 7244 20358 7246 20410
rect 7246 20358 7298 20410
rect 7298 20358 7300 20410
rect 7244 20356 7300 20358
rect 6972 20188 7028 20244
rect 6748 19292 6804 19348
rect 5516 18284 5572 18340
rect 5068 17836 5124 17892
rect 6300 18396 6356 18452
rect 5628 17612 5684 17668
rect 5740 17836 5796 17892
rect 5180 17052 5236 17108
rect 5292 16658 5348 16660
rect 5292 16606 5294 16658
rect 5294 16606 5346 16658
rect 5346 16606 5348 16658
rect 5292 16604 5348 16606
rect 4956 15932 5012 15988
rect 4620 15372 4676 15428
rect 5292 15820 5348 15876
rect 5964 17106 6020 17108
rect 5964 17054 5966 17106
rect 5966 17054 6018 17106
rect 6018 17054 6020 17106
rect 5964 17052 6020 17054
rect 6524 18226 6580 18228
rect 6524 18174 6526 18226
rect 6526 18174 6578 18226
rect 6578 18174 6580 18226
rect 6524 18172 6580 18174
rect 7980 20188 8036 20244
rect 9100 21532 9156 21588
rect 8092 20076 8148 20132
rect 6860 19180 6916 19236
rect 7036 18842 7092 18844
rect 7036 18790 7038 18842
rect 7038 18790 7090 18842
rect 7090 18790 7092 18842
rect 7036 18788 7092 18790
rect 7140 18842 7196 18844
rect 7140 18790 7142 18842
rect 7142 18790 7194 18842
rect 7194 18790 7196 18842
rect 7140 18788 7196 18790
rect 7244 18842 7300 18844
rect 7244 18790 7246 18842
rect 7246 18790 7298 18842
rect 7298 18790 7300 18842
rect 7244 18788 7300 18790
rect 7308 18450 7364 18452
rect 7308 18398 7310 18450
rect 7310 18398 7362 18450
rect 7362 18398 7364 18450
rect 7308 18396 7364 18398
rect 7868 19852 7924 19908
rect 7980 19234 8036 19236
rect 7980 19182 7982 19234
rect 7982 19182 8034 19234
rect 8034 19182 8036 19234
rect 7980 19180 8036 19182
rect 8876 20188 8932 20244
rect 8764 20076 8820 20132
rect 8652 20018 8708 20020
rect 8652 19966 8654 20018
rect 8654 19966 8706 20018
rect 8706 19966 8708 20018
rect 8652 19964 8708 19966
rect 8764 19794 8820 19796
rect 8764 19742 8766 19794
rect 8766 19742 8818 19794
rect 8818 19742 8820 19794
rect 8764 19740 8820 19742
rect 8316 19628 8372 19684
rect 8316 19292 8372 19348
rect 8428 19068 8484 19124
rect 7308 18172 7364 18228
rect 8204 18732 8260 18788
rect 9884 21586 9940 21588
rect 9884 21534 9886 21586
rect 9886 21534 9938 21586
rect 9938 21534 9940 21586
rect 9884 21532 9940 21534
rect 13244 21586 13300 21588
rect 13244 21534 13246 21586
rect 13246 21534 13298 21586
rect 13298 21534 13300 21586
rect 13244 21532 13300 21534
rect 9948 21194 10004 21196
rect 9948 21142 9950 21194
rect 9950 21142 10002 21194
rect 10002 21142 10004 21194
rect 9948 21140 10004 21142
rect 10052 21194 10108 21196
rect 10052 21142 10054 21194
rect 10054 21142 10106 21194
rect 10106 21142 10108 21194
rect 10052 21140 10108 21142
rect 10156 21194 10212 21196
rect 10156 21142 10158 21194
rect 10158 21142 10210 21194
rect 10210 21142 10212 21194
rect 10156 21140 10212 21142
rect 9100 19122 9156 19124
rect 9100 19070 9102 19122
rect 9102 19070 9154 19122
rect 9154 19070 9156 19122
rect 9100 19068 9156 19070
rect 8092 18562 8148 18564
rect 8092 18510 8094 18562
rect 8094 18510 8146 18562
rect 8146 18510 8148 18562
rect 8092 18508 8148 18510
rect 7756 18396 7812 18452
rect 7036 17274 7092 17276
rect 7036 17222 7038 17274
rect 7038 17222 7090 17274
rect 7090 17222 7092 17274
rect 7036 17220 7092 17222
rect 7140 17274 7196 17276
rect 7140 17222 7142 17274
rect 7142 17222 7194 17274
rect 7194 17222 7196 17274
rect 7140 17220 7196 17222
rect 7244 17274 7300 17276
rect 7244 17222 7246 17274
rect 7246 17222 7298 17274
rect 7298 17222 7300 17274
rect 7244 17220 7300 17222
rect 5628 16044 5684 16100
rect 5516 15708 5572 15764
rect 6076 16098 6132 16100
rect 6076 16046 6078 16098
rect 6078 16046 6130 16098
rect 6130 16046 6132 16098
rect 6076 16044 6132 16046
rect 6636 16604 6692 16660
rect 6076 15708 6132 15764
rect 5852 15484 5908 15540
rect 4508 14252 4564 14308
rect 5068 14140 5124 14196
rect 4396 13580 4452 13636
rect 5964 14140 6020 14196
rect 6300 15708 6356 15764
rect 6188 15372 6244 15428
rect 4620 13468 4676 13524
rect 4124 13354 4180 13356
rect 4124 13302 4126 13354
rect 4126 13302 4178 13354
rect 4178 13302 4180 13354
rect 4124 13300 4180 13302
rect 4228 13354 4284 13356
rect 4228 13302 4230 13354
rect 4230 13302 4282 13354
rect 4282 13302 4284 13354
rect 4228 13300 4284 13302
rect 4332 13354 4388 13356
rect 4332 13302 4334 13354
rect 4334 13302 4386 13354
rect 4386 13302 4388 13354
rect 4332 13300 4388 13302
rect 5404 13468 5460 13524
rect 6412 15314 6468 15316
rect 6412 15262 6414 15314
rect 6414 15262 6466 15314
rect 6466 15262 6468 15314
rect 6412 15260 6468 15262
rect 8764 18508 8820 18564
rect 8652 18396 8708 18452
rect 7756 16940 7812 16996
rect 8204 18172 8260 18228
rect 7644 16882 7700 16884
rect 7644 16830 7646 16882
rect 7646 16830 7698 16882
rect 7698 16830 7700 16882
rect 7644 16828 7700 16830
rect 8092 16882 8148 16884
rect 8092 16830 8094 16882
rect 8094 16830 8146 16882
rect 8146 16830 8148 16882
rect 8092 16828 8148 16830
rect 7420 16098 7476 16100
rect 7420 16046 7422 16098
rect 7422 16046 7474 16098
rect 7474 16046 7476 16098
rect 7420 16044 7476 16046
rect 7308 15820 7364 15876
rect 6636 15260 6692 15316
rect 6748 15708 6804 15764
rect 7036 15706 7092 15708
rect 7036 15654 7038 15706
rect 7038 15654 7090 15706
rect 7090 15654 7092 15706
rect 7036 15652 7092 15654
rect 7140 15706 7196 15708
rect 7140 15654 7142 15706
rect 7142 15654 7194 15706
rect 7194 15654 7196 15706
rect 7140 15652 7196 15654
rect 7244 15706 7300 15708
rect 7244 15654 7246 15706
rect 7246 15654 7298 15706
rect 7298 15654 7300 15706
rect 7244 15652 7300 15654
rect 6748 15372 6804 15428
rect 8652 18060 8708 18116
rect 10108 20802 10164 20804
rect 10108 20750 10110 20802
rect 10110 20750 10162 20802
rect 10162 20750 10164 20802
rect 10108 20748 10164 20750
rect 10332 20076 10388 20132
rect 9548 19740 9604 19796
rect 9884 19794 9940 19796
rect 9884 19742 9886 19794
rect 9886 19742 9938 19794
rect 9938 19742 9940 19794
rect 9884 19740 9940 19742
rect 9948 19626 10004 19628
rect 9948 19574 9950 19626
rect 9950 19574 10002 19626
rect 10002 19574 10004 19626
rect 9948 19572 10004 19574
rect 10052 19626 10108 19628
rect 10052 19574 10054 19626
rect 10054 19574 10106 19626
rect 10106 19574 10108 19626
rect 10052 19572 10108 19574
rect 10156 19626 10212 19628
rect 10156 19574 10158 19626
rect 10158 19574 10210 19626
rect 10210 19574 10212 19626
rect 10156 19572 10212 19574
rect 10780 20076 10836 20132
rect 10892 19404 10948 19460
rect 11228 19740 11284 19796
rect 9324 18732 9380 18788
rect 9884 18396 9940 18452
rect 9548 18172 9604 18228
rect 8876 17778 8932 17780
rect 8876 17726 8878 17778
rect 8878 17726 8930 17778
rect 8930 17726 8932 17778
rect 8876 17724 8932 17726
rect 9212 17724 9268 17780
rect 8540 16994 8596 16996
rect 8540 16942 8542 16994
rect 8542 16942 8594 16994
rect 8594 16942 8596 16994
rect 8540 16940 8596 16942
rect 6524 14924 6580 14980
rect 9548 16940 9604 16996
rect 9436 16882 9492 16884
rect 9436 16830 9438 16882
rect 9438 16830 9490 16882
rect 9490 16830 9492 16882
rect 9436 16828 9492 16830
rect 10444 18562 10500 18564
rect 10444 18510 10446 18562
rect 10446 18510 10498 18562
rect 10498 18510 10500 18562
rect 10444 18508 10500 18510
rect 12012 19458 12068 19460
rect 12012 19406 12014 19458
rect 12014 19406 12066 19458
rect 12066 19406 12068 19458
rect 12012 19404 12068 19406
rect 12860 20410 12916 20412
rect 12860 20358 12862 20410
rect 12862 20358 12914 20410
rect 12914 20358 12916 20410
rect 12860 20356 12916 20358
rect 12964 20410 13020 20412
rect 12964 20358 12966 20410
rect 12966 20358 13018 20410
rect 13018 20358 13020 20410
rect 12964 20356 13020 20358
rect 13068 20410 13124 20412
rect 13068 20358 13070 20410
rect 13070 20358 13122 20410
rect 13122 20358 13124 20410
rect 13068 20356 13124 20358
rect 15596 21532 15652 21588
rect 15148 21420 15204 21476
rect 12796 19404 12852 19460
rect 11900 19122 11956 19124
rect 11900 19070 11902 19122
rect 11902 19070 11954 19122
rect 11954 19070 11956 19122
rect 11900 19068 11956 19070
rect 11340 19010 11396 19012
rect 11340 18958 11342 19010
rect 11342 18958 11394 19010
rect 11394 18958 11396 19010
rect 11340 18956 11396 18958
rect 10892 18620 10948 18676
rect 11004 18732 11060 18788
rect 10780 18508 10836 18564
rect 12012 18956 12068 19012
rect 12348 19068 12404 19124
rect 11564 18674 11620 18676
rect 11564 18622 11566 18674
rect 11566 18622 11618 18674
rect 11618 18622 11620 18674
rect 11564 18620 11620 18622
rect 11228 18508 11284 18564
rect 10220 18172 10276 18228
rect 9948 18058 10004 18060
rect 9948 18006 9950 18058
rect 9950 18006 10002 18058
rect 10002 18006 10004 18058
rect 9948 18004 10004 18006
rect 10052 18058 10108 18060
rect 10052 18006 10054 18058
rect 10054 18006 10106 18058
rect 10106 18006 10108 18058
rect 10052 18004 10108 18006
rect 10156 18058 10212 18060
rect 10156 18006 10158 18058
rect 10158 18006 10210 18058
rect 10210 18006 10212 18058
rect 10156 18004 10212 18006
rect 10892 17724 10948 17780
rect 10332 16940 10388 16996
rect 9948 16490 10004 16492
rect 9948 16438 9950 16490
rect 9950 16438 10002 16490
rect 10002 16438 10004 16490
rect 9948 16436 10004 16438
rect 10052 16490 10108 16492
rect 10052 16438 10054 16490
rect 10054 16438 10106 16490
rect 10106 16438 10108 16490
rect 10052 16436 10108 16438
rect 10156 16490 10212 16492
rect 10156 16438 10158 16490
rect 10158 16438 10210 16490
rect 10210 16438 10212 16490
rect 10156 16436 10212 16438
rect 9212 16044 9268 16100
rect 8652 15426 8708 15428
rect 8652 15374 8654 15426
rect 8654 15374 8706 15426
rect 8706 15374 8708 15426
rect 8652 15372 8708 15374
rect 8092 14924 8148 14980
rect 12236 18450 12292 18452
rect 12236 18398 12238 18450
rect 12238 18398 12290 18450
rect 12290 18398 12292 18450
rect 12236 18396 12292 18398
rect 11452 17052 11508 17108
rect 12124 16940 12180 16996
rect 11564 16828 11620 16884
rect 11564 16268 11620 16324
rect 12684 19234 12740 19236
rect 12684 19182 12686 19234
rect 12686 19182 12738 19234
rect 12738 19182 12740 19234
rect 12684 19180 12740 19182
rect 12860 18842 12916 18844
rect 12860 18790 12862 18842
rect 12862 18790 12914 18842
rect 12914 18790 12916 18842
rect 12860 18788 12916 18790
rect 12964 18842 13020 18844
rect 12964 18790 12966 18842
rect 12966 18790 13018 18842
rect 13018 18790 13020 18842
rect 12964 18788 13020 18790
rect 13068 18842 13124 18844
rect 13068 18790 13070 18842
rect 13070 18790 13122 18842
rect 13122 18790 13124 18842
rect 13068 18788 13124 18790
rect 12460 18620 12516 18676
rect 13804 19122 13860 19124
rect 13804 19070 13806 19122
rect 13806 19070 13858 19122
rect 13858 19070 13860 19122
rect 13804 19068 13860 19070
rect 16044 21474 16100 21476
rect 16044 21422 16046 21474
rect 16046 21422 16098 21474
rect 16098 21422 16100 21474
rect 16044 21420 16100 21422
rect 15772 21194 15828 21196
rect 15772 21142 15774 21194
rect 15774 21142 15826 21194
rect 15826 21142 15828 21194
rect 15772 21140 15828 21142
rect 15876 21194 15932 21196
rect 15876 21142 15878 21194
rect 15878 21142 15930 21194
rect 15930 21142 15932 21194
rect 15876 21140 15932 21142
rect 15980 21194 16036 21196
rect 15980 21142 15982 21194
rect 15982 21142 16034 21194
rect 16034 21142 16036 21194
rect 15980 21140 16036 21142
rect 15596 20802 15652 20804
rect 15596 20750 15598 20802
rect 15598 20750 15650 20802
rect 15650 20750 15652 20802
rect 15596 20748 15652 20750
rect 14476 19122 14532 19124
rect 14476 19070 14478 19122
rect 14478 19070 14530 19122
rect 14530 19070 14532 19122
rect 14476 19068 14532 19070
rect 12684 18284 12740 18340
rect 14252 18956 14308 19012
rect 15036 18956 15092 19012
rect 14924 18844 14980 18900
rect 13356 18396 13412 18452
rect 12908 18172 12964 18228
rect 14812 18674 14868 18676
rect 14812 18622 14814 18674
rect 14814 18622 14866 18674
rect 14866 18622 14868 18674
rect 14812 18620 14868 18622
rect 14924 18508 14980 18564
rect 14924 18338 14980 18340
rect 14924 18286 14926 18338
rect 14926 18286 14978 18338
rect 14978 18286 14980 18338
rect 14924 18284 14980 18286
rect 13692 18172 13748 18228
rect 14364 18226 14420 18228
rect 14364 18174 14366 18226
rect 14366 18174 14418 18226
rect 14418 18174 14420 18226
rect 14364 18172 14420 18174
rect 12908 17500 12964 17556
rect 12860 17274 12916 17276
rect 12860 17222 12862 17274
rect 12862 17222 12914 17274
rect 12914 17222 12916 17274
rect 12860 17220 12916 17222
rect 12964 17274 13020 17276
rect 12964 17222 12966 17274
rect 12966 17222 13018 17274
rect 13018 17222 13020 17274
rect 12964 17220 13020 17222
rect 13068 17274 13124 17276
rect 13068 17222 13070 17274
rect 13070 17222 13122 17274
rect 13122 17222 13124 17274
rect 13068 17220 13124 17222
rect 12684 16828 12740 16884
rect 13804 16492 13860 16548
rect 12684 16268 12740 16324
rect 12236 15986 12292 15988
rect 12236 15934 12238 15986
rect 12238 15934 12290 15986
rect 12290 15934 12292 15986
rect 12236 15932 12292 15934
rect 12860 15706 12916 15708
rect 12860 15654 12862 15706
rect 12862 15654 12914 15706
rect 12914 15654 12916 15706
rect 12860 15652 12916 15654
rect 12964 15706 13020 15708
rect 12964 15654 12966 15706
rect 12966 15654 13018 15706
rect 13018 15654 13020 15706
rect 12964 15652 13020 15654
rect 13068 15706 13124 15708
rect 13068 15654 13070 15706
rect 13070 15654 13122 15706
rect 13122 15654 13124 15706
rect 13068 15652 13124 15654
rect 12012 15036 12068 15092
rect 9948 14922 10004 14924
rect 9948 14870 9950 14922
rect 9950 14870 10002 14922
rect 10002 14870 10004 14922
rect 9948 14868 10004 14870
rect 10052 14922 10108 14924
rect 10052 14870 10054 14922
rect 10054 14870 10106 14922
rect 10106 14870 10108 14922
rect 10052 14868 10108 14870
rect 10156 14922 10212 14924
rect 10156 14870 10158 14922
rect 10158 14870 10210 14922
rect 10210 14870 10212 14922
rect 10156 14868 10212 14870
rect 7036 14138 7092 14140
rect 7036 14086 7038 14138
rect 7038 14086 7090 14138
rect 7090 14086 7092 14138
rect 7036 14084 7092 14086
rect 7140 14138 7196 14140
rect 7140 14086 7142 14138
rect 7142 14086 7194 14138
rect 7194 14086 7196 14138
rect 7140 14084 7196 14086
rect 7244 14138 7300 14140
rect 7244 14086 7246 14138
rect 7246 14086 7298 14138
rect 7298 14086 7300 14138
rect 7244 14084 7300 14086
rect 4124 11786 4180 11788
rect 4124 11734 4126 11786
rect 4126 11734 4178 11786
rect 4178 11734 4180 11786
rect 4124 11732 4180 11734
rect 4228 11786 4284 11788
rect 4228 11734 4230 11786
rect 4230 11734 4282 11786
rect 4282 11734 4284 11786
rect 4228 11732 4284 11734
rect 4332 11786 4388 11788
rect 4332 11734 4334 11786
rect 4334 11734 4386 11786
rect 4386 11734 4388 11786
rect 4332 11732 4388 11734
rect 4732 11676 4788 11732
rect 3388 11564 3444 11620
rect 1820 10556 1876 10612
rect 3500 10668 3556 10724
rect 3612 8428 3668 8484
rect 4124 10218 4180 10220
rect 4124 10166 4126 10218
rect 4126 10166 4178 10218
rect 4178 10166 4180 10218
rect 4124 10164 4180 10166
rect 4228 10218 4284 10220
rect 4228 10166 4230 10218
rect 4230 10166 4282 10218
rect 4282 10166 4284 10218
rect 4228 10164 4284 10166
rect 4332 10218 4388 10220
rect 4332 10166 4334 10218
rect 4334 10166 4386 10218
rect 4386 10166 4388 10218
rect 4332 10164 4388 10166
rect 4620 10668 4676 10724
rect 4732 10610 4788 10612
rect 4732 10558 4734 10610
rect 4734 10558 4786 10610
rect 4786 10558 4788 10610
rect 4732 10556 4788 10558
rect 4620 9100 4676 9156
rect 4124 8650 4180 8652
rect 4124 8598 4126 8650
rect 4126 8598 4178 8650
rect 4178 8598 4180 8650
rect 4124 8596 4180 8598
rect 4228 8650 4284 8652
rect 4228 8598 4230 8650
rect 4230 8598 4282 8650
rect 4282 8598 4284 8650
rect 4228 8596 4284 8598
rect 4332 8650 4388 8652
rect 4332 8598 4334 8650
rect 4334 8598 4386 8650
rect 4386 8598 4388 8650
rect 4332 8596 4388 8598
rect 5516 11676 5572 11732
rect 5404 9154 5460 9156
rect 5404 9102 5406 9154
rect 5406 9102 5458 9154
rect 5458 9102 5460 9154
rect 5404 9100 5460 9102
rect 4620 8428 4676 8484
rect 7036 12570 7092 12572
rect 7036 12518 7038 12570
rect 7038 12518 7090 12570
rect 7090 12518 7092 12570
rect 7036 12516 7092 12518
rect 7140 12570 7196 12572
rect 7140 12518 7142 12570
rect 7142 12518 7194 12570
rect 7194 12518 7196 12570
rect 7140 12516 7196 12518
rect 7244 12570 7300 12572
rect 7244 12518 7246 12570
rect 7246 12518 7298 12570
rect 7298 12518 7300 12570
rect 7244 12516 7300 12518
rect 5852 11452 5908 11508
rect 6748 11506 6804 11508
rect 6748 11454 6750 11506
rect 6750 11454 6802 11506
rect 6802 11454 6804 11506
rect 6748 11452 6804 11454
rect 7036 11002 7092 11004
rect 7036 10950 7038 11002
rect 7038 10950 7090 11002
rect 7090 10950 7092 11002
rect 7036 10948 7092 10950
rect 7140 11002 7196 11004
rect 7140 10950 7142 11002
rect 7142 10950 7194 11002
rect 7194 10950 7196 11002
rect 7140 10948 7196 10950
rect 7244 11002 7300 11004
rect 7244 10950 7246 11002
rect 7246 10950 7298 11002
rect 7298 10950 7300 11002
rect 7244 10948 7300 10950
rect 5852 10556 5908 10612
rect 8092 14364 8148 14420
rect 8428 13804 8484 13860
rect 9436 13804 9492 13860
rect 9212 13692 9268 13748
rect 11340 13746 11396 13748
rect 11340 13694 11342 13746
rect 11342 13694 11394 13746
rect 11394 13694 11396 13746
rect 11340 13692 11396 13694
rect 8652 13580 8708 13636
rect 9948 13354 10004 13356
rect 9948 13302 9950 13354
rect 9950 13302 10002 13354
rect 10002 13302 10004 13354
rect 9948 13300 10004 13302
rect 10052 13354 10108 13356
rect 10052 13302 10054 13354
rect 10054 13302 10106 13354
rect 10106 13302 10108 13354
rect 10052 13300 10108 13302
rect 10156 13354 10212 13356
rect 10156 13302 10158 13354
rect 10158 13302 10210 13354
rect 10210 13302 10212 13354
rect 10156 13300 10212 13302
rect 11340 12796 11396 12852
rect 8764 12066 8820 12068
rect 8764 12014 8766 12066
rect 8766 12014 8818 12066
rect 8818 12014 8820 12066
rect 8764 12012 8820 12014
rect 7868 11452 7924 11508
rect 9100 11900 9156 11956
rect 9100 11452 9156 11508
rect 7036 9434 7092 9436
rect 7036 9382 7038 9434
rect 7038 9382 7090 9434
rect 7090 9382 7092 9434
rect 7036 9380 7092 9382
rect 7140 9434 7196 9436
rect 7140 9382 7142 9434
rect 7142 9382 7194 9434
rect 7194 9382 7196 9434
rect 7140 9380 7196 9382
rect 7244 9434 7300 9436
rect 7244 9382 7246 9434
rect 7246 9382 7298 9434
rect 7298 9382 7300 9434
rect 7244 9380 7300 9382
rect 5628 8204 5684 8260
rect 5852 8092 5908 8148
rect 4396 7980 4452 8036
rect 5740 8034 5796 8036
rect 5740 7982 5742 8034
rect 5742 7982 5794 8034
rect 5794 7982 5796 8034
rect 5740 7980 5796 7982
rect 4172 7474 4228 7476
rect 4172 7422 4174 7474
rect 4174 7422 4226 7474
rect 4226 7422 4228 7474
rect 4172 7420 4228 7422
rect 4508 7196 4564 7252
rect 4124 7082 4180 7084
rect 4124 7030 4126 7082
rect 4126 7030 4178 7082
rect 4178 7030 4180 7082
rect 4124 7028 4180 7030
rect 4228 7082 4284 7084
rect 4228 7030 4230 7082
rect 4230 7030 4282 7082
rect 4282 7030 4284 7082
rect 4228 7028 4284 7030
rect 4332 7082 4388 7084
rect 4332 7030 4334 7082
rect 4334 7030 4386 7082
rect 4386 7030 4388 7082
rect 4332 7028 4388 7030
rect 5516 7250 5572 7252
rect 5516 7198 5518 7250
rect 5518 7198 5570 7250
rect 5570 7198 5572 7250
rect 5516 7196 5572 7198
rect 9996 12236 10052 12292
rect 11340 12236 11396 12292
rect 10444 12066 10500 12068
rect 10444 12014 10446 12066
rect 10446 12014 10498 12066
rect 10498 12014 10500 12066
rect 10444 12012 10500 12014
rect 9948 11786 10004 11788
rect 9948 11734 9950 11786
rect 9950 11734 10002 11786
rect 10002 11734 10004 11786
rect 9948 11732 10004 11734
rect 10052 11786 10108 11788
rect 10052 11734 10054 11786
rect 10054 11734 10106 11786
rect 10106 11734 10108 11786
rect 10052 11732 10108 11734
rect 10156 11786 10212 11788
rect 10156 11734 10158 11786
rect 10158 11734 10210 11786
rect 10210 11734 10212 11786
rect 10156 11732 10212 11734
rect 9772 10668 9828 10724
rect 9948 10218 10004 10220
rect 9948 10166 9950 10218
rect 9950 10166 10002 10218
rect 10002 10166 10004 10218
rect 9948 10164 10004 10166
rect 10052 10218 10108 10220
rect 10052 10166 10054 10218
rect 10054 10166 10106 10218
rect 10106 10166 10108 10218
rect 10052 10164 10108 10166
rect 10156 10218 10212 10220
rect 10156 10166 10158 10218
rect 10158 10166 10210 10218
rect 10210 10166 10212 10218
rect 10156 10164 10212 10166
rect 11228 11900 11284 11956
rect 11564 11394 11620 11396
rect 11564 11342 11566 11394
rect 11566 11342 11618 11394
rect 11618 11342 11620 11394
rect 11564 11340 11620 11342
rect 11004 9884 11060 9940
rect 9996 9042 10052 9044
rect 9996 8990 9998 9042
rect 9998 8990 10050 9042
rect 10050 8990 10052 9042
rect 9996 8988 10052 8990
rect 6860 8258 6916 8260
rect 6860 8206 6862 8258
rect 6862 8206 6914 8258
rect 6914 8206 6916 8258
rect 6860 8204 6916 8206
rect 6636 8146 6692 8148
rect 6636 8094 6638 8146
rect 6638 8094 6690 8146
rect 6690 8094 6692 8146
rect 6636 8092 6692 8094
rect 6300 7980 6356 8036
rect 7036 7866 7092 7868
rect 7036 7814 7038 7866
rect 7038 7814 7090 7866
rect 7090 7814 7092 7866
rect 7036 7812 7092 7814
rect 7140 7866 7196 7868
rect 7140 7814 7142 7866
rect 7142 7814 7194 7866
rect 7194 7814 7196 7866
rect 7140 7812 7196 7814
rect 7244 7866 7300 7868
rect 7244 7814 7246 7866
rect 7246 7814 7298 7866
rect 7298 7814 7300 7866
rect 7244 7812 7300 7814
rect 6860 7644 6916 7700
rect 6524 7586 6580 7588
rect 6524 7534 6526 7586
rect 6526 7534 6578 7586
rect 6578 7534 6580 7586
rect 6524 7532 6580 7534
rect 7196 7586 7252 7588
rect 7196 7534 7198 7586
rect 7198 7534 7250 7586
rect 7250 7534 7252 7586
rect 7196 7532 7252 7534
rect 6300 7474 6356 7476
rect 6300 7422 6302 7474
rect 6302 7422 6354 7474
rect 6354 7422 6356 7474
rect 6300 7420 6356 7422
rect 8204 7644 8260 7700
rect 8316 7586 8372 7588
rect 8316 7534 8318 7586
rect 8318 7534 8370 7586
rect 8370 7534 8372 7586
rect 8316 7532 8372 7534
rect 9948 8650 10004 8652
rect 9948 8598 9950 8650
rect 9950 8598 10002 8650
rect 10002 8598 10004 8650
rect 9948 8596 10004 8598
rect 10052 8650 10108 8652
rect 10052 8598 10054 8650
rect 10054 8598 10106 8650
rect 10106 8598 10108 8650
rect 10052 8596 10108 8598
rect 10156 8650 10212 8652
rect 10156 8598 10158 8650
rect 10158 8598 10210 8650
rect 10210 8598 10212 8650
rect 10156 8596 10212 8598
rect 9436 7980 9492 8036
rect 11004 8988 11060 9044
rect 14140 15932 14196 15988
rect 13132 15314 13188 15316
rect 13132 15262 13134 15314
rect 13134 15262 13186 15314
rect 13186 15262 13188 15314
rect 13132 15260 13188 15262
rect 13356 15314 13412 15316
rect 13356 15262 13358 15314
rect 13358 15262 13410 15314
rect 13410 15262 13412 15314
rect 13356 15260 13412 15262
rect 14252 15314 14308 15316
rect 14252 15262 14254 15314
rect 14254 15262 14306 15314
rect 14306 15262 14308 15314
rect 14252 15260 14308 15262
rect 18396 22316 18452 22372
rect 21596 22762 21652 22764
rect 21596 22710 21598 22762
rect 21598 22710 21650 22762
rect 21650 22710 21652 22762
rect 21596 22708 21652 22710
rect 21700 22762 21756 22764
rect 21700 22710 21702 22762
rect 21702 22710 21754 22762
rect 21754 22710 21756 22762
rect 21700 22708 21756 22710
rect 21804 22762 21860 22764
rect 21804 22710 21806 22762
rect 21806 22710 21858 22762
rect 21858 22710 21860 22762
rect 21804 22708 21860 22710
rect 21308 22540 21364 22596
rect 22428 22594 22484 22596
rect 22428 22542 22430 22594
rect 22430 22542 22482 22594
rect 22482 22542 22484 22594
rect 22428 22540 22484 22542
rect 21420 22370 21476 22372
rect 21420 22318 21422 22370
rect 21422 22318 21474 22370
rect 21474 22318 21476 22370
rect 21420 22316 21476 22318
rect 20860 22204 20916 22260
rect 21308 22204 21364 22260
rect 20188 22146 20244 22148
rect 20188 22094 20190 22146
rect 20190 22094 20242 22146
rect 20242 22094 20244 22146
rect 20188 22092 20244 22094
rect 18684 21978 18740 21980
rect 18684 21926 18686 21978
rect 18686 21926 18738 21978
rect 18738 21926 18740 21978
rect 18684 21924 18740 21926
rect 18788 21978 18844 21980
rect 18788 21926 18790 21978
rect 18790 21926 18842 21978
rect 18842 21926 18844 21978
rect 18788 21924 18844 21926
rect 18892 21978 18948 21980
rect 18892 21926 18894 21978
rect 18894 21926 18946 21978
rect 18946 21926 18948 21978
rect 18892 21924 18948 21926
rect 21084 21868 21140 21924
rect 17836 20748 17892 20804
rect 16492 20130 16548 20132
rect 16492 20078 16494 20130
rect 16494 20078 16546 20130
rect 16546 20078 16548 20130
rect 16492 20076 16548 20078
rect 16044 19740 16100 19796
rect 15772 19626 15828 19628
rect 15772 19574 15774 19626
rect 15774 19574 15826 19626
rect 15826 19574 15828 19626
rect 15772 19572 15828 19574
rect 15876 19626 15932 19628
rect 15876 19574 15878 19626
rect 15878 19574 15930 19626
rect 15930 19574 15932 19626
rect 15876 19572 15932 19574
rect 15980 19626 16036 19628
rect 15980 19574 15982 19626
rect 15982 19574 16034 19626
rect 16034 19574 16036 19626
rect 15980 19572 16036 19574
rect 15596 19404 15652 19460
rect 15260 19234 15316 19236
rect 15260 19182 15262 19234
rect 15262 19182 15314 19234
rect 15314 19182 15316 19234
rect 15260 19180 15316 19182
rect 17724 20130 17780 20132
rect 17724 20078 17726 20130
rect 17726 20078 17778 20130
rect 17778 20078 17780 20130
rect 17724 20076 17780 20078
rect 15484 19122 15540 19124
rect 15484 19070 15486 19122
rect 15486 19070 15538 19122
rect 15538 19070 15540 19122
rect 15484 19068 15540 19070
rect 15372 18956 15428 19012
rect 15372 18226 15428 18228
rect 15372 18174 15374 18226
rect 15374 18174 15426 18226
rect 15426 18174 15428 18226
rect 15372 18172 15428 18174
rect 16156 18284 16212 18340
rect 15772 18058 15828 18060
rect 15772 18006 15774 18058
rect 15774 18006 15826 18058
rect 15826 18006 15828 18058
rect 15772 18004 15828 18006
rect 15876 18058 15932 18060
rect 15876 18006 15878 18058
rect 15878 18006 15930 18058
rect 15930 18006 15932 18058
rect 15876 18004 15932 18006
rect 15980 18058 16036 18060
rect 15980 18006 15982 18058
rect 15982 18006 16034 18058
rect 16034 18006 16036 18058
rect 15980 18004 16036 18006
rect 16156 17836 16212 17892
rect 15932 17554 15988 17556
rect 15932 17502 15934 17554
rect 15934 17502 15986 17554
rect 15986 17502 15988 17554
rect 15932 17500 15988 17502
rect 15260 17276 15316 17332
rect 14812 16492 14868 16548
rect 15772 16490 15828 16492
rect 15772 16438 15774 16490
rect 15774 16438 15826 16490
rect 15826 16438 15828 16490
rect 15772 16436 15828 16438
rect 15876 16490 15932 16492
rect 15876 16438 15878 16490
rect 15878 16438 15930 16490
rect 15930 16438 15932 16490
rect 15876 16436 15932 16438
rect 15980 16490 16036 16492
rect 15980 16438 15982 16490
rect 15982 16438 16034 16490
rect 16034 16438 16036 16490
rect 15980 16436 16036 16438
rect 16268 17500 16324 17556
rect 14700 15148 14756 15204
rect 12796 14642 12852 14644
rect 12796 14590 12798 14642
rect 12798 14590 12850 14642
rect 12850 14590 12852 14642
rect 12796 14588 12852 14590
rect 12572 14530 12628 14532
rect 12572 14478 12574 14530
rect 12574 14478 12626 14530
rect 12626 14478 12628 14530
rect 12572 14476 12628 14478
rect 13468 14530 13524 14532
rect 13468 14478 13470 14530
rect 13470 14478 13522 14530
rect 13522 14478 13524 14530
rect 13468 14476 13524 14478
rect 12860 14138 12916 14140
rect 12860 14086 12862 14138
rect 12862 14086 12914 14138
rect 12914 14086 12916 14138
rect 12860 14084 12916 14086
rect 12964 14138 13020 14140
rect 12964 14086 12966 14138
rect 12966 14086 13018 14138
rect 13018 14086 13020 14138
rect 12964 14084 13020 14086
rect 13068 14138 13124 14140
rect 13068 14086 13070 14138
rect 13070 14086 13122 14138
rect 13122 14086 13124 14138
rect 13068 14084 13124 14086
rect 14924 14588 14980 14644
rect 14252 13634 14308 13636
rect 14252 13582 14254 13634
rect 14254 13582 14306 13634
rect 14306 13582 14308 13634
rect 14252 13580 14308 13582
rect 14924 13580 14980 13636
rect 13692 13468 13748 13524
rect 14588 13522 14644 13524
rect 14588 13470 14590 13522
rect 14590 13470 14642 13522
rect 14642 13470 14644 13522
rect 14588 13468 14644 13470
rect 14028 13074 14084 13076
rect 14028 13022 14030 13074
rect 14030 13022 14082 13074
rect 14082 13022 14084 13074
rect 14028 13020 14084 13022
rect 12860 12570 12916 12572
rect 12860 12518 12862 12570
rect 12862 12518 12914 12570
rect 12914 12518 12916 12570
rect 12860 12516 12916 12518
rect 12964 12570 13020 12572
rect 12964 12518 12966 12570
rect 12966 12518 13018 12570
rect 13018 12518 13020 12570
rect 12964 12516 13020 12518
rect 13068 12570 13124 12572
rect 13068 12518 13070 12570
rect 13070 12518 13122 12570
rect 13122 12518 13124 12570
rect 13068 12516 13124 12518
rect 12572 11564 12628 11620
rect 13580 11618 13636 11620
rect 13580 11566 13582 11618
rect 13582 11566 13634 11618
rect 13634 11566 13636 11618
rect 13580 11564 13636 11566
rect 11900 11228 11956 11284
rect 12860 11002 12916 11004
rect 12860 10950 12862 11002
rect 12862 10950 12914 11002
rect 12914 10950 12916 11002
rect 12860 10948 12916 10950
rect 12964 11002 13020 11004
rect 12964 10950 12966 11002
rect 12966 10950 13018 11002
rect 13018 10950 13020 11002
rect 12964 10948 13020 10950
rect 13068 11002 13124 11004
rect 13068 10950 13070 11002
rect 13070 10950 13122 11002
rect 13122 10950 13124 11002
rect 13068 10948 13124 10950
rect 12012 9938 12068 9940
rect 12012 9886 12014 9938
rect 12014 9886 12066 9938
rect 12066 9886 12068 9938
rect 12012 9884 12068 9886
rect 12860 9434 12916 9436
rect 12860 9382 12862 9434
rect 12862 9382 12914 9434
rect 12914 9382 12916 9434
rect 12860 9380 12916 9382
rect 12964 9434 13020 9436
rect 12964 9382 12966 9434
rect 12966 9382 13018 9434
rect 13018 9382 13020 9434
rect 12964 9380 13020 9382
rect 13068 9434 13124 9436
rect 13068 9382 13070 9434
rect 13070 9382 13122 9434
rect 13122 9382 13124 9434
rect 13068 9380 13124 9382
rect 12796 8988 12852 9044
rect 11564 8258 11620 8260
rect 11564 8206 11566 8258
rect 11566 8206 11618 8258
rect 11618 8206 11620 8258
rect 11564 8204 11620 8206
rect 15708 15372 15764 15428
rect 15596 15314 15652 15316
rect 15596 15262 15598 15314
rect 15598 15262 15650 15314
rect 15650 15262 15652 15314
rect 15596 15260 15652 15262
rect 15484 15202 15540 15204
rect 15484 15150 15486 15202
rect 15486 15150 15538 15202
rect 15538 15150 15540 15202
rect 15484 15148 15540 15150
rect 15372 15036 15428 15092
rect 15772 14922 15828 14924
rect 15772 14870 15774 14922
rect 15774 14870 15826 14922
rect 15826 14870 15828 14922
rect 15772 14868 15828 14870
rect 15876 14922 15932 14924
rect 15876 14870 15878 14922
rect 15878 14870 15930 14922
rect 15930 14870 15932 14922
rect 15876 14868 15932 14870
rect 15980 14922 16036 14924
rect 15980 14870 15982 14922
rect 15982 14870 16034 14922
rect 16034 14870 16036 14922
rect 15980 14868 16036 14870
rect 16604 18844 16660 18900
rect 16492 18396 16548 18452
rect 17388 19740 17444 19796
rect 17164 19234 17220 19236
rect 17164 19182 17166 19234
rect 17166 19182 17218 19234
rect 17218 19182 17220 19234
rect 17164 19180 17220 19182
rect 16828 17554 16884 17556
rect 16828 17502 16830 17554
rect 16830 17502 16882 17554
rect 16882 17502 16884 17554
rect 16828 17500 16884 17502
rect 16940 17442 16996 17444
rect 16940 17390 16942 17442
rect 16942 17390 16994 17442
rect 16994 17390 16996 17442
rect 16940 17388 16996 17390
rect 16828 17276 16884 17332
rect 16492 15820 16548 15876
rect 18684 20410 18740 20412
rect 18684 20358 18686 20410
rect 18686 20358 18738 20410
rect 18738 20358 18740 20410
rect 18684 20356 18740 20358
rect 18788 20410 18844 20412
rect 18788 20358 18790 20410
rect 18790 20358 18842 20410
rect 18842 20358 18844 20410
rect 18788 20356 18844 20358
rect 18892 20410 18948 20412
rect 18892 20358 18894 20410
rect 18894 20358 18946 20410
rect 18946 20358 18948 20410
rect 18892 20356 18948 20358
rect 17388 18562 17444 18564
rect 17388 18510 17390 18562
rect 17390 18510 17442 18562
rect 17442 18510 17444 18562
rect 17388 18508 17444 18510
rect 17612 18844 17668 18900
rect 17500 17666 17556 17668
rect 17500 17614 17502 17666
rect 17502 17614 17554 17666
rect 17554 17614 17556 17666
rect 17500 17612 17556 17614
rect 17164 17442 17220 17444
rect 17164 17390 17166 17442
rect 17166 17390 17218 17442
rect 17218 17390 17220 17442
rect 17164 17388 17220 17390
rect 17052 16604 17108 16660
rect 17052 15484 17108 15540
rect 17164 16828 17220 16884
rect 16604 15372 16660 15428
rect 16156 13804 16212 13860
rect 15772 13354 15828 13356
rect 15772 13302 15774 13354
rect 15774 13302 15826 13354
rect 15826 13302 15828 13354
rect 15772 13300 15828 13302
rect 15876 13354 15932 13356
rect 15876 13302 15878 13354
rect 15878 13302 15930 13354
rect 15930 13302 15932 13354
rect 15876 13300 15932 13302
rect 15980 13354 16036 13356
rect 15980 13302 15982 13354
rect 15982 13302 16034 13354
rect 16034 13302 16036 13354
rect 15980 13300 16036 13302
rect 15260 13020 15316 13076
rect 14364 12348 14420 12404
rect 15596 12684 15652 12740
rect 15708 12348 15764 12404
rect 14140 12124 14196 12180
rect 15148 12178 15204 12180
rect 15148 12126 15150 12178
rect 15150 12126 15202 12178
rect 15202 12126 15204 12178
rect 15148 12124 15204 12126
rect 15484 12066 15540 12068
rect 15484 12014 15486 12066
rect 15486 12014 15538 12066
rect 15538 12014 15540 12066
rect 15484 12012 15540 12014
rect 14700 11452 14756 11508
rect 14476 11282 14532 11284
rect 14476 11230 14478 11282
rect 14478 11230 14530 11282
rect 14530 11230 14532 11282
rect 14476 11228 14532 11230
rect 16604 13020 16660 13076
rect 16492 12850 16548 12852
rect 16492 12798 16494 12850
rect 16494 12798 16546 12850
rect 16546 12798 16548 12850
rect 16492 12796 16548 12798
rect 16380 12684 16436 12740
rect 15772 11786 15828 11788
rect 15772 11734 15774 11786
rect 15774 11734 15826 11786
rect 15826 11734 15828 11786
rect 15772 11732 15828 11734
rect 15876 11786 15932 11788
rect 15876 11734 15878 11786
rect 15878 11734 15930 11786
rect 15930 11734 15932 11786
rect 15876 11732 15932 11734
rect 15980 11786 16036 11788
rect 15980 11734 15982 11786
rect 15982 11734 16034 11786
rect 16034 11734 16036 11786
rect 15980 11732 16036 11734
rect 15596 11452 15652 11508
rect 15260 10780 15316 10836
rect 14812 9212 14868 9268
rect 16492 12402 16548 12404
rect 16492 12350 16494 12402
rect 16494 12350 16546 12402
rect 16546 12350 16548 12402
rect 16492 12348 16548 12350
rect 16492 10834 16548 10836
rect 16492 10782 16494 10834
rect 16494 10782 16546 10834
rect 16546 10782 16548 10834
rect 16492 10780 16548 10782
rect 15484 8988 15540 9044
rect 13692 8204 13748 8260
rect 10444 7980 10500 8036
rect 10892 8092 10948 8148
rect 9996 7756 10052 7812
rect 8988 7420 9044 7476
rect 9100 7532 9156 7588
rect 8092 6578 8148 6580
rect 8092 6526 8094 6578
rect 8094 6526 8146 6578
rect 8146 6526 8148 6578
rect 8092 6524 8148 6526
rect 8764 6578 8820 6580
rect 8764 6526 8766 6578
rect 8766 6526 8818 6578
rect 8818 6526 8820 6578
rect 8764 6524 8820 6526
rect 7036 6298 7092 6300
rect 7036 6246 7038 6298
rect 7038 6246 7090 6298
rect 7090 6246 7092 6298
rect 7036 6244 7092 6246
rect 7140 6298 7196 6300
rect 7140 6246 7142 6298
rect 7142 6246 7194 6298
rect 7194 6246 7196 6298
rect 7140 6244 7196 6246
rect 7244 6298 7300 6300
rect 7244 6246 7246 6298
rect 7246 6246 7298 6298
rect 7298 6246 7300 6298
rect 7244 6244 7300 6246
rect 10892 7644 10948 7700
rect 10332 7474 10388 7476
rect 10332 7422 10334 7474
rect 10334 7422 10386 7474
rect 10386 7422 10388 7474
rect 10332 7420 10388 7422
rect 11116 7586 11172 7588
rect 11116 7534 11118 7586
rect 11118 7534 11170 7586
rect 11170 7534 11172 7586
rect 11116 7532 11172 7534
rect 9948 7082 10004 7084
rect 9948 7030 9950 7082
rect 9950 7030 10002 7082
rect 10002 7030 10004 7082
rect 9948 7028 10004 7030
rect 10052 7082 10108 7084
rect 10052 7030 10054 7082
rect 10054 7030 10106 7082
rect 10106 7030 10108 7082
rect 10052 7028 10108 7030
rect 10156 7082 10212 7084
rect 10156 7030 10158 7082
rect 10158 7030 10210 7082
rect 10210 7030 10212 7082
rect 10156 7028 10212 7030
rect 13468 8146 13524 8148
rect 13468 8094 13470 8146
rect 13470 8094 13522 8146
rect 13522 8094 13524 8146
rect 13468 8092 13524 8094
rect 12012 7532 12068 7588
rect 12860 7866 12916 7868
rect 12860 7814 12862 7866
rect 12862 7814 12914 7866
rect 12914 7814 12916 7866
rect 12860 7812 12916 7814
rect 12964 7866 13020 7868
rect 12964 7814 12966 7866
rect 12966 7814 13018 7866
rect 13018 7814 13020 7866
rect 12964 7812 13020 7814
rect 13068 7866 13124 7868
rect 13068 7814 13070 7866
rect 13070 7814 13122 7866
rect 13122 7814 13124 7866
rect 13068 7812 13124 7814
rect 12796 7532 12852 7588
rect 15772 10218 15828 10220
rect 15772 10166 15774 10218
rect 15774 10166 15826 10218
rect 15826 10166 15828 10218
rect 15772 10164 15828 10166
rect 15876 10218 15932 10220
rect 15876 10166 15878 10218
rect 15878 10166 15930 10218
rect 15930 10166 15932 10218
rect 15876 10164 15932 10166
rect 15980 10218 16036 10220
rect 15980 10166 15982 10218
rect 15982 10166 16034 10218
rect 16034 10166 16036 10218
rect 15980 10164 16036 10166
rect 17724 17836 17780 17892
rect 19292 19852 19348 19908
rect 19740 20802 19796 20804
rect 19740 20750 19742 20802
rect 19742 20750 19794 20802
rect 19794 20750 19796 20802
rect 19740 20748 19796 20750
rect 20748 20748 20804 20804
rect 20748 20188 20804 20244
rect 19292 19180 19348 19236
rect 18684 18842 18740 18844
rect 18684 18790 18686 18842
rect 18686 18790 18738 18842
rect 18738 18790 18740 18842
rect 18684 18788 18740 18790
rect 18788 18842 18844 18844
rect 18788 18790 18790 18842
rect 18790 18790 18842 18842
rect 18842 18790 18844 18842
rect 18788 18788 18844 18790
rect 18892 18842 18948 18844
rect 18892 18790 18894 18842
rect 18894 18790 18946 18842
rect 18946 18790 18948 18842
rect 18892 18788 18948 18790
rect 20076 19852 20132 19908
rect 20300 19404 20356 19460
rect 19740 18562 19796 18564
rect 19740 18510 19742 18562
rect 19742 18510 19794 18562
rect 19794 18510 19796 18562
rect 19740 18508 19796 18510
rect 18060 18450 18116 18452
rect 18060 18398 18062 18450
rect 18062 18398 18114 18450
rect 18114 18398 18116 18450
rect 18060 18396 18116 18398
rect 18396 18284 18452 18340
rect 19516 18450 19572 18452
rect 19516 18398 19518 18450
rect 19518 18398 19570 18450
rect 19570 18398 19572 18450
rect 19516 18396 19572 18398
rect 17836 17612 17892 17668
rect 17612 15484 17668 15540
rect 20076 18338 20132 18340
rect 20076 18286 20078 18338
rect 20078 18286 20130 18338
rect 20130 18286 20132 18338
rect 20076 18284 20132 18286
rect 23660 22092 23716 22148
rect 23548 21868 23604 21924
rect 21596 21194 21652 21196
rect 21596 21142 21598 21194
rect 21598 21142 21650 21194
rect 21650 21142 21652 21194
rect 21596 21140 21652 21142
rect 21700 21194 21756 21196
rect 21700 21142 21702 21194
rect 21702 21142 21754 21194
rect 21754 21142 21756 21194
rect 21700 21140 21756 21142
rect 21804 21194 21860 21196
rect 21804 21142 21806 21194
rect 21806 21142 21858 21194
rect 21858 21142 21860 21194
rect 21804 21140 21860 21142
rect 22540 20860 22596 20916
rect 21980 20188 22036 20244
rect 21196 18508 21252 18564
rect 20412 17836 20468 17892
rect 20636 18172 20692 18228
rect 19068 17388 19124 17444
rect 18684 17274 18740 17276
rect 18684 17222 18686 17274
rect 18686 17222 18738 17274
rect 18738 17222 18740 17274
rect 18684 17220 18740 17222
rect 18788 17274 18844 17276
rect 18788 17222 18790 17274
rect 18790 17222 18842 17274
rect 18842 17222 18844 17274
rect 18788 17220 18844 17222
rect 18892 17274 18948 17276
rect 18892 17222 18894 17274
rect 18894 17222 18946 17274
rect 18946 17222 18948 17274
rect 18892 17220 18948 17222
rect 18284 15874 18340 15876
rect 18284 15822 18286 15874
rect 18286 15822 18338 15874
rect 18338 15822 18340 15874
rect 18284 15820 18340 15822
rect 18684 15706 18740 15708
rect 18172 15484 18228 15540
rect 18508 15596 18564 15652
rect 18684 15654 18686 15706
rect 18686 15654 18738 15706
rect 18738 15654 18740 15706
rect 18684 15652 18740 15654
rect 18788 15706 18844 15708
rect 18788 15654 18790 15706
rect 18790 15654 18842 15706
rect 18842 15654 18844 15706
rect 18788 15652 18844 15654
rect 18892 15706 18948 15708
rect 18892 15654 18894 15706
rect 18894 15654 18946 15706
rect 18946 15654 18948 15706
rect 18892 15652 18948 15654
rect 18844 15426 18900 15428
rect 18844 15374 18846 15426
rect 18846 15374 18898 15426
rect 18898 15374 18900 15426
rect 18844 15372 18900 15374
rect 17500 13746 17556 13748
rect 17500 13694 17502 13746
rect 17502 13694 17554 13746
rect 17554 13694 17556 13746
rect 17500 13692 17556 13694
rect 18172 14476 18228 14532
rect 18172 14252 18228 14308
rect 19068 14306 19124 14308
rect 19068 14254 19070 14306
rect 19070 14254 19122 14306
rect 19122 14254 19124 14306
rect 19068 14252 19124 14254
rect 18684 14138 18740 14140
rect 18684 14086 18686 14138
rect 18686 14086 18738 14138
rect 18738 14086 18740 14138
rect 18684 14084 18740 14086
rect 18788 14138 18844 14140
rect 18788 14086 18790 14138
rect 18790 14086 18842 14138
rect 18842 14086 18844 14138
rect 18788 14084 18844 14086
rect 18892 14138 18948 14140
rect 18892 14086 18894 14138
rect 18894 14086 18946 14138
rect 18946 14086 18948 14138
rect 18892 14084 18948 14086
rect 17724 13468 17780 13524
rect 18396 13468 18452 13524
rect 17388 12796 17444 12852
rect 19516 15484 19572 15540
rect 19852 15314 19908 15316
rect 19852 15262 19854 15314
rect 19854 15262 19906 15314
rect 19906 15262 19908 15314
rect 19852 15260 19908 15262
rect 20972 17612 21028 17668
rect 20636 17164 20692 17220
rect 20524 15932 20580 15988
rect 20524 15260 20580 15316
rect 20076 15036 20132 15092
rect 20188 14588 20244 14644
rect 19292 14530 19348 14532
rect 19292 14478 19294 14530
rect 19294 14478 19346 14530
rect 19346 14478 19348 14530
rect 19292 14476 19348 14478
rect 20748 16156 20804 16212
rect 20860 15036 20916 15092
rect 20636 13746 20692 13748
rect 20636 13694 20638 13746
rect 20638 13694 20690 13746
rect 20690 13694 20692 13746
rect 20636 13692 20692 13694
rect 19404 13580 19460 13636
rect 18956 12850 19012 12852
rect 18956 12798 18958 12850
rect 18958 12798 19010 12850
rect 19010 12798 19012 12850
rect 18956 12796 19012 12798
rect 18684 12570 18740 12572
rect 18684 12518 18686 12570
rect 18686 12518 18738 12570
rect 18738 12518 18740 12570
rect 18684 12516 18740 12518
rect 18788 12570 18844 12572
rect 18788 12518 18790 12570
rect 18790 12518 18842 12570
rect 18842 12518 18844 12570
rect 18788 12516 18844 12518
rect 18892 12570 18948 12572
rect 18892 12518 18894 12570
rect 18894 12518 18946 12570
rect 18946 12518 18948 12570
rect 18892 12516 18948 12518
rect 18956 12236 19012 12292
rect 17500 12066 17556 12068
rect 17500 12014 17502 12066
rect 17502 12014 17554 12066
rect 17554 12014 17556 12066
rect 17500 12012 17556 12014
rect 16940 11394 16996 11396
rect 16940 11342 16942 11394
rect 16942 11342 16994 11394
rect 16994 11342 16996 11394
rect 16940 11340 16996 11342
rect 18684 11002 18740 11004
rect 18684 10950 18686 11002
rect 18686 10950 18738 11002
rect 18738 10950 18740 11002
rect 18684 10948 18740 10950
rect 18788 11002 18844 11004
rect 18788 10950 18790 11002
rect 18790 10950 18842 11002
rect 18842 10950 18844 11002
rect 18788 10948 18844 10950
rect 18892 11002 18948 11004
rect 18892 10950 18894 11002
rect 18894 10950 18946 11002
rect 18946 10950 18948 11002
rect 18892 10948 18948 10950
rect 17388 10108 17444 10164
rect 16604 9266 16660 9268
rect 16604 9214 16606 9266
rect 16606 9214 16658 9266
rect 16658 9214 16660 9266
rect 16604 9212 16660 9214
rect 16044 9042 16100 9044
rect 16044 8990 16046 9042
rect 16046 8990 16098 9042
rect 16098 8990 16100 9042
rect 16044 8988 16100 8990
rect 15708 8764 15764 8820
rect 15772 8650 15828 8652
rect 15772 8598 15774 8650
rect 15774 8598 15826 8650
rect 15826 8598 15828 8650
rect 15772 8596 15828 8598
rect 15876 8650 15932 8652
rect 15876 8598 15878 8650
rect 15878 8598 15930 8650
rect 15930 8598 15932 8650
rect 15876 8596 15932 8598
rect 15980 8650 16036 8652
rect 15980 8598 15982 8650
rect 15982 8598 16034 8650
rect 16034 8598 16036 8650
rect 15980 8596 16036 8598
rect 15484 7532 15540 7588
rect 11452 7308 11508 7364
rect 13916 7362 13972 7364
rect 13916 7310 13918 7362
rect 13918 7310 13970 7362
rect 13970 7310 13972 7362
rect 13916 7308 13972 7310
rect 18284 9996 18340 10052
rect 19292 11676 19348 11732
rect 19740 12290 19796 12292
rect 19740 12238 19742 12290
rect 19742 12238 19794 12290
rect 19794 12238 19796 12290
rect 19740 12236 19796 12238
rect 19964 12684 20020 12740
rect 19516 11452 19572 11508
rect 19068 9996 19124 10052
rect 20300 13020 20356 13076
rect 20076 12178 20132 12180
rect 20076 12126 20078 12178
rect 20078 12126 20130 12178
rect 20130 12126 20132 12178
rect 20076 12124 20132 12126
rect 19964 11340 20020 11396
rect 20524 10780 20580 10836
rect 20636 12236 20692 12292
rect 16492 7308 16548 7364
rect 16828 8764 16884 8820
rect 17388 8764 17444 8820
rect 21868 19964 21924 20020
rect 23212 20690 23268 20692
rect 23212 20638 23214 20690
rect 23214 20638 23266 20690
rect 23266 20638 23268 20690
rect 23212 20636 23268 20638
rect 23212 20188 23268 20244
rect 21596 19626 21652 19628
rect 21596 19574 21598 19626
rect 21598 19574 21650 19626
rect 21650 19574 21652 19626
rect 21596 19572 21652 19574
rect 21700 19626 21756 19628
rect 21700 19574 21702 19626
rect 21702 19574 21754 19626
rect 21754 19574 21756 19626
rect 21700 19572 21756 19574
rect 21804 19626 21860 19628
rect 21804 19574 21806 19626
rect 21806 19574 21858 19626
rect 21858 19574 21860 19626
rect 21804 19572 21860 19574
rect 24508 21978 24564 21980
rect 24508 21926 24510 21978
rect 24510 21926 24562 21978
rect 24562 21926 24564 21978
rect 24508 21924 24564 21926
rect 24612 21978 24668 21980
rect 24612 21926 24614 21978
rect 24614 21926 24666 21978
rect 24666 21926 24668 21978
rect 24612 21924 24668 21926
rect 24716 21978 24772 21980
rect 24716 21926 24718 21978
rect 24718 21926 24770 21978
rect 24770 21926 24772 21978
rect 24716 21924 24772 21926
rect 23996 20914 24052 20916
rect 23996 20862 23998 20914
rect 23998 20862 24050 20914
rect 24050 20862 24052 20914
rect 23996 20860 24052 20862
rect 24508 20410 24564 20412
rect 24508 20358 24510 20410
rect 24510 20358 24562 20410
rect 24562 20358 24564 20410
rect 24508 20356 24564 20358
rect 24612 20410 24668 20412
rect 24612 20358 24614 20410
rect 24614 20358 24666 20410
rect 24666 20358 24668 20410
rect 24612 20356 24668 20358
rect 24716 20410 24772 20412
rect 24716 20358 24718 20410
rect 24718 20358 24770 20410
rect 24770 20358 24772 20410
rect 24716 20356 24772 20358
rect 22876 19906 22932 19908
rect 22876 19854 22878 19906
rect 22878 19854 22930 19906
rect 22930 19854 22932 19906
rect 22876 19852 22932 19854
rect 22204 19404 22260 19460
rect 21596 18058 21652 18060
rect 21596 18006 21598 18058
rect 21598 18006 21650 18058
rect 21650 18006 21652 18058
rect 21596 18004 21652 18006
rect 21700 18058 21756 18060
rect 21700 18006 21702 18058
rect 21702 18006 21754 18058
rect 21754 18006 21756 18058
rect 21700 18004 21756 18006
rect 21804 18058 21860 18060
rect 21804 18006 21806 18058
rect 21806 18006 21858 18058
rect 21858 18006 21860 18058
rect 21804 18004 21860 18006
rect 21308 17890 21364 17892
rect 21308 17838 21310 17890
rect 21310 17838 21362 17890
rect 21362 17838 21364 17890
rect 21308 17836 21364 17838
rect 22092 18172 22148 18228
rect 22316 18396 22372 18452
rect 22652 17890 22708 17892
rect 22652 17838 22654 17890
rect 22654 17838 22706 17890
rect 22706 17838 22708 17890
rect 22652 17836 22708 17838
rect 21868 17164 21924 17220
rect 21980 16828 22036 16884
rect 21308 15932 21364 15988
rect 21420 16604 21476 16660
rect 21596 16490 21652 16492
rect 21596 16438 21598 16490
rect 21598 16438 21650 16490
rect 21650 16438 21652 16490
rect 21596 16436 21652 16438
rect 21700 16490 21756 16492
rect 21700 16438 21702 16490
rect 21702 16438 21754 16490
rect 21754 16438 21756 16490
rect 21700 16436 21756 16438
rect 21804 16490 21860 16492
rect 21804 16438 21806 16490
rect 21806 16438 21858 16490
rect 21858 16438 21860 16490
rect 21804 16436 21860 16438
rect 21868 16098 21924 16100
rect 21868 16046 21870 16098
rect 21870 16046 21922 16098
rect 21922 16046 21924 16098
rect 21868 16044 21924 16046
rect 21644 15148 21700 15204
rect 21532 15036 21588 15092
rect 21596 14922 21652 14924
rect 21596 14870 21598 14922
rect 21598 14870 21650 14922
rect 21650 14870 21652 14922
rect 21596 14868 21652 14870
rect 21700 14922 21756 14924
rect 21700 14870 21702 14922
rect 21702 14870 21754 14922
rect 21754 14870 21756 14922
rect 21700 14868 21756 14870
rect 21804 14922 21860 14924
rect 21804 14870 21806 14922
rect 21806 14870 21858 14922
rect 21858 14870 21860 14922
rect 21804 14868 21860 14870
rect 21532 14306 21588 14308
rect 21532 14254 21534 14306
rect 21534 14254 21586 14306
rect 21586 14254 21588 14306
rect 21532 14252 21588 14254
rect 23212 17164 23268 17220
rect 23884 17164 23940 17220
rect 22428 16156 22484 16212
rect 23100 16882 23156 16884
rect 23100 16830 23102 16882
rect 23102 16830 23154 16882
rect 23154 16830 23156 16882
rect 23100 16828 23156 16830
rect 22876 16604 22932 16660
rect 22092 15372 22148 15428
rect 22988 15426 23044 15428
rect 22988 15374 22990 15426
rect 22990 15374 23042 15426
rect 23042 15374 23044 15426
rect 22988 15372 23044 15374
rect 22428 15036 22484 15092
rect 21420 13634 21476 13636
rect 21420 13582 21422 13634
rect 21422 13582 21474 13634
rect 21474 13582 21476 13634
rect 21420 13580 21476 13582
rect 21596 13354 21652 13356
rect 21596 13302 21598 13354
rect 21598 13302 21650 13354
rect 21650 13302 21652 13354
rect 21596 13300 21652 13302
rect 21700 13354 21756 13356
rect 21700 13302 21702 13354
rect 21702 13302 21754 13354
rect 21754 13302 21756 13354
rect 21700 13300 21756 13302
rect 21804 13354 21860 13356
rect 21804 13302 21806 13354
rect 21806 13302 21858 13354
rect 21858 13302 21860 13354
rect 21804 13300 21860 13302
rect 21644 12738 21700 12740
rect 21644 12686 21646 12738
rect 21646 12686 21698 12738
rect 21698 12686 21700 12738
rect 21644 12684 21700 12686
rect 21420 12236 21476 12292
rect 21644 12290 21700 12292
rect 21644 12238 21646 12290
rect 21646 12238 21698 12290
rect 21698 12238 21700 12290
rect 21644 12236 21700 12238
rect 21308 11506 21364 11508
rect 21308 11454 21310 11506
rect 21310 11454 21362 11506
rect 21362 11454 21364 11506
rect 21308 11452 21364 11454
rect 22092 13020 22148 13076
rect 22652 14642 22708 14644
rect 22652 14590 22654 14642
rect 22654 14590 22706 14642
rect 22706 14590 22708 14642
rect 22652 14588 22708 14590
rect 23100 14364 23156 14420
rect 23100 13804 23156 13860
rect 23100 12684 23156 12740
rect 21868 11900 21924 11956
rect 22204 12348 22260 12404
rect 21596 11786 21652 11788
rect 21596 11734 21598 11786
rect 21598 11734 21650 11786
rect 21650 11734 21652 11786
rect 21596 11732 21652 11734
rect 21700 11786 21756 11788
rect 21700 11734 21702 11786
rect 21702 11734 21754 11786
rect 21754 11734 21756 11786
rect 21700 11732 21756 11734
rect 21804 11786 21860 11788
rect 21804 11734 21806 11786
rect 21806 11734 21858 11786
rect 21858 11734 21860 11786
rect 21804 11732 21860 11734
rect 22540 12236 22596 12292
rect 22092 11900 22148 11956
rect 20748 10556 20804 10612
rect 21756 10556 21812 10612
rect 18684 9434 18740 9436
rect 18684 9382 18686 9434
rect 18686 9382 18738 9434
rect 18738 9382 18740 9434
rect 18684 9380 18740 9382
rect 18788 9434 18844 9436
rect 18788 9382 18790 9434
rect 18790 9382 18842 9434
rect 18842 9382 18844 9434
rect 18788 9380 18844 9382
rect 18892 9434 18948 9436
rect 18892 9382 18894 9434
rect 18894 9382 18946 9434
rect 18946 9382 18948 9434
rect 20860 9436 20916 9492
rect 18892 9380 18948 9382
rect 19740 8988 19796 9044
rect 18508 8428 18564 8484
rect 19628 8428 19684 8484
rect 15772 7082 15828 7084
rect 15772 7030 15774 7082
rect 15774 7030 15826 7082
rect 15826 7030 15828 7082
rect 15772 7028 15828 7030
rect 15876 7082 15932 7084
rect 15876 7030 15878 7082
rect 15878 7030 15930 7082
rect 15930 7030 15932 7082
rect 15876 7028 15932 7030
rect 15980 7082 16036 7084
rect 15980 7030 15982 7082
rect 15982 7030 16034 7082
rect 16034 7030 16036 7082
rect 15980 7028 16036 7030
rect 18284 8034 18340 8036
rect 18284 7982 18286 8034
rect 18286 7982 18338 8034
rect 18338 7982 18340 8034
rect 18284 7980 18340 7982
rect 18684 7866 18740 7868
rect 18684 7814 18686 7866
rect 18686 7814 18738 7866
rect 18738 7814 18740 7866
rect 18684 7812 18740 7814
rect 18788 7866 18844 7868
rect 18788 7814 18790 7866
rect 18790 7814 18842 7866
rect 18842 7814 18844 7866
rect 18788 7812 18844 7814
rect 18892 7866 18948 7868
rect 18892 7814 18894 7866
rect 18894 7814 18946 7866
rect 18946 7814 18948 7866
rect 19516 7868 19572 7924
rect 18892 7812 18948 7814
rect 20300 8988 20356 9044
rect 22092 10780 22148 10836
rect 21868 10332 21924 10388
rect 21596 10218 21652 10220
rect 21308 10108 21364 10164
rect 21596 10166 21598 10218
rect 21598 10166 21650 10218
rect 21650 10166 21652 10218
rect 21596 10164 21652 10166
rect 21700 10218 21756 10220
rect 21700 10166 21702 10218
rect 21702 10166 21754 10218
rect 21754 10166 21756 10218
rect 21700 10164 21756 10166
rect 21804 10218 21860 10220
rect 21804 10166 21806 10218
rect 21806 10166 21858 10218
rect 21858 10166 21860 10218
rect 21804 10164 21860 10166
rect 21980 10108 22036 10164
rect 21644 9436 21700 9492
rect 21084 9042 21140 9044
rect 21084 8990 21086 9042
rect 21086 8990 21138 9042
rect 21138 8990 21140 9042
rect 21084 8988 21140 8990
rect 21420 8540 21476 8596
rect 21596 8650 21652 8652
rect 21596 8598 21598 8650
rect 21598 8598 21650 8650
rect 21650 8598 21652 8650
rect 21596 8596 21652 8598
rect 21700 8650 21756 8652
rect 21700 8598 21702 8650
rect 21702 8598 21754 8650
rect 21754 8598 21756 8650
rect 21700 8596 21756 8598
rect 21804 8650 21860 8652
rect 21804 8598 21806 8650
rect 21806 8598 21858 8650
rect 21858 8598 21860 8650
rect 21804 8596 21860 8598
rect 20972 8316 21028 8372
rect 20076 8092 20132 8148
rect 18956 7474 19012 7476
rect 18956 7422 18958 7474
rect 18958 7422 19010 7474
rect 19010 7422 19012 7474
rect 18956 7420 19012 7422
rect 20412 8034 20468 8036
rect 20412 7982 20414 8034
rect 20414 7982 20466 8034
rect 20466 7982 20468 8034
rect 20412 7980 20468 7982
rect 20524 7868 20580 7924
rect 20748 7756 20804 7812
rect 20076 7420 20132 7476
rect 20524 7420 20580 7476
rect 16828 6636 16884 6692
rect 12012 6466 12068 6468
rect 12012 6414 12014 6466
rect 12014 6414 12066 6466
rect 12066 6414 12068 6466
rect 12012 6412 12068 6414
rect 13468 6412 13524 6468
rect 12860 6298 12916 6300
rect 12860 6246 12862 6298
rect 12862 6246 12914 6298
rect 12914 6246 12916 6298
rect 12860 6244 12916 6246
rect 12964 6298 13020 6300
rect 12964 6246 12966 6298
rect 12966 6246 13018 6298
rect 13018 6246 13020 6298
rect 12964 6244 13020 6246
rect 13068 6298 13124 6300
rect 13068 6246 13070 6298
rect 13070 6246 13122 6298
rect 13122 6246 13124 6298
rect 13068 6244 13124 6246
rect 14252 5906 14308 5908
rect 14252 5854 14254 5906
rect 14254 5854 14306 5906
rect 14306 5854 14308 5906
rect 14252 5852 14308 5854
rect 17724 6690 17780 6692
rect 17724 6638 17726 6690
rect 17726 6638 17778 6690
rect 17778 6638 17780 6690
rect 17724 6636 17780 6638
rect 18684 6298 18740 6300
rect 18684 6246 18686 6298
rect 18686 6246 18738 6298
rect 18738 6246 18740 6298
rect 18684 6244 18740 6246
rect 18788 6298 18844 6300
rect 18788 6246 18790 6298
rect 18790 6246 18842 6298
rect 18842 6246 18844 6298
rect 18788 6244 18844 6246
rect 18892 6298 18948 6300
rect 18892 6246 18894 6298
rect 18894 6246 18946 6298
rect 18946 6246 18948 6298
rect 18892 6244 18948 6246
rect 22764 11394 22820 11396
rect 22764 11342 22766 11394
rect 22766 11342 22818 11394
rect 22818 11342 22820 11394
rect 22764 11340 22820 11342
rect 22316 10556 22372 10612
rect 22540 10780 22596 10836
rect 21644 8428 21700 8484
rect 21084 8092 21140 8148
rect 20972 7420 21028 7476
rect 21308 7980 21364 8036
rect 21532 8146 21588 8148
rect 21532 8094 21534 8146
rect 21534 8094 21586 8146
rect 21586 8094 21588 8146
rect 21532 8092 21588 8094
rect 21420 7868 21476 7924
rect 21644 7756 21700 7812
rect 21420 7474 21476 7476
rect 21420 7422 21422 7474
rect 21422 7422 21474 7474
rect 21474 7422 21476 7474
rect 21420 7420 21476 7422
rect 22092 8370 22148 8372
rect 22092 8318 22094 8370
rect 22094 8318 22146 8370
rect 22146 8318 22148 8370
rect 22092 8316 22148 8318
rect 22652 7644 22708 7700
rect 21596 7082 21652 7084
rect 21596 7030 21598 7082
rect 21598 7030 21650 7082
rect 21650 7030 21652 7082
rect 21596 7028 21652 7030
rect 21700 7082 21756 7084
rect 21700 7030 21702 7082
rect 21702 7030 21754 7082
rect 21754 7030 21756 7082
rect 21700 7028 21756 7030
rect 21804 7082 21860 7084
rect 21804 7030 21806 7082
rect 21806 7030 21858 7082
rect 21858 7030 21860 7082
rect 21804 7028 21860 7030
rect 16828 5852 16884 5908
rect 21308 6690 21364 6692
rect 21308 6638 21310 6690
rect 21310 6638 21362 6690
rect 21362 6638 21364 6690
rect 21308 6636 21364 6638
rect 4124 5514 4180 5516
rect 4124 5462 4126 5514
rect 4126 5462 4178 5514
rect 4178 5462 4180 5514
rect 4124 5460 4180 5462
rect 4228 5514 4284 5516
rect 4228 5462 4230 5514
rect 4230 5462 4282 5514
rect 4282 5462 4284 5514
rect 4228 5460 4284 5462
rect 4332 5514 4388 5516
rect 4332 5462 4334 5514
rect 4334 5462 4386 5514
rect 4386 5462 4388 5514
rect 4332 5460 4388 5462
rect 9948 5514 10004 5516
rect 9948 5462 9950 5514
rect 9950 5462 10002 5514
rect 10002 5462 10004 5514
rect 9948 5460 10004 5462
rect 10052 5514 10108 5516
rect 10052 5462 10054 5514
rect 10054 5462 10106 5514
rect 10106 5462 10108 5514
rect 10052 5460 10108 5462
rect 10156 5514 10212 5516
rect 10156 5462 10158 5514
rect 10158 5462 10210 5514
rect 10210 5462 10212 5514
rect 10156 5460 10212 5462
rect 15772 5514 15828 5516
rect 15772 5462 15774 5514
rect 15774 5462 15826 5514
rect 15826 5462 15828 5514
rect 15772 5460 15828 5462
rect 15876 5514 15932 5516
rect 15876 5462 15878 5514
rect 15878 5462 15930 5514
rect 15930 5462 15932 5514
rect 15876 5460 15932 5462
rect 15980 5514 16036 5516
rect 15980 5462 15982 5514
rect 15982 5462 16034 5514
rect 16034 5462 16036 5514
rect 15980 5460 16036 5462
rect 23324 16044 23380 16100
rect 23996 16268 24052 16324
rect 24220 19852 24276 19908
rect 24508 18842 24564 18844
rect 24508 18790 24510 18842
rect 24510 18790 24562 18842
rect 24562 18790 24564 18842
rect 24508 18788 24564 18790
rect 24612 18842 24668 18844
rect 24612 18790 24614 18842
rect 24614 18790 24666 18842
rect 24666 18790 24668 18842
rect 24612 18788 24668 18790
rect 24716 18842 24772 18844
rect 24716 18790 24718 18842
rect 24718 18790 24770 18842
rect 24770 18790 24772 18842
rect 24716 18788 24772 18790
rect 24220 17948 24276 18004
rect 24508 17274 24564 17276
rect 24508 17222 24510 17274
rect 24510 17222 24562 17274
rect 24562 17222 24564 17274
rect 24508 17220 24564 17222
rect 24612 17274 24668 17276
rect 24612 17222 24614 17274
rect 24614 17222 24666 17274
rect 24666 17222 24668 17274
rect 24612 17220 24668 17222
rect 24716 17274 24772 17276
rect 24716 17222 24718 17274
rect 24718 17222 24770 17274
rect 24770 17222 24772 17274
rect 24716 17220 24772 17222
rect 23548 15820 23604 15876
rect 23324 14588 23380 14644
rect 24332 15932 24388 15988
rect 23884 14418 23940 14420
rect 23884 14366 23886 14418
rect 23886 14366 23938 14418
rect 23938 14366 23940 14418
rect 23884 14364 23940 14366
rect 23884 13858 23940 13860
rect 23884 13806 23886 13858
rect 23886 13806 23938 13858
rect 23938 13806 23940 13858
rect 23884 13804 23940 13806
rect 23324 13074 23380 13076
rect 23324 13022 23326 13074
rect 23326 13022 23378 13074
rect 23378 13022 23380 13074
rect 23324 13020 23380 13022
rect 23884 12738 23940 12740
rect 23884 12686 23886 12738
rect 23886 12686 23938 12738
rect 23938 12686 23940 12738
rect 23884 12684 23940 12686
rect 23548 12124 23604 12180
rect 23324 9042 23380 9044
rect 23324 8990 23326 9042
rect 23326 8990 23378 9042
rect 23378 8990 23380 9042
rect 23324 8988 23380 8990
rect 22876 8034 22932 8036
rect 22876 7982 22878 8034
rect 22878 7982 22930 8034
rect 22930 7982 22932 8034
rect 22876 7980 22932 7982
rect 23324 7980 23380 8036
rect 22876 7420 22932 7476
rect 22988 5964 23044 6020
rect 23324 5852 23380 5908
rect 21596 5514 21652 5516
rect 21596 5462 21598 5514
rect 21598 5462 21650 5514
rect 21650 5462 21652 5514
rect 21596 5460 21652 5462
rect 21700 5514 21756 5516
rect 21700 5462 21702 5514
rect 21702 5462 21754 5514
rect 21754 5462 21756 5514
rect 21700 5460 21756 5462
rect 21804 5514 21860 5516
rect 21804 5462 21806 5514
rect 21806 5462 21858 5514
rect 21858 5462 21860 5514
rect 21804 5460 21860 5462
rect 20972 5180 21028 5236
rect 23548 5234 23604 5236
rect 23548 5182 23550 5234
rect 23550 5182 23602 5234
rect 23602 5182 23604 5234
rect 23548 5180 23604 5182
rect 23884 9436 23940 9492
rect 24508 15706 24564 15708
rect 24508 15654 24510 15706
rect 24510 15654 24562 15706
rect 24562 15654 24564 15706
rect 24508 15652 24564 15654
rect 24612 15706 24668 15708
rect 24612 15654 24614 15706
rect 24614 15654 24666 15706
rect 24666 15654 24668 15706
rect 24612 15652 24668 15654
rect 24716 15706 24772 15708
rect 24716 15654 24718 15706
rect 24718 15654 24770 15706
rect 24770 15654 24772 15706
rect 24716 15652 24772 15654
rect 24220 14252 24276 14308
rect 24508 14138 24564 14140
rect 24508 14086 24510 14138
rect 24510 14086 24562 14138
rect 24562 14086 24564 14138
rect 24508 14084 24564 14086
rect 24612 14138 24668 14140
rect 24612 14086 24614 14138
rect 24614 14086 24666 14138
rect 24666 14086 24668 14138
rect 24612 14084 24668 14086
rect 24716 14138 24772 14140
rect 24716 14086 24718 14138
rect 24718 14086 24770 14138
rect 24770 14086 24772 14138
rect 24716 14084 24772 14086
rect 24220 13916 24276 13972
rect 24220 12850 24276 12852
rect 24220 12798 24222 12850
rect 24222 12798 24274 12850
rect 24274 12798 24276 12850
rect 24220 12796 24276 12798
rect 24220 11900 24276 11956
rect 24508 12570 24564 12572
rect 24508 12518 24510 12570
rect 24510 12518 24562 12570
rect 24562 12518 24564 12570
rect 24508 12516 24564 12518
rect 24612 12570 24668 12572
rect 24612 12518 24614 12570
rect 24614 12518 24666 12570
rect 24666 12518 24668 12570
rect 24612 12516 24668 12518
rect 24716 12570 24772 12572
rect 24716 12518 24718 12570
rect 24718 12518 24770 12570
rect 24770 12518 24772 12570
rect 24716 12516 24772 12518
rect 24508 11002 24564 11004
rect 24508 10950 24510 11002
rect 24510 10950 24562 11002
rect 24562 10950 24564 11002
rect 24508 10948 24564 10950
rect 24612 11002 24668 11004
rect 24612 10950 24614 11002
rect 24614 10950 24666 11002
rect 24666 10950 24668 11002
rect 24612 10948 24668 10950
rect 24716 11002 24772 11004
rect 24716 10950 24718 11002
rect 24718 10950 24770 11002
rect 24770 10950 24772 11002
rect 24716 10948 24772 10950
rect 24220 9436 24276 9492
rect 24332 9884 24388 9940
rect 24108 7756 24164 7812
rect 24508 9434 24564 9436
rect 24508 9382 24510 9434
rect 24510 9382 24562 9434
rect 24562 9382 24564 9434
rect 24508 9380 24564 9382
rect 24612 9434 24668 9436
rect 24612 9382 24614 9434
rect 24614 9382 24666 9434
rect 24666 9382 24668 9434
rect 24612 9380 24668 9382
rect 24716 9434 24772 9436
rect 24716 9382 24718 9434
rect 24718 9382 24770 9434
rect 24770 9382 24772 9434
rect 24716 9380 24772 9382
rect 24508 7866 24564 7868
rect 24508 7814 24510 7866
rect 24510 7814 24562 7866
rect 24562 7814 24564 7866
rect 24508 7812 24564 7814
rect 24612 7866 24668 7868
rect 24612 7814 24614 7866
rect 24614 7814 24666 7866
rect 24666 7814 24668 7866
rect 24612 7812 24668 7814
rect 24716 7866 24772 7868
rect 24716 7814 24718 7866
rect 24718 7814 24770 7866
rect 24770 7814 24772 7866
rect 24716 7812 24772 7814
rect 24220 7420 24276 7476
rect 24508 6298 24564 6300
rect 24508 6246 24510 6298
rect 24510 6246 24562 6298
rect 24562 6246 24564 6298
rect 24508 6244 24564 6246
rect 24612 6298 24668 6300
rect 24612 6246 24614 6298
rect 24614 6246 24666 6298
rect 24666 6246 24668 6298
rect 24612 6244 24668 6246
rect 24716 6298 24772 6300
rect 24716 6246 24718 6298
rect 24718 6246 24770 6298
rect 24770 6246 24772 6298
rect 24716 6244 24772 6246
rect 7036 4730 7092 4732
rect 7036 4678 7038 4730
rect 7038 4678 7090 4730
rect 7090 4678 7092 4730
rect 7036 4676 7092 4678
rect 7140 4730 7196 4732
rect 7140 4678 7142 4730
rect 7142 4678 7194 4730
rect 7194 4678 7196 4730
rect 7140 4676 7196 4678
rect 7244 4730 7300 4732
rect 7244 4678 7246 4730
rect 7246 4678 7298 4730
rect 7298 4678 7300 4730
rect 7244 4676 7300 4678
rect 12860 4730 12916 4732
rect 12860 4678 12862 4730
rect 12862 4678 12914 4730
rect 12914 4678 12916 4730
rect 12860 4676 12916 4678
rect 12964 4730 13020 4732
rect 12964 4678 12966 4730
rect 12966 4678 13018 4730
rect 13018 4678 13020 4730
rect 12964 4676 13020 4678
rect 13068 4730 13124 4732
rect 13068 4678 13070 4730
rect 13070 4678 13122 4730
rect 13122 4678 13124 4730
rect 13068 4676 13124 4678
rect 18684 4730 18740 4732
rect 18684 4678 18686 4730
rect 18686 4678 18738 4730
rect 18738 4678 18740 4730
rect 18684 4676 18740 4678
rect 18788 4730 18844 4732
rect 18788 4678 18790 4730
rect 18790 4678 18842 4730
rect 18842 4678 18844 4730
rect 18788 4676 18844 4678
rect 18892 4730 18948 4732
rect 18892 4678 18894 4730
rect 18894 4678 18946 4730
rect 18946 4678 18948 4730
rect 18892 4676 18948 4678
rect 4124 3946 4180 3948
rect 4124 3894 4126 3946
rect 4126 3894 4178 3946
rect 4178 3894 4180 3946
rect 4124 3892 4180 3894
rect 4228 3946 4284 3948
rect 4228 3894 4230 3946
rect 4230 3894 4282 3946
rect 4282 3894 4284 3946
rect 4228 3892 4284 3894
rect 4332 3946 4388 3948
rect 4332 3894 4334 3946
rect 4334 3894 4386 3946
rect 4386 3894 4388 3946
rect 4332 3892 4388 3894
rect 9948 3946 10004 3948
rect 9948 3894 9950 3946
rect 9950 3894 10002 3946
rect 10002 3894 10004 3946
rect 9948 3892 10004 3894
rect 10052 3946 10108 3948
rect 10052 3894 10054 3946
rect 10054 3894 10106 3946
rect 10106 3894 10108 3946
rect 10052 3892 10108 3894
rect 10156 3946 10212 3948
rect 10156 3894 10158 3946
rect 10158 3894 10210 3946
rect 10210 3894 10212 3946
rect 10156 3892 10212 3894
rect 15772 3946 15828 3948
rect 15772 3894 15774 3946
rect 15774 3894 15826 3946
rect 15826 3894 15828 3946
rect 15772 3892 15828 3894
rect 15876 3946 15932 3948
rect 15876 3894 15878 3946
rect 15878 3894 15930 3946
rect 15930 3894 15932 3946
rect 15876 3892 15932 3894
rect 15980 3946 16036 3948
rect 15980 3894 15982 3946
rect 15982 3894 16034 3946
rect 16034 3894 16036 3946
rect 15980 3892 16036 3894
rect 21596 3946 21652 3948
rect 21596 3894 21598 3946
rect 21598 3894 21650 3946
rect 21650 3894 21652 3946
rect 21596 3892 21652 3894
rect 21700 3946 21756 3948
rect 21700 3894 21702 3946
rect 21702 3894 21754 3946
rect 21754 3894 21756 3946
rect 21700 3892 21756 3894
rect 21804 3946 21860 3948
rect 21804 3894 21806 3946
rect 21806 3894 21858 3946
rect 21858 3894 21860 3946
rect 21804 3892 21860 3894
rect 23436 3442 23492 3444
rect 23436 3390 23438 3442
rect 23438 3390 23490 3442
rect 23490 3390 23492 3442
rect 23436 3388 23492 3390
rect 24508 4730 24564 4732
rect 24508 4678 24510 4730
rect 24510 4678 24562 4730
rect 24562 4678 24564 4730
rect 24508 4676 24564 4678
rect 24612 4730 24668 4732
rect 24612 4678 24614 4730
rect 24614 4678 24666 4730
rect 24666 4678 24668 4730
rect 24612 4676 24668 4678
rect 24716 4730 24772 4732
rect 24716 4678 24718 4730
rect 24718 4678 24770 4730
rect 24770 4678 24772 4730
rect 24716 4676 24772 4678
rect 24220 3836 24276 3892
rect 23884 3388 23940 3444
rect 7036 3162 7092 3164
rect 7036 3110 7038 3162
rect 7038 3110 7090 3162
rect 7090 3110 7092 3162
rect 7036 3108 7092 3110
rect 7140 3162 7196 3164
rect 7140 3110 7142 3162
rect 7142 3110 7194 3162
rect 7194 3110 7196 3162
rect 7140 3108 7196 3110
rect 7244 3162 7300 3164
rect 7244 3110 7246 3162
rect 7246 3110 7298 3162
rect 7298 3110 7300 3162
rect 7244 3108 7300 3110
rect 12860 3162 12916 3164
rect 12860 3110 12862 3162
rect 12862 3110 12914 3162
rect 12914 3110 12916 3162
rect 12860 3108 12916 3110
rect 12964 3162 13020 3164
rect 12964 3110 12966 3162
rect 12966 3110 13018 3162
rect 13018 3110 13020 3162
rect 12964 3108 13020 3110
rect 13068 3162 13124 3164
rect 13068 3110 13070 3162
rect 13070 3110 13122 3162
rect 13122 3110 13124 3162
rect 13068 3108 13124 3110
rect 18684 3162 18740 3164
rect 18684 3110 18686 3162
rect 18686 3110 18738 3162
rect 18738 3110 18740 3162
rect 18684 3108 18740 3110
rect 18788 3162 18844 3164
rect 18788 3110 18790 3162
rect 18790 3110 18842 3162
rect 18842 3110 18844 3162
rect 18788 3108 18844 3110
rect 18892 3162 18948 3164
rect 18892 3110 18894 3162
rect 18894 3110 18946 3162
rect 18946 3110 18948 3162
rect 18892 3108 18948 3110
rect 24508 3162 24564 3164
rect 24508 3110 24510 3162
rect 24510 3110 24562 3162
rect 24562 3110 24564 3162
rect 24508 3108 24564 3110
rect 24612 3162 24668 3164
rect 24612 3110 24614 3162
rect 24614 3110 24666 3162
rect 24666 3110 24668 3162
rect 24612 3108 24668 3110
rect 24716 3162 24772 3164
rect 24716 3110 24718 3162
rect 24718 3110 24770 3162
rect 24770 3110 24772 3162
rect 24716 3108 24772 3110
rect 23996 1820 24052 1876
<< metal3 >>
rect 25200 24052 26000 24080
rect 20290 23996 20300 24052
rect 20356 23996 26000 24052
rect 25200 23968 26000 23996
rect 4114 22708 4124 22764
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4388 22708 4398 22764
rect 9938 22708 9948 22764
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 10212 22708 10222 22764
rect 15762 22708 15772 22764
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 16036 22708 16046 22764
rect 21586 22708 21596 22764
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21860 22708 21870 22764
rect 21298 22540 21308 22596
rect 21364 22540 22428 22596
rect 22484 22540 22494 22596
rect 17490 22316 17500 22372
rect 17556 22316 18396 22372
rect 18452 22316 21420 22372
rect 21476 22316 21486 22372
rect 20850 22204 20860 22260
rect 20916 22204 21308 22260
rect 21364 22204 24948 22260
rect 20178 22092 20188 22148
rect 20244 22092 23660 22148
rect 23716 22092 23726 22148
rect 24892 22036 24948 22204
rect 25200 22036 26000 22064
rect 24892 21980 26000 22036
rect 7026 21924 7036 21980
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7300 21924 7310 21980
rect 12850 21924 12860 21980
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 13124 21924 13134 21980
rect 18674 21924 18684 21980
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18948 21924 18958 21980
rect 24498 21924 24508 21980
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24772 21924 24782 21980
rect 25200 21952 26000 21980
rect 21074 21868 21084 21924
rect 21140 21868 23548 21924
rect 23604 21868 23614 21924
rect 5058 21532 5068 21588
rect 5124 21532 9100 21588
rect 9156 21532 9884 21588
rect 9940 21532 9950 21588
rect 13234 21532 13244 21588
rect 13300 21532 15596 21588
rect 15652 21532 15662 21588
rect 15138 21420 15148 21476
rect 15204 21420 16044 21476
rect 16100 21420 16110 21476
rect 4114 21140 4124 21196
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4388 21140 4398 21196
rect 9938 21140 9948 21196
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 10212 21140 10222 21196
rect 15762 21140 15772 21196
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 16036 21140 16046 21196
rect 21586 21140 21596 21196
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21860 21140 21870 21196
rect 22530 20860 22540 20916
rect 22596 20860 23996 20916
rect 24052 20860 24062 20916
rect 7970 20748 7980 20804
rect 8036 20748 8428 20804
rect 8484 20748 10108 20804
rect 10164 20748 10174 20804
rect 15586 20748 15596 20804
rect 15652 20748 17836 20804
rect 17892 20748 17902 20804
rect 19730 20748 19740 20804
rect 19796 20748 20748 20804
rect 20804 20748 20814 20804
rect 23174 20636 23212 20692
rect 23268 20636 23278 20692
rect 7026 20356 7036 20412
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7300 20356 7310 20412
rect 12850 20356 12860 20412
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 13124 20356 13134 20412
rect 18674 20356 18684 20412
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18948 20356 18958 20412
rect 24498 20356 24508 20412
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24772 20356 24782 20412
rect 6962 20188 6972 20244
rect 7028 20188 7980 20244
rect 8036 20188 8876 20244
rect 8932 20188 8942 20244
rect 20738 20188 20748 20244
rect 20804 20188 21980 20244
rect 22036 20188 23212 20244
rect 23268 20188 23278 20244
rect 3490 20076 3500 20132
rect 3556 20076 5068 20132
rect 5124 20076 5134 20132
rect 8082 20076 8092 20132
rect 8148 20076 8764 20132
rect 8820 20076 10332 20132
rect 10388 20076 10780 20132
rect 10836 20076 10846 20132
rect 16482 20076 16492 20132
rect 16548 20076 17724 20132
rect 17780 20076 17790 20132
rect 25200 20020 26000 20048
rect 8642 19964 8652 20020
rect 8708 19964 8718 20020
rect 21858 19964 21868 20020
rect 21924 19964 26000 20020
rect 8652 19908 8708 19964
rect 25200 19936 26000 19964
rect 7858 19852 7868 19908
rect 7924 19852 8708 19908
rect 19282 19852 19292 19908
rect 19348 19852 20076 19908
rect 20132 19852 20142 19908
rect 22866 19852 22876 19908
rect 22932 19852 24220 19908
rect 24276 19852 24286 19908
rect 8316 19684 8372 19852
rect 8754 19740 8764 19796
rect 8820 19740 9548 19796
rect 9604 19740 9614 19796
rect 9874 19740 9884 19796
rect 9940 19740 11228 19796
rect 11284 19740 11294 19796
rect 16034 19740 16044 19796
rect 16100 19740 17388 19796
rect 17444 19740 17454 19796
rect 8306 19628 8316 19684
rect 8372 19628 8382 19684
rect 4114 19572 4124 19628
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4388 19572 4398 19628
rect 9938 19572 9948 19628
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 10212 19572 10222 19628
rect 15762 19572 15772 19628
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 16036 19572 16046 19628
rect 21586 19572 21596 19628
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21860 19572 21870 19628
rect 10882 19404 10892 19460
rect 10948 19404 12012 19460
rect 12068 19404 12078 19460
rect 12786 19404 12796 19460
rect 12852 19404 15596 19460
rect 15652 19404 15662 19460
rect 20290 19404 20300 19460
rect 20356 19404 22204 19460
rect 22260 19404 22270 19460
rect 4610 19292 4620 19348
rect 4676 19292 6748 19348
rect 6804 19292 8316 19348
rect 8372 19292 8382 19348
rect 1810 19180 1820 19236
rect 1876 19180 3500 19236
rect 3556 19180 3566 19236
rect 6850 19180 6860 19236
rect 6916 19180 7980 19236
rect 8036 19180 8046 19236
rect 12674 19180 12684 19236
rect 12740 19180 15260 19236
rect 15316 19180 15326 19236
rect 17154 19180 17164 19236
rect 17220 19180 19292 19236
rect 19348 19180 19358 19236
rect 8418 19068 8428 19124
rect 8484 19068 9100 19124
rect 9156 19068 9166 19124
rect 11890 19068 11900 19124
rect 11956 19068 12348 19124
rect 12404 19068 13300 19124
rect 13794 19068 13804 19124
rect 13860 19068 14476 19124
rect 14532 19068 15484 19124
rect 15540 19068 15550 19124
rect 11330 18956 11340 19012
rect 11396 18956 12012 19012
rect 12068 18956 12078 19012
rect 7026 18788 7036 18844
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7300 18788 7310 18844
rect 12850 18788 12860 18844
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 13124 18788 13134 18844
rect 13244 18788 13300 19068
rect 14242 18956 14252 19012
rect 14308 18956 15036 19012
rect 15092 18956 15372 19012
rect 15428 18956 15438 19012
rect 14914 18844 14924 18900
rect 14980 18844 16604 18900
rect 16660 18844 17612 18900
rect 17668 18844 17678 18900
rect 18674 18788 18684 18844
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18948 18788 18958 18844
rect 24498 18788 24508 18844
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24772 18788 24782 18844
rect 8194 18732 8204 18788
rect 8260 18732 9324 18788
rect 9380 18732 11004 18788
rect 11060 18732 11070 18788
rect 13244 18732 15148 18788
rect 10882 18620 10892 18676
rect 10948 18620 11564 18676
rect 11620 18620 11630 18676
rect 12450 18620 12460 18676
rect 12516 18620 14812 18676
rect 14868 18620 14878 18676
rect 15092 18564 15148 18732
rect 8082 18508 8092 18564
rect 8148 18508 8764 18564
rect 8820 18508 10444 18564
rect 10500 18508 10510 18564
rect 10770 18508 10780 18564
rect 10836 18508 11228 18564
rect 11284 18508 11294 18564
rect 14588 18508 14924 18564
rect 14980 18508 14990 18564
rect 15092 18508 17388 18564
rect 17444 18508 17454 18564
rect 19730 18508 19740 18564
rect 19796 18508 21196 18564
rect 21252 18508 21262 18564
rect 3938 18396 3948 18452
rect 4004 18396 4396 18452
rect 4452 18396 6300 18452
rect 6356 18396 6366 18452
rect 7298 18396 7308 18452
rect 7364 18396 7756 18452
rect 7812 18396 7822 18452
rect 8642 18396 8652 18452
rect 8708 18396 9884 18452
rect 9940 18396 9950 18452
rect 12226 18396 12236 18452
rect 12292 18396 13356 18452
rect 13412 18396 13422 18452
rect 14588 18340 14644 18508
rect 16482 18396 16492 18452
rect 16548 18396 18060 18452
rect 18116 18396 18126 18452
rect 19506 18396 19516 18452
rect 19572 18396 22316 18452
rect 22372 18396 22382 18452
rect 3602 18284 3612 18340
rect 3668 18284 4844 18340
rect 4900 18284 5012 18340
rect 5506 18284 5516 18340
rect 5572 18284 12684 18340
rect 12740 18284 14644 18340
rect 14914 18284 14924 18340
rect 14980 18284 16156 18340
rect 16212 18284 16222 18340
rect 18386 18284 18396 18340
rect 18452 18284 20076 18340
rect 20132 18284 20142 18340
rect 3836 18228 3892 18284
rect 4956 18228 5012 18284
rect 3826 18172 3836 18228
rect 3892 18172 3902 18228
rect 4956 18172 6020 18228
rect 6514 18172 6524 18228
rect 6580 18172 7308 18228
rect 7364 18172 8204 18228
rect 8260 18172 8270 18228
rect 9538 18172 9548 18228
rect 9604 18172 10220 18228
rect 10276 18172 10286 18228
rect 12898 18172 12908 18228
rect 12964 18172 13692 18228
rect 13748 18172 13758 18228
rect 14354 18172 14364 18228
rect 14420 18172 15372 18228
rect 15428 18172 15438 18228
rect 20626 18172 20636 18228
rect 20692 18172 22092 18228
rect 22148 18172 22158 18228
rect 5964 18116 6020 18172
rect 5964 18060 8652 18116
rect 8708 18060 8718 18116
rect 4114 18004 4124 18060
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4388 18004 4398 18060
rect 9938 18004 9948 18060
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 10212 18004 10222 18060
rect 15762 18004 15772 18060
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 16036 18004 16046 18060
rect 21586 18004 21596 18060
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21860 18004 21870 18060
rect 25200 18004 26000 18032
rect 24210 17948 24220 18004
rect 24276 17948 26000 18004
rect 25200 17920 26000 17948
rect 4610 17836 4620 17892
rect 4676 17836 5068 17892
rect 5124 17836 5740 17892
rect 5796 17836 5806 17892
rect 16146 17836 16156 17892
rect 16212 17836 17724 17892
rect 17780 17836 17790 17892
rect 20402 17836 20412 17892
rect 20468 17836 21308 17892
rect 21364 17836 22652 17892
rect 22708 17836 22718 17892
rect 8866 17724 8876 17780
rect 8932 17724 9212 17780
rect 9268 17724 10892 17780
rect 10948 17724 10958 17780
rect 2370 17612 2380 17668
rect 2436 17612 2828 17668
rect 2884 17612 3276 17668
rect 3332 17612 3342 17668
rect 4722 17612 4732 17668
rect 4788 17612 5628 17668
rect 5684 17612 5694 17668
rect 17490 17612 17500 17668
rect 17556 17612 17836 17668
rect 17892 17612 20972 17668
rect 21028 17612 21038 17668
rect 3378 17500 3388 17556
rect 3444 17500 4620 17556
rect 4676 17500 12908 17556
rect 12964 17500 15148 17556
rect 15922 17500 15932 17556
rect 15988 17500 16268 17556
rect 16324 17500 16828 17556
rect 16884 17500 16894 17556
rect 15092 17444 15148 17500
rect 15092 17388 16940 17444
rect 16996 17388 17006 17444
rect 17154 17388 17164 17444
rect 17220 17388 19068 17444
rect 19124 17388 19134 17444
rect 15250 17276 15260 17332
rect 15316 17276 16828 17332
rect 16884 17276 16894 17332
rect 7026 17220 7036 17276
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7300 17220 7310 17276
rect 12850 17220 12860 17276
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 13124 17220 13134 17276
rect 18674 17220 18684 17276
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18948 17220 18958 17276
rect 24498 17220 24508 17276
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24772 17220 24782 17276
rect 20626 17164 20636 17220
rect 20692 17164 21868 17220
rect 21924 17164 23212 17220
rect 23268 17164 23884 17220
rect 23940 17164 23950 17220
rect 5170 17052 5180 17108
rect 5236 17052 5964 17108
rect 6020 17052 11452 17108
rect 11508 17052 11518 17108
rect 7746 16940 7756 16996
rect 7812 16940 8540 16996
rect 8596 16940 9548 16996
rect 9604 16940 9940 16996
rect 10322 16940 10332 16996
rect 10388 16940 12124 16996
rect 12180 16940 12190 16996
rect 9884 16884 9940 16940
rect 7634 16828 7644 16884
rect 7700 16828 8092 16884
rect 8148 16828 9436 16884
rect 9492 16828 9502 16884
rect 9884 16828 11564 16884
rect 11620 16828 11630 16884
rect 12674 16828 12684 16884
rect 12740 16828 17164 16884
rect 17220 16828 17230 16884
rect 21970 16828 21980 16884
rect 22036 16828 23100 16884
rect 23156 16828 23166 16884
rect 5282 16604 5292 16660
rect 5348 16604 6636 16660
rect 6692 16604 6702 16660
rect 15092 16604 17052 16660
rect 17108 16604 17118 16660
rect 21410 16604 21420 16660
rect 21476 16604 22876 16660
rect 22932 16604 22942 16660
rect 15092 16548 15148 16604
rect 13794 16492 13804 16548
rect 13860 16492 14812 16548
rect 14868 16492 15148 16548
rect 4114 16436 4124 16492
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4388 16436 4398 16492
rect 9938 16436 9948 16492
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 10212 16436 10222 16492
rect 15762 16436 15772 16492
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 16036 16436 16046 16492
rect 21586 16436 21596 16492
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21860 16436 21870 16492
rect 2146 16268 2156 16324
rect 2212 16268 2828 16324
rect 2884 16268 2894 16324
rect 11554 16268 11564 16324
rect 11620 16268 12684 16324
rect 12740 16268 23996 16324
rect 24052 16268 24062 16324
rect 20738 16156 20748 16212
rect 20804 16156 22428 16212
rect 22484 16156 22494 16212
rect 3154 16044 3164 16100
rect 3220 16044 4844 16100
rect 4900 16044 5628 16100
rect 5684 16044 6076 16100
rect 6132 16044 6142 16100
rect 7410 16044 7420 16100
rect 7476 16044 9212 16100
rect 9268 16044 9278 16100
rect 21858 16044 21868 16100
rect 21924 16044 23324 16100
rect 23380 16044 23390 16100
rect 25200 15988 26000 16016
rect 2706 15932 2716 15988
rect 2772 15932 4060 15988
rect 4116 15932 4126 15988
rect 4274 15932 4284 15988
rect 4340 15932 4956 15988
rect 5012 15932 5022 15988
rect 12226 15932 12236 15988
rect 12292 15932 14140 15988
rect 14196 15932 14206 15988
rect 20514 15932 20524 15988
rect 20580 15932 21308 15988
rect 21364 15932 21374 15988
rect 24322 15932 24332 15988
rect 24388 15932 26000 15988
rect 4284 15876 4340 15932
rect 25200 15904 26000 15932
rect 3388 15820 4340 15876
rect 4610 15820 4620 15876
rect 4676 15820 5292 15876
rect 5348 15820 7308 15876
rect 7364 15820 7374 15876
rect 16482 15820 16492 15876
rect 16548 15820 18284 15876
rect 18340 15820 23548 15876
rect 23604 15820 23614 15876
rect 3388 15764 3444 15820
rect 3378 15708 3388 15764
rect 3444 15708 3454 15764
rect 4386 15708 4396 15764
rect 4452 15708 4844 15764
rect 4900 15708 4910 15764
rect 5506 15708 5516 15764
rect 5572 15708 6076 15764
rect 6132 15708 6300 15764
rect 6356 15708 6748 15764
rect 6804 15708 6814 15764
rect 7026 15652 7036 15708
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7300 15652 7310 15708
rect 12850 15652 12860 15708
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 13124 15652 13134 15708
rect 18674 15652 18684 15708
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18948 15652 18958 15708
rect 24498 15652 24508 15708
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24772 15652 24782 15708
rect 17612 15596 18508 15652
rect 18564 15596 18574 15652
rect 17612 15540 17668 15596
rect 2258 15484 2268 15540
rect 2324 15484 5852 15540
rect 5908 15484 5918 15540
rect 17042 15484 17052 15540
rect 17108 15484 17612 15540
rect 17668 15484 17678 15540
rect 18162 15484 18172 15540
rect 18228 15484 19516 15540
rect 19572 15484 19582 15540
rect 2818 15372 2828 15428
rect 2884 15372 3500 15428
rect 3556 15372 4620 15428
rect 4676 15372 4686 15428
rect 5404 15372 6188 15428
rect 6244 15372 6254 15428
rect 6738 15372 6748 15428
rect 6804 15372 8652 15428
rect 8708 15372 8718 15428
rect 15698 15372 15708 15428
rect 15764 15372 16604 15428
rect 16660 15372 18844 15428
rect 18900 15372 22092 15428
rect 22148 15372 22158 15428
rect 22950 15372 22988 15428
rect 23044 15372 23054 15428
rect 5404 15316 5460 15372
rect 2034 15260 2044 15316
rect 2100 15260 2604 15316
rect 2660 15260 5460 15316
rect 6402 15260 6412 15316
rect 6468 15260 6636 15316
rect 6692 15260 6702 15316
rect 13122 15260 13132 15316
rect 13188 15260 13198 15316
rect 13346 15260 13356 15316
rect 13412 15260 14252 15316
rect 14308 15260 15596 15316
rect 15652 15260 15662 15316
rect 19842 15260 19852 15316
rect 19908 15260 20524 15316
rect 20580 15260 20590 15316
rect 13132 15092 13188 15260
rect 14690 15148 14700 15204
rect 14756 15148 15484 15204
rect 15540 15148 15550 15204
rect 21308 15148 21644 15204
rect 21700 15148 21710 15204
rect 21308 15092 21364 15148
rect 12002 15036 12012 15092
rect 12068 15036 15372 15092
rect 15428 15036 15438 15092
rect 20066 15036 20076 15092
rect 20132 15036 20860 15092
rect 20916 15036 21364 15092
rect 21522 15036 21532 15092
rect 21588 15036 22428 15092
rect 22484 15036 22494 15092
rect 6514 14924 6524 14980
rect 6580 14924 8092 14980
rect 8148 14924 8158 14980
rect 4114 14868 4124 14924
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4388 14868 4398 14924
rect 9938 14868 9948 14924
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 10212 14868 10222 14924
rect 15762 14868 15772 14924
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 16036 14868 16046 14924
rect 21586 14868 21596 14924
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21860 14868 21870 14924
rect 12786 14588 12796 14644
rect 12852 14588 14924 14644
rect 14980 14588 14990 14644
rect 20178 14588 20188 14644
rect 20244 14588 22652 14644
rect 22708 14588 23324 14644
rect 23380 14588 23390 14644
rect 2594 14476 2604 14532
rect 2660 14476 3276 14532
rect 3332 14476 3342 14532
rect 8372 14476 12572 14532
rect 12628 14476 13468 14532
rect 13524 14476 13534 14532
rect 18162 14476 18172 14532
rect 18228 14476 19292 14532
rect 19348 14476 19358 14532
rect 2706 14364 2716 14420
rect 2772 14364 8092 14420
rect 8148 14364 8158 14420
rect 8372 14308 8428 14476
rect 23090 14364 23100 14420
rect 23156 14364 23884 14420
rect 23940 14364 23950 14420
rect 4498 14252 4508 14308
rect 4564 14252 8428 14308
rect 18162 14252 18172 14308
rect 18228 14252 19068 14308
rect 19124 14252 19134 14308
rect 21522 14252 21532 14308
rect 21588 14252 24220 14308
rect 24276 14252 24286 14308
rect 5058 14140 5068 14196
rect 5124 14140 5964 14196
rect 6020 14140 6030 14196
rect 7026 14084 7036 14140
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7300 14084 7310 14140
rect 12850 14084 12860 14140
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 13124 14084 13134 14140
rect 18674 14084 18684 14140
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18948 14084 18958 14140
rect 24498 14084 24508 14140
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24772 14084 24782 14140
rect 25200 13972 26000 14000
rect 24210 13916 24220 13972
rect 24276 13916 26000 13972
rect 25200 13888 26000 13916
rect 8418 13804 8428 13860
rect 8484 13804 9436 13860
rect 9492 13804 9502 13860
rect 15092 13804 16156 13860
rect 16212 13804 16222 13860
rect 23090 13804 23100 13860
rect 23156 13804 23884 13860
rect 23940 13804 23950 13860
rect 9202 13692 9212 13748
rect 9268 13692 11340 13748
rect 11396 13692 11406 13748
rect 4386 13580 4396 13636
rect 4452 13580 8652 13636
rect 8708 13580 8718 13636
rect 14242 13580 14252 13636
rect 14308 13580 14924 13636
rect 14980 13580 14990 13636
rect 15092 13524 15148 13804
rect 17490 13692 17500 13748
rect 17556 13692 20636 13748
rect 20692 13692 20702 13748
rect 19394 13580 19404 13636
rect 19460 13580 21420 13636
rect 21476 13580 21486 13636
rect 4610 13468 4620 13524
rect 4676 13468 5404 13524
rect 5460 13468 5470 13524
rect 13682 13468 13692 13524
rect 13748 13468 14588 13524
rect 14644 13468 15148 13524
rect 17714 13468 17724 13524
rect 17780 13468 18396 13524
rect 18452 13468 18462 13524
rect 4114 13300 4124 13356
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4388 13300 4398 13356
rect 9938 13300 9948 13356
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 10212 13300 10222 13356
rect 15762 13300 15772 13356
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 16036 13300 16046 13356
rect 21586 13300 21596 13356
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21860 13300 21870 13356
rect 14018 13020 14028 13076
rect 14084 13020 15260 13076
rect 15316 13020 16604 13076
rect 16660 13020 16670 13076
rect 20290 13020 20300 13076
rect 20356 13020 22092 13076
rect 22148 13020 23324 13076
rect 23380 13020 23390 13076
rect 14028 12852 14084 13020
rect 11330 12796 11340 12852
rect 11396 12796 14084 12852
rect 16482 12796 16492 12852
rect 16548 12796 17388 12852
rect 17444 12796 17454 12852
rect 18946 12796 18956 12852
rect 19012 12796 24220 12852
rect 24276 12796 24286 12852
rect 15092 12684 15596 12740
rect 15652 12684 16380 12740
rect 16436 12684 16446 12740
rect 19954 12684 19964 12740
rect 20020 12684 21644 12740
rect 21700 12684 21710 12740
rect 23090 12684 23100 12740
rect 23156 12684 23884 12740
rect 23940 12684 23950 12740
rect 7026 12516 7036 12572
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7300 12516 7310 12572
rect 12850 12516 12860 12572
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 13124 12516 13134 12572
rect 15092 12404 15148 12684
rect 18674 12516 18684 12572
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18948 12516 18958 12572
rect 24498 12516 24508 12572
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24772 12516 24782 12572
rect 14354 12348 14364 12404
rect 14420 12348 15148 12404
rect 15698 12348 15708 12404
rect 15764 12348 16492 12404
rect 16548 12348 16558 12404
rect 22194 12348 22204 12404
rect 22260 12348 23212 12404
rect 23268 12348 23278 12404
rect 9986 12236 9996 12292
rect 10052 12236 11340 12292
rect 11396 12236 11406 12292
rect 18946 12236 18956 12292
rect 19012 12236 19740 12292
rect 19796 12236 20636 12292
rect 20692 12236 21420 12292
rect 21476 12236 21486 12292
rect 21634 12236 21644 12292
rect 21700 12236 22540 12292
rect 22596 12236 22606 12292
rect 14130 12124 14140 12180
rect 14196 12124 15148 12180
rect 15204 12124 15214 12180
rect 20066 12124 20076 12180
rect 20132 12124 23548 12180
rect 23604 12124 23614 12180
rect 8754 12012 8764 12068
rect 8820 12012 10444 12068
rect 10500 12012 10510 12068
rect 15474 12012 15484 12068
rect 15540 12012 17500 12068
rect 17556 12012 17566 12068
rect 25200 11956 26000 11984
rect 9090 11900 9100 11956
rect 9156 11900 11228 11956
rect 11284 11900 11294 11956
rect 21420 11900 21868 11956
rect 21924 11900 22092 11956
rect 22148 11900 22158 11956
rect 24210 11900 24220 11956
rect 24276 11900 26000 11956
rect 4114 11732 4124 11788
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4388 11732 4398 11788
rect 9938 11732 9948 11788
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 10212 11732 10222 11788
rect 15762 11732 15772 11788
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 16036 11732 16046 11788
rect 21420 11732 21476 11900
rect 25200 11872 26000 11900
rect 21586 11732 21596 11788
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21860 11732 21870 11788
rect 4722 11676 4732 11732
rect 4788 11676 5516 11732
rect 5572 11676 5582 11732
rect 19282 11676 19292 11732
rect 19348 11676 21476 11732
rect 4732 11620 4788 11676
rect 3378 11564 3388 11620
rect 3444 11564 4788 11620
rect 12562 11564 12572 11620
rect 12628 11564 13580 11620
rect 13636 11564 13646 11620
rect 5842 11452 5852 11508
rect 5908 11452 6748 11508
rect 6804 11452 7868 11508
rect 7924 11452 9100 11508
rect 9156 11452 9166 11508
rect 14690 11452 14700 11508
rect 14756 11452 15596 11508
rect 15652 11452 15662 11508
rect 19506 11452 19516 11508
rect 19572 11452 21308 11508
rect 21364 11452 21374 11508
rect 11554 11340 11564 11396
rect 11620 11340 16940 11396
rect 16996 11340 17006 11396
rect 19954 11340 19964 11396
rect 20020 11340 22764 11396
rect 22820 11340 22830 11396
rect 11890 11228 11900 11284
rect 11956 11228 14476 11284
rect 14532 11228 14542 11284
rect 7026 10948 7036 11004
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7300 10948 7310 11004
rect 12850 10948 12860 11004
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 13124 10948 13134 11004
rect 18674 10948 18684 11004
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18948 10948 18958 11004
rect 24498 10948 24508 11004
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24772 10948 24782 11004
rect 15250 10780 15260 10836
rect 15316 10780 16492 10836
rect 16548 10780 16558 10836
rect 20514 10780 20524 10836
rect 20580 10780 22092 10836
rect 22148 10780 22540 10836
rect 22596 10780 22606 10836
rect 3490 10668 3500 10724
rect 3556 10668 4620 10724
rect 4676 10668 9772 10724
rect 9828 10668 9838 10724
rect 1810 10556 1820 10612
rect 1876 10556 4732 10612
rect 4788 10556 5852 10612
rect 5908 10556 5918 10612
rect 20738 10556 20748 10612
rect 20804 10556 21756 10612
rect 21812 10556 22316 10612
rect 22372 10556 22382 10612
rect 21858 10332 21868 10388
rect 21924 10332 22036 10388
rect 4114 10164 4124 10220
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4388 10164 4398 10220
rect 9938 10164 9948 10220
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 10212 10164 10222 10220
rect 15762 10164 15772 10220
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 16036 10164 16046 10220
rect 21586 10164 21596 10220
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21860 10164 21870 10220
rect 21980 10164 22036 10332
rect 17378 10108 17388 10164
rect 17444 10108 21308 10164
rect 21364 10108 21374 10164
rect 21970 10108 21980 10164
rect 22036 10108 22046 10164
rect 18274 9996 18284 10052
rect 18340 9996 19068 10052
rect 19124 9996 19134 10052
rect 25200 9940 26000 9968
rect 10994 9884 11004 9940
rect 11060 9884 12012 9940
rect 12068 9884 12078 9940
rect 24322 9884 24332 9940
rect 24388 9884 26000 9940
rect 25200 9856 26000 9884
rect 20850 9436 20860 9492
rect 20916 9436 21644 9492
rect 21700 9436 23884 9492
rect 23940 9436 24220 9492
rect 24276 9436 24286 9492
rect 7026 9380 7036 9436
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7300 9380 7310 9436
rect 12850 9380 12860 9436
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 13124 9380 13134 9436
rect 18674 9380 18684 9436
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18948 9380 18958 9436
rect 24498 9380 24508 9436
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24772 9380 24782 9436
rect 14802 9212 14812 9268
rect 14868 9212 16604 9268
rect 16660 9212 16670 9268
rect 4610 9100 4620 9156
rect 4676 9100 5404 9156
rect 5460 9100 5470 9156
rect 9986 8988 9996 9044
rect 10052 8988 11004 9044
rect 11060 8988 11070 9044
rect 12786 8988 12796 9044
rect 12852 8988 15484 9044
rect 15540 8988 16044 9044
rect 16100 8988 16110 9044
rect 19730 8988 19740 9044
rect 19796 8988 20300 9044
rect 20356 8988 21084 9044
rect 21140 8988 23324 9044
rect 23380 8988 23390 9044
rect 15698 8764 15708 8820
rect 15764 8764 16828 8820
rect 16884 8764 17388 8820
rect 17444 8764 17454 8820
rect 4114 8596 4124 8652
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4388 8596 4398 8652
rect 9938 8596 9948 8652
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 10212 8596 10222 8652
rect 15762 8596 15772 8652
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 16036 8596 16046 8652
rect 21586 8596 21596 8652
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21860 8596 21870 8652
rect 21410 8540 21420 8596
rect 21476 8540 21486 8596
rect 21420 8484 21476 8540
rect 3602 8428 3612 8484
rect 3668 8428 4620 8484
rect 4676 8428 4686 8484
rect 18498 8428 18508 8484
rect 18564 8428 19628 8484
rect 19684 8428 19694 8484
rect 21420 8428 21644 8484
rect 21700 8428 21710 8484
rect 20962 8316 20972 8372
rect 21028 8316 22092 8372
rect 22148 8316 22158 8372
rect 5618 8204 5628 8260
rect 5684 8204 6860 8260
rect 6916 8204 6926 8260
rect 11554 8204 11564 8260
rect 11620 8204 13692 8260
rect 13748 8204 13758 8260
rect 5842 8092 5852 8148
rect 5908 8092 6636 8148
rect 6692 8092 6702 8148
rect 10882 8092 10892 8148
rect 10948 8092 13468 8148
rect 13524 8092 13534 8148
rect 20066 8092 20076 8148
rect 20132 8092 21084 8148
rect 21140 8092 21532 8148
rect 21588 8092 21598 8148
rect 4386 7980 4396 8036
rect 4452 7980 5740 8036
rect 5796 7980 5806 8036
rect 6290 7980 6300 8036
rect 6356 7980 9436 8036
rect 9492 7980 10444 8036
rect 10500 7980 10510 8036
rect 18274 7980 18284 8036
rect 18340 7980 19572 8036
rect 20402 7980 20412 8036
rect 20468 7980 21308 8036
rect 21364 7980 21374 8036
rect 22866 7980 22876 8036
rect 22932 7980 23324 8036
rect 23380 7980 23390 8036
rect 19516 7924 19572 7980
rect 25200 7924 26000 7952
rect 19506 7868 19516 7924
rect 19572 7868 20524 7924
rect 20580 7868 21420 7924
rect 21476 7868 21486 7924
rect 24892 7868 26000 7924
rect 7026 7812 7036 7868
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7300 7812 7310 7868
rect 12850 7812 12860 7868
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 13124 7812 13134 7868
rect 18674 7812 18684 7868
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18948 7812 18958 7868
rect 24498 7812 24508 7868
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24772 7812 24782 7868
rect 9986 7756 9996 7812
rect 10052 7756 11172 7812
rect 20738 7756 20748 7812
rect 20804 7756 21644 7812
rect 21700 7756 24108 7812
rect 24164 7756 24174 7812
rect 11116 7700 11172 7756
rect 24892 7700 24948 7868
rect 25200 7840 26000 7868
rect 6850 7644 6860 7700
rect 6916 7644 8204 7700
rect 8260 7644 10892 7700
rect 10948 7644 10958 7700
rect 11116 7644 12852 7700
rect 22642 7644 22652 7700
rect 22708 7644 24948 7700
rect 12796 7588 12852 7644
rect 6514 7532 6524 7588
rect 6580 7532 7196 7588
rect 7252 7532 7262 7588
rect 8306 7532 8316 7588
rect 8372 7532 9100 7588
rect 9156 7532 9166 7588
rect 11106 7532 11116 7588
rect 11172 7532 12012 7588
rect 12068 7532 12078 7588
rect 12786 7532 12796 7588
rect 12852 7532 15484 7588
rect 15540 7532 15550 7588
rect 4162 7420 4172 7476
rect 4228 7420 6300 7476
rect 6356 7420 6366 7476
rect 8978 7420 8988 7476
rect 9044 7420 10332 7476
rect 10388 7420 10398 7476
rect 18946 7420 18956 7476
rect 19012 7420 20076 7476
rect 20132 7420 20524 7476
rect 20580 7420 20590 7476
rect 20962 7420 20972 7476
rect 21028 7420 21420 7476
rect 21476 7420 21486 7476
rect 22866 7420 22876 7476
rect 22932 7420 24220 7476
rect 24276 7420 24286 7476
rect 11442 7308 11452 7364
rect 11508 7308 13916 7364
rect 13972 7308 16492 7364
rect 16548 7308 16558 7364
rect 4498 7196 4508 7252
rect 4564 7196 5516 7252
rect 5572 7196 5582 7252
rect 4114 7028 4124 7084
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4388 7028 4398 7084
rect 9938 7028 9948 7084
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 10212 7028 10222 7084
rect 15762 7028 15772 7084
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 16036 7028 16046 7084
rect 21586 7028 21596 7084
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21860 7028 21870 7084
rect 16818 6636 16828 6692
rect 16884 6636 17724 6692
rect 17780 6636 21308 6692
rect 21364 6636 21374 6692
rect 8082 6524 8092 6580
rect 8148 6524 8764 6580
rect 8820 6524 8830 6580
rect 12002 6412 12012 6468
rect 12068 6412 13468 6468
rect 13524 6412 13534 6468
rect 7026 6244 7036 6300
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7300 6244 7310 6300
rect 12850 6244 12860 6300
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 13124 6244 13134 6300
rect 18674 6244 18684 6300
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18948 6244 18958 6300
rect 24498 6244 24508 6300
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24772 6244 24782 6300
rect 22950 5964 22988 6020
rect 23044 5964 23054 6020
rect 25200 5908 26000 5936
rect 14242 5852 14252 5908
rect 14308 5852 16828 5908
rect 16884 5852 16894 5908
rect 23314 5852 23324 5908
rect 23380 5852 26000 5908
rect 25200 5824 26000 5852
rect 4114 5460 4124 5516
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4388 5460 4398 5516
rect 9938 5460 9948 5516
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 10212 5460 10222 5516
rect 15762 5460 15772 5516
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 16036 5460 16046 5516
rect 21586 5460 21596 5516
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21860 5460 21870 5516
rect 20962 5180 20972 5236
rect 21028 5180 23548 5236
rect 23604 5180 23614 5236
rect 7026 4676 7036 4732
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7300 4676 7310 4732
rect 12850 4676 12860 4732
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 13124 4676 13134 4732
rect 18674 4676 18684 4732
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18948 4676 18958 4732
rect 24498 4676 24508 4732
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24772 4676 24782 4732
rect 4114 3892 4124 3948
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4388 3892 4398 3948
rect 9938 3892 9948 3948
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 10212 3892 10222 3948
rect 15762 3892 15772 3948
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 16036 3892 16046 3948
rect 21586 3892 21596 3948
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21860 3892 21870 3948
rect 25200 3892 26000 3920
rect 24210 3836 24220 3892
rect 24276 3836 26000 3892
rect 25200 3808 26000 3836
rect 23426 3388 23436 3444
rect 23492 3388 23884 3444
rect 23940 3388 23950 3444
rect 7026 3108 7036 3164
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7300 3108 7310 3164
rect 12850 3108 12860 3164
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 13124 3108 13134 3164
rect 18674 3108 18684 3164
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18948 3108 18958 3164
rect 24498 3108 24508 3164
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24772 3108 24782 3164
rect 25200 1876 26000 1904
rect 23986 1820 23996 1876
rect 24052 1820 26000 1876
rect 25200 1792 26000 1820
<< via3 >>
rect 4124 22708 4180 22764
rect 4228 22708 4284 22764
rect 4332 22708 4388 22764
rect 9948 22708 10004 22764
rect 10052 22708 10108 22764
rect 10156 22708 10212 22764
rect 15772 22708 15828 22764
rect 15876 22708 15932 22764
rect 15980 22708 16036 22764
rect 21596 22708 21652 22764
rect 21700 22708 21756 22764
rect 21804 22708 21860 22764
rect 7036 21924 7092 21980
rect 7140 21924 7196 21980
rect 7244 21924 7300 21980
rect 12860 21924 12916 21980
rect 12964 21924 13020 21980
rect 13068 21924 13124 21980
rect 18684 21924 18740 21980
rect 18788 21924 18844 21980
rect 18892 21924 18948 21980
rect 24508 21924 24564 21980
rect 24612 21924 24668 21980
rect 24716 21924 24772 21980
rect 4124 21140 4180 21196
rect 4228 21140 4284 21196
rect 4332 21140 4388 21196
rect 9948 21140 10004 21196
rect 10052 21140 10108 21196
rect 10156 21140 10212 21196
rect 15772 21140 15828 21196
rect 15876 21140 15932 21196
rect 15980 21140 16036 21196
rect 21596 21140 21652 21196
rect 21700 21140 21756 21196
rect 21804 21140 21860 21196
rect 23212 20636 23268 20692
rect 7036 20356 7092 20412
rect 7140 20356 7196 20412
rect 7244 20356 7300 20412
rect 12860 20356 12916 20412
rect 12964 20356 13020 20412
rect 13068 20356 13124 20412
rect 18684 20356 18740 20412
rect 18788 20356 18844 20412
rect 18892 20356 18948 20412
rect 24508 20356 24564 20412
rect 24612 20356 24668 20412
rect 24716 20356 24772 20412
rect 4124 19572 4180 19628
rect 4228 19572 4284 19628
rect 4332 19572 4388 19628
rect 9948 19572 10004 19628
rect 10052 19572 10108 19628
rect 10156 19572 10212 19628
rect 15772 19572 15828 19628
rect 15876 19572 15932 19628
rect 15980 19572 16036 19628
rect 21596 19572 21652 19628
rect 21700 19572 21756 19628
rect 21804 19572 21860 19628
rect 7036 18788 7092 18844
rect 7140 18788 7196 18844
rect 7244 18788 7300 18844
rect 12860 18788 12916 18844
rect 12964 18788 13020 18844
rect 13068 18788 13124 18844
rect 18684 18788 18740 18844
rect 18788 18788 18844 18844
rect 18892 18788 18948 18844
rect 24508 18788 24564 18844
rect 24612 18788 24668 18844
rect 24716 18788 24772 18844
rect 4124 18004 4180 18060
rect 4228 18004 4284 18060
rect 4332 18004 4388 18060
rect 9948 18004 10004 18060
rect 10052 18004 10108 18060
rect 10156 18004 10212 18060
rect 15772 18004 15828 18060
rect 15876 18004 15932 18060
rect 15980 18004 16036 18060
rect 21596 18004 21652 18060
rect 21700 18004 21756 18060
rect 21804 18004 21860 18060
rect 7036 17220 7092 17276
rect 7140 17220 7196 17276
rect 7244 17220 7300 17276
rect 12860 17220 12916 17276
rect 12964 17220 13020 17276
rect 13068 17220 13124 17276
rect 18684 17220 18740 17276
rect 18788 17220 18844 17276
rect 18892 17220 18948 17276
rect 24508 17220 24564 17276
rect 24612 17220 24668 17276
rect 24716 17220 24772 17276
rect 4124 16436 4180 16492
rect 4228 16436 4284 16492
rect 4332 16436 4388 16492
rect 9948 16436 10004 16492
rect 10052 16436 10108 16492
rect 10156 16436 10212 16492
rect 15772 16436 15828 16492
rect 15876 16436 15932 16492
rect 15980 16436 16036 16492
rect 21596 16436 21652 16492
rect 21700 16436 21756 16492
rect 21804 16436 21860 16492
rect 7036 15652 7092 15708
rect 7140 15652 7196 15708
rect 7244 15652 7300 15708
rect 12860 15652 12916 15708
rect 12964 15652 13020 15708
rect 13068 15652 13124 15708
rect 18684 15652 18740 15708
rect 18788 15652 18844 15708
rect 18892 15652 18948 15708
rect 24508 15652 24564 15708
rect 24612 15652 24668 15708
rect 24716 15652 24772 15708
rect 22988 15372 23044 15428
rect 4124 14868 4180 14924
rect 4228 14868 4284 14924
rect 4332 14868 4388 14924
rect 9948 14868 10004 14924
rect 10052 14868 10108 14924
rect 10156 14868 10212 14924
rect 15772 14868 15828 14924
rect 15876 14868 15932 14924
rect 15980 14868 16036 14924
rect 21596 14868 21652 14924
rect 21700 14868 21756 14924
rect 21804 14868 21860 14924
rect 7036 14084 7092 14140
rect 7140 14084 7196 14140
rect 7244 14084 7300 14140
rect 12860 14084 12916 14140
rect 12964 14084 13020 14140
rect 13068 14084 13124 14140
rect 18684 14084 18740 14140
rect 18788 14084 18844 14140
rect 18892 14084 18948 14140
rect 24508 14084 24564 14140
rect 24612 14084 24668 14140
rect 24716 14084 24772 14140
rect 4124 13300 4180 13356
rect 4228 13300 4284 13356
rect 4332 13300 4388 13356
rect 9948 13300 10004 13356
rect 10052 13300 10108 13356
rect 10156 13300 10212 13356
rect 15772 13300 15828 13356
rect 15876 13300 15932 13356
rect 15980 13300 16036 13356
rect 21596 13300 21652 13356
rect 21700 13300 21756 13356
rect 21804 13300 21860 13356
rect 7036 12516 7092 12572
rect 7140 12516 7196 12572
rect 7244 12516 7300 12572
rect 12860 12516 12916 12572
rect 12964 12516 13020 12572
rect 13068 12516 13124 12572
rect 18684 12516 18740 12572
rect 18788 12516 18844 12572
rect 18892 12516 18948 12572
rect 24508 12516 24564 12572
rect 24612 12516 24668 12572
rect 24716 12516 24772 12572
rect 23212 12348 23268 12404
rect 4124 11732 4180 11788
rect 4228 11732 4284 11788
rect 4332 11732 4388 11788
rect 9948 11732 10004 11788
rect 10052 11732 10108 11788
rect 10156 11732 10212 11788
rect 15772 11732 15828 11788
rect 15876 11732 15932 11788
rect 15980 11732 16036 11788
rect 21596 11732 21652 11788
rect 21700 11732 21756 11788
rect 21804 11732 21860 11788
rect 7036 10948 7092 11004
rect 7140 10948 7196 11004
rect 7244 10948 7300 11004
rect 12860 10948 12916 11004
rect 12964 10948 13020 11004
rect 13068 10948 13124 11004
rect 18684 10948 18740 11004
rect 18788 10948 18844 11004
rect 18892 10948 18948 11004
rect 24508 10948 24564 11004
rect 24612 10948 24668 11004
rect 24716 10948 24772 11004
rect 4124 10164 4180 10220
rect 4228 10164 4284 10220
rect 4332 10164 4388 10220
rect 9948 10164 10004 10220
rect 10052 10164 10108 10220
rect 10156 10164 10212 10220
rect 15772 10164 15828 10220
rect 15876 10164 15932 10220
rect 15980 10164 16036 10220
rect 21596 10164 21652 10220
rect 21700 10164 21756 10220
rect 21804 10164 21860 10220
rect 7036 9380 7092 9436
rect 7140 9380 7196 9436
rect 7244 9380 7300 9436
rect 12860 9380 12916 9436
rect 12964 9380 13020 9436
rect 13068 9380 13124 9436
rect 18684 9380 18740 9436
rect 18788 9380 18844 9436
rect 18892 9380 18948 9436
rect 24508 9380 24564 9436
rect 24612 9380 24668 9436
rect 24716 9380 24772 9436
rect 4124 8596 4180 8652
rect 4228 8596 4284 8652
rect 4332 8596 4388 8652
rect 9948 8596 10004 8652
rect 10052 8596 10108 8652
rect 10156 8596 10212 8652
rect 15772 8596 15828 8652
rect 15876 8596 15932 8652
rect 15980 8596 16036 8652
rect 21596 8596 21652 8652
rect 21700 8596 21756 8652
rect 21804 8596 21860 8652
rect 7036 7812 7092 7868
rect 7140 7812 7196 7868
rect 7244 7812 7300 7868
rect 12860 7812 12916 7868
rect 12964 7812 13020 7868
rect 13068 7812 13124 7868
rect 18684 7812 18740 7868
rect 18788 7812 18844 7868
rect 18892 7812 18948 7868
rect 24508 7812 24564 7868
rect 24612 7812 24668 7868
rect 24716 7812 24772 7868
rect 4124 7028 4180 7084
rect 4228 7028 4284 7084
rect 4332 7028 4388 7084
rect 9948 7028 10004 7084
rect 10052 7028 10108 7084
rect 10156 7028 10212 7084
rect 15772 7028 15828 7084
rect 15876 7028 15932 7084
rect 15980 7028 16036 7084
rect 21596 7028 21652 7084
rect 21700 7028 21756 7084
rect 21804 7028 21860 7084
rect 7036 6244 7092 6300
rect 7140 6244 7196 6300
rect 7244 6244 7300 6300
rect 12860 6244 12916 6300
rect 12964 6244 13020 6300
rect 13068 6244 13124 6300
rect 18684 6244 18740 6300
rect 18788 6244 18844 6300
rect 18892 6244 18948 6300
rect 24508 6244 24564 6300
rect 24612 6244 24668 6300
rect 24716 6244 24772 6300
rect 22988 5964 23044 6020
rect 4124 5460 4180 5516
rect 4228 5460 4284 5516
rect 4332 5460 4388 5516
rect 9948 5460 10004 5516
rect 10052 5460 10108 5516
rect 10156 5460 10212 5516
rect 15772 5460 15828 5516
rect 15876 5460 15932 5516
rect 15980 5460 16036 5516
rect 21596 5460 21652 5516
rect 21700 5460 21756 5516
rect 21804 5460 21860 5516
rect 7036 4676 7092 4732
rect 7140 4676 7196 4732
rect 7244 4676 7300 4732
rect 12860 4676 12916 4732
rect 12964 4676 13020 4732
rect 13068 4676 13124 4732
rect 18684 4676 18740 4732
rect 18788 4676 18844 4732
rect 18892 4676 18948 4732
rect 24508 4676 24564 4732
rect 24612 4676 24668 4732
rect 24716 4676 24772 4732
rect 4124 3892 4180 3948
rect 4228 3892 4284 3948
rect 4332 3892 4388 3948
rect 9948 3892 10004 3948
rect 10052 3892 10108 3948
rect 10156 3892 10212 3948
rect 15772 3892 15828 3948
rect 15876 3892 15932 3948
rect 15980 3892 16036 3948
rect 21596 3892 21652 3948
rect 21700 3892 21756 3948
rect 21804 3892 21860 3948
rect 7036 3108 7092 3164
rect 7140 3108 7196 3164
rect 7244 3108 7300 3164
rect 12860 3108 12916 3164
rect 12964 3108 13020 3164
rect 13068 3108 13124 3164
rect 18684 3108 18740 3164
rect 18788 3108 18844 3164
rect 18892 3108 18948 3164
rect 24508 3108 24564 3164
rect 24612 3108 24668 3164
rect 24716 3108 24772 3164
<< metal4 >>
rect 4096 22764 4416 22796
rect 4096 22708 4124 22764
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4388 22708 4416 22764
rect 4096 21196 4416 22708
rect 4096 21140 4124 21196
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4388 21140 4416 21196
rect 4096 19628 4416 21140
rect 4096 19572 4124 19628
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4388 19572 4416 19628
rect 4096 18060 4416 19572
rect 4096 18004 4124 18060
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4388 18004 4416 18060
rect 4096 16492 4416 18004
rect 4096 16436 4124 16492
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4388 16436 4416 16492
rect 4096 14924 4416 16436
rect 4096 14868 4124 14924
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4388 14868 4416 14924
rect 4096 13356 4416 14868
rect 4096 13300 4124 13356
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4388 13300 4416 13356
rect 4096 11788 4416 13300
rect 4096 11732 4124 11788
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4388 11732 4416 11788
rect 4096 10220 4416 11732
rect 4096 10164 4124 10220
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4388 10164 4416 10220
rect 4096 8652 4416 10164
rect 4096 8596 4124 8652
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4388 8596 4416 8652
rect 4096 7084 4416 8596
rect 4096 7028 4124 7084
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4388 7028 4416 7084
rect 4096 5516 4416 7028
rect 4096 5460 4124 5516
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4388 5460 4416 5516
rect 4096 3948 4416 5460
rect 4096 3892 4124 3948
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4388 3892 4416 3948
rect 4096 3076 4416 3892
rect 7008 21980 7328 22796
rect 7008 21924 7036 21980
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7300 21924 7328 21980
rect 7008 20412 7328 21924
rect 7008 20356 7036 20412
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7300 20356 7328 20412
rect 7008 18844 7328 20356
rect 7008 18788 7036 18844
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7300 18788 7328 18844
rect 7008 17276 7328 18788
rect 7008 17220 7036 17276
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7300 17220 7328 17276
rect 7008 15708 7328 17220
rect 7008 15652 7036 15708
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7300 15652 7328 15708
rect 7008 14140 7328 15652
rect 7008 14084 7036 14140
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7300 14084 7328 14140
rect 7008 12572 7328 14084
rect 7008 12516 7036 12572
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7300 12516 7328 12572
rect 7008 11004 7328 12516
rect 7008 10948 7036 11004
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7300 10948 7328 11004
rect 7008 9436 7328 10948
rect 7008 9380 7036 9436
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7300 9380 7328 9436
rect 7008 7868 7328 9380
rect 7008 7812 7036 7868
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7300 7812 7328 7868
rect 7008 6300 7328 7812
rect 7008 6244 7036 6300
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7300 6244 7328 6300
rect 7008 4732 7328 6244
rect 7008 4676 7036 4732
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7300 4676 7328 4732
rect 7008 3164 7328 4676
rect 7008 3108 7036 3164
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7300 3108 7328 3164
rect 7008 3076 7328 3108
rect 9920 22764 10240 22796
rect 9920 22708 9948 22764
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 10212 22708 10240 22764
rect 9920 21196 10240 22708
rect 9920 21140 9948 21196
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 10212 21140 10240 21196
rect 9920 19628 10240 21140
rect 9920 19572 9948 19628
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 10212 19572 10240 19628
rect 9920 18060 10240 19572
rect 9920 18004 9948 18060
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 10212 18004 10240 18060
rect 9920 16492 10240 18004
rect 9920 16436 9948 16492
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 10212 16436 10240 16492
rect 9920 14924 10240 16436
rect 9920 14868 9948 14924
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 10212 14868 10240 14924
rect 9920 13356 10240 14868
rect 9920 13300 9948 13356
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 10212 13300 10240 13356
rect 9920 11788 10240 13300
rect 9920 11732 9948 11788
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 10212 11732 10240 11788
rect 9920 10220 10240 11732
rect 9920 10164 9948 10220
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 10212 10164 10240 10220
rect 9920 8652 10240 10164
rect 9920 8596 9948 8652
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 10212 8596 10240 8652
rect 9920 7084 10240 8596
rect 9920 7028 9948 7084
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 10212 7028 10240 7084
rect 9920 5516 10240 7028
rect 9920 5460 9948 5516
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 10212 5460 10240 5516
rect 9920 3948 10240 5460
rect 9920 3892 9948 3948
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 10212 3892 10240 3948
rect 9920 3076 10240 3892
rect 12832 21980 13152 22796
rect 12832 21924 12860 21980
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 13124 21924 13152 21980
rect 12832 20412 13152 21924
rect 12832 20356 12860 20412
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 13124 20356 13152 20412
rect 12832 18844 13152 20356
rect 12832 18788 12860 18844
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 13124 18788 13152 18844
rect 12832 17276 13152 18788
rect 12832 17220 12860 17276
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 13124 17220 13152 17276
rect 12832 15708 13152 17220
rect 12832 15652 12860 15708
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 13124 15652 13152 15708
rect 12832 14140 13152 15652
rect 12832 14084 12860 14140
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 13124 14084 13152 14140
rect 12832 12572 13152 14084
rect 12832 12516 12860 12572
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 13124 12516 13152 12572
rect 12832 11004 13152 12516
rect 12832 10948 12860 11004
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 13124 10948 13152 11004
rect 12832 9436 13152 10948
rect 12832 9380 12860 9436
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 13124 9380 13152 9436
rect 12832 7868 13152 9380
rect 12832 7812 12860 7868
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 13124 7812 13152 7868
rect 12832 6300 13152 7812
rect 12832 6244 12860 6300
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 13124 6244 13152 6300
rect 12832 4732 13152 6244
rect 12832 4676 12860 4732
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 13124 4676 13152 4732
rect 12832 3164 13152 4676
rect 12832 3108 12860 3164
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 13124 3108 13152 3164
rect 12832 3076 13152 3108
rect 15744 22764 16064 22796
rect 15744 22708 15772 22764
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 16036 22708 16064 22764
rect 15744 21196 16064 22708
rect 15744 21140 15772 21196
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 16036 21140 16064 21196
rect 15744 19628 16064 21140
rect 15744 19572 15772 19628
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 16036 19572 16064 19628
rect 15744 18060 16064 19572
rect 15744 18004 15772 18060
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 16036 18004 16064 18060
rect 15744 16492 16064 18004
rect 15744 16436 15772 16492
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 16036 16436 16064 16492
rect 15744 14924 16064 16436
rect 15744 14868 15772 14924
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 16036 14868 16064 14924
rect 15744 13356 16064 14868
rect 15744 13300 15772 13356
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 16036 13300 16064 13356
rect 15744 11788 16064 13300
rect 15744 11732 15772 11788
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 16036 11732 16064 11788
rect 15744 10220 16064 11732
rect 15744 10164 15772 10220
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 16036 10164 16064 10220
rect 15744 8652 16064 10164
rect 15744 8596 15772 8652
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 16036 8596 16064 8652
rect 15744 7084 16064 8596
rect 15744 7028 15772 7084
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 16036 7028 16064 7084
rect 15744 5516 16064 7028
rect 15744 5460 15772 5516
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 16036 5460 16064 5516
rect 15744 3948 16064 5460
rect 15744 3892 15772 3948
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 16036 3892 16064 3948
rect 15744 3076 16064 3892
rect 18656 21980 18976 22796
rect 18656 21924 18684 21980
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18948 21924 18976 21980
rect 18656 20412 18976 21924
rect 18656 20356 18684 20412
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18948 20356 18976 20412
rect 18656 18844 18976 20356
rect 18656 18788 18684 18844
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18948 18788 18976 18844
rect 18656 17276 18976 18788
rect 18656 17220 18684 17276
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18948 17220 18976 17276
rect 18656 15708 18976 17220
rect 18656 15652 18684 15708
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18948 15652 18976 15708
rect 18656 14140 18976 15652
rect 18656 14084 18684 14140
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18948 14084 18976 14140
rect 18656 12572 18976 14084
rect 18656 12516 18684 12572
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18948 12516 18976 12572
rect 18656 11004 18976 12516
rect 18656 10948 18684 11004
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18948 10948 18976 11004
rect 18656 9436 18976 10948
rect 18656 9380 18684 9436
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18948 9380 18976 9436
rect 18656 7868 18976 9380
rect 18656 7812 18684 7868
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18948 7812 18976 7868
rect 18656 6300 18976 7812
rect 18656 6244 18684 6300
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18948 6244 18976 6300
rect 18656 4732 18976 6244
rect 18656 4676 18684 4732
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18948 4676 18976 4732
rect 18656 3164 18976 4676
rect 18656 3108 18684 3164
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18948 3108 18976 3164
rect 18656 3076 18976 3108
rect 21568 22764 21888 22796
rect 21568 22708 21596 22764
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21860 22708 21888 22764
rect 21568 21196 21888 22708
rect 21568 21140 21596 21196
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21860 21140 21888 21196
rect 21568 19628 21888 21140
rect 24480 21980 24800 22796
rect 24480 21924 24508 21980
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24772 21924 24800 21980
rect 21568 19572 21596 19628
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21860 19572 21888 19628
rect 21568 18060 21888 19572
rect 21568 18004 21596 18060
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21860 18004 21888 18060
rect 21568 16492 21888 18004
rect 21568 16436 21596 16492
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21860 16436 21888 16492
rect 21568 14924 21888 16436
rect 23212 20692 23268 20702
rect 21568 14868 21596 14924
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21860 14868 21888 14924
rect 21568 13356 21888 14868
rect 21568 13300 21596 13356
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21860 13300 21888 13356
rect 21568 11788 21888 13300
rect 21568 11732 21596 11788
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21860 11732 21888 11788
rect 21568 10220 21888 11732
rect 21568 10164 21596 10220
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21860 10164 21888 10220
rect 21568 8652 21888 10164
rect 21568 8596 21596 8652
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21860 8596 21888 8652
rect 21568 7084 21888 8596
rect 21568 7028 21596 7084
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21860 7028 21888 7084
rect 21568 5516 21888 7028
rect 22988 15428 23044 15438
rect 22988 6020 23044 15372
rect 23212 12404 23268 20636
rect 23212 12338 23268 12348
rect 24480 20412 24800 21924
rect 24480 20356 24508 20412
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24772 20356 24800 20412
rect 24480 18844 24800 20356
rect 24480 18788 24508 18844
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24772 18788 24800 18844
rect 24480 17276 24800 18788
rect 24480 17220 24508 17276
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24772 17220 24800 17276
rect 24480 15708 24800 17220
rect 24480 15652 24508 15708
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24772 15652 24800 15708
rect 24480 14140 24800 15652
rect 24480 14084 24508 14140
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24772 14084 24800 14140
rect 24480 12572 24800 14084
rect 24480 12516 24508 12572
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24772 12516 24800 12572
rect 22988 5954 23044 5964
rect 24480 11004 24800 12516
rect 24480 10948 24508 11004
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24772 10948 24800 11004
rect 24480 9436 24800 10948
rect 24480 9380 24508 9436
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24772 9380 24800 9436
rect 24480 7868 24800 9380
rect 24480 7812 24508 7868
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24772 7812 24800 7868
rect 24480 6300 24800 7812
rect 24480 6244 24508 6300
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24772 6244 24800 6300
rect 21568 5460 21596 5516
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21860 5460 21888 5516
rect 21568 3948 21888 5460
rect 21568 3892 21596 3948
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21860 3892 21888 3948
rect 21568 3076 21888 3892
rect 24480 4732 24800 6244
rect 24480 4676 24508 4732
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24772 4676 24800 4732
rect 24480 3164 24800 4676
rect 24480 3108 24508 3164
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24772 3108 24800 3164
rect 24480 3076 24800 3108
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _177_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 21168 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _178_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 20048 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _179_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 21056 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _180_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 21280 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _181_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 20944 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _182_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 22848 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _183_
timestamp 1694700623
transform 1 0 21280 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _184_
timestamp 1694700623
transform -1 0 17920 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _185_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 19040 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _186_
timestamp 1694700623
transform -1 0 20272 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _187_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 19600 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _188_
timestamp 1694700623
transform 1 0 17248 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _189_
timestamp 1694700623
transform -1 0 19600 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 20944 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _191_
timestamp 1694700623
transform -1 0 20384 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _192_
timestamp 1694700623
transform -1 0 18704 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _193_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 22064 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _194_
timestamp 1694700623
transform -1 0 22512 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1694700623
transform -1 0 19712 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _196_
timestamp 1694700623
transform 1 0 19712 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _197_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 22064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _198_
timestamp 1694700623
transform -1 0 20272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _199_
timestamp 1694700623
transform -1 0 20272 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1694700623
transform 1 0 20272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _201_
timestamp 1694700623
transform -1 0 22064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _202_
timestamp 1694700623
transform -1 0 22960 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _203_
timestamp 1694700623
transform -1 0 20608 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1694700623
transform -1 0 20608 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _205_
timestamp 1694700623
transform -1 0 17248 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _206_
timestamp 1694700623
transform 1 0 17920 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _207_
timestamp 1694700623
transform 1 0 19040 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _208_
timestamp 1694700623
transform -1 0 20048 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _209_
timestamp 1694700623
transform 1 0 21616 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _210_
timestamp 1694700623
transform -1 0 23072 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _211_
timestamp 1694700623
transform -1 0 21616 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _212_
timestamp 1694700623
transform -1 0 16688 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _213_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _214_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 12208 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _215_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 15232 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _216_
timestamp 1694700623
transform 1 0 16016 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _217_
timestamp 1694700623
transform 1 0 13328 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _218_
timestamp 1694700623
transform -1 0 12768 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _219_
timestamp 1694700623
transform -1 0 11088 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _220_
timestamp 1694700623
transform -1 0 16240 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _221_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 10192 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _222_
timestamp 1694700623
transform 1 0 9408 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _223_
timestamp 1694700623
transform 1 0 8288 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _224_
timestamp 1694700623
transform -1 0 14224 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _225_
timestamp 1694700623
transform 1 0 4256 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _226_
timestamp 1694700623
transform 1 0 2912 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _227_
timestamp 1694700623
transform 1 0 2016 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _228_
timestamp 1694700623
transform 1 0 5488 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _229_
timestamp 1694700623
transform 1 0 3024 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _230_
timestamp 1694700623
transform 1 0 2016 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _231_
timestamp 1694700623
transform 1 0 6944 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _232_
timestamp 1694700623
transform 1 0 5264 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _233_
timestamp 1694700623
transform -1 0 4704 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _234_
timestamp 1694700623
transform 1 0 9744 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _235_
timestamp 1694700623
transform 1 0 8512 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _236_
timestamp 1694700623
transform -1 0 8288 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _237_
timestamp 1694700623
transform -1 0 12656 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _238_
timestamp 1694700623
transform 1 0 11424 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _239_
timestamp 1694700623
transform 1 0 11536 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _240_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 15680 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _241_
timestamp 1694700623
transform 1 0 16240 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _242_
timestamp 1694700623
transform 1 0 14672 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _243_
timestamp 1694700623
transform 1 0 16240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _244_
timestamp 1694700623
transform 1 0 15792 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _245_
timestamp 1694700623
transform 1 0 17248 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _246_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 17024 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _247_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 15008 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _248_
timestamp 1694700623
transform -1 0 17696 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _249_
timestamp 1694700623
transform 1 0 15904 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _250_
timestamp 1694700623
transform 1 0 15680 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _251_
timestamp 1694700623
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _252_
timestamp 1694700623
transform 1 0 14448 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _253_
timestamp 1694700623
transform 1 0 15344 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _254_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 14000 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _255_
timestamp 1694700623
transform -1 0 15344 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _256_
timestamp 1694700623
transform -1 0 12432 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _257_
timestamp 1694700623
transform -1 0 15456 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _258_
timestamp 1694700623
transform 1 0 14000 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _259_
timestamp 1694700623
transform 1 0 15232 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _260_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 14112 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _261_
timestamp 1694700623
transform 1 0 13776 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _262_
timestamp 1694700623
transform 1 0 13664 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _263_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 14112 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _264_
timestamp 1694700623
transform 1 0 15008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _265_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 11760 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _266_
timestamp 1694700623
transform -1 0 12432 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _267_
timestamp 1694700623
transform -1 0 24304 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _268_
timestamp 1694700623
transform 1 0 22400 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _269_
timestamp 1694700623
transform -1 0 23744 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _270_
timestamp 1694700623
transform -1 0 23632 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _271_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 20272 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _272_
timestamp 1694700623
transform -1 0 24304 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _273_
timestamp 1694700623
transform -1 0 24416 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _274_
timestamp 1694700623
transform -1 0 24080 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _275_
timestamp 1694700623
transform 1 0 22512 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _276_
timestamp 1694700623
transform -1 0 24416 0 -1 12544
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _277_
timestamp 1694700623
transform 1 0 22960 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _278_
timestamp 1694700623
transform 1 0 22960 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _279_
timestamp 1694700623
transform -1 0 24304 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _280_
timestamp 1694700623
transform -1 0 24304 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _281_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 22400 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _282_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 15904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _283_
timestamp 1694700623
transform 1 0 14000 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _284_
timestamp 1694700623
transform 1 0 14448 0 1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _285_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 22848 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _286_
timestamp 1694700623
transform -1 0 11760 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _287_
timestamp 1694700623
transform 1 0 8064 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _288_
timestamp 1694700623
transform 1 0 7840 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _289_
timestamp 1694700623
transform 1 0 10304 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _290_
timestamp 1694700623
transform 1 0 6720 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _291_
timestamp 1694700623
transform 1 0 7728 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _292_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 9968 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _293_
timestamp 1694700623
transform 1 0 7952 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _294_
timestamp 1694700623
transform 1 0 8960 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _295_
timestamp 1694700623
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _296_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 10528 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _297_
timestamp 1694700623
transform -1 0 7840 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _298_
timestamp 1694700623
transform 1 0 13216 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _299_
timestamp 1694700623
transform 1 0 8512 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _300_
timestamp 1694700623
transform -1 0 8512 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _301_
timestamp 1694700623
transform 1 0 5936 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _302_
timestamp 1694700623
transform -1 0 4928 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _303_
timestamp 1694700623
transform -1 0 5264 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _304_
timestamp 1694700623
transform -1 0 9184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _305_
timestamp 1694700623
transform -1 0 7504 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _306_
timestamp 1694700623
transform -1 0 4032 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _307_
timestamp 1694700623
transform 1 0 2688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _308_
timestamp 1694700623
transform -1 0 13216 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _309_
timestamp 1694700623
transform -1 0 5824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _310_
timestamp 1694700623
transform 1 0 10192 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _311_
timestamp 1694700623
transform -1 0 10976 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _312_
timestamp 1694700623
transform 1 0 9968 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _313_
timestamp 1694700623
transform -1 0 10192 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _314_
timestamp 1694700623
transform 1 0 11088 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _315_
timestamp 1694700623
transform 1 0 11200 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _316_
timestamp 1694700623
transform -1 0 6160 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _317_
timestamp 1694700623
transform 1 0 3920 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _318_
timestamp 1694700623
transform -1 0 4032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _319_
timestamp 1694700623
transform 1 0 3584 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _320_
timestamp 1694700623
transform 1 0 4144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _321_
timestamp 1694700623
transform -1 0 8288 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _322_
timestamp 1694700623
transform 1 0 7616 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _323_
timestamp 1694700623
transform 1 0 5488 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _324_
timestamp 1694700623
transform 1 0 5040 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _325_
timestamp 1694700623
transform -1 0 6832 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _326_
timestamp 1694700623
transform 1 0 5712 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _327_
timestamp 1694700623
transform 1 0 4816 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _328_
timestamp 1694700623
transform 1 0 6048 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _329_
timestamp 1694700623
transform -1 0 2688 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _330_
timestamp 1694700623
transform 1 0 5600 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _331_
timestamp 1694700623
transform -1 0 5264 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _332_
timestamp 1694700623
transform 1 0 2464 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _333_
timestamp 1694700623
transform 1 0 2912 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _334_
timestamp 1694700623
transform -1 0 8848 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _335_
timestamp 1694700623
transform 1 0 2240 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _336_
timestamp 1694700623
transform -1 0 3808 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _337_
timestamp 1694700623
transform -1 0 2464 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _338_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2128 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _339_
timestamp 1694700623
transform 1 0 5712 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _340_
timestamp 1694700623
transform 1 0 6048 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _341_
timestamp 1694700623
transform -1 0 7392 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _342_
timestamp 1694700623
transform 1 0 7728 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _343_
timestamp 1694700623
transform 1 0 9408 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _344_
timestamp 1694700623
transform -1 0 20048 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _345_
timestamp 1694700623
transform -1 0 22400 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _346_
timestamp 1694700623
transform -1 0 16800 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _347_
timestamp 1694700623
transform 1 0 16688 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _348_
timestamp 1694700623
transform -1 0 19264 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _349_
timestamp 1694700623
transform -1 0 18704 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _350_
timestamp 1694700623
transform -1 0 21168 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _351_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 17920 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _352_
timestamp 1694700623
transform 1 0 19376 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _353_
timestamp 1694700623
transform 1 0 19264 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _354_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 8960 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _355_
timestamp 1694700623
transform 1 0 17248 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _356_
timestamp 1694700623
transform 1 0 17584 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _357_
timestamp 1694700623
transform 1 0 21168 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _358_
timestamp 1694700623
transform 1 0 21168 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _359_
timestamp 1694700623
transform 1 0 17248 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _360_
timestamp 1694700623
transform 1 0 17248 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _361_
timestamp 1694700623
transform 1 0 20496 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _362_
timestamp 1694700623
transform 1 0 17248 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _363_
timestamp 1694700623
transform 1 0 20832 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _364_
timestamp 1694700623
transform 1 0 17248 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _365_
timestamp 1694700623
transform 1 0 17696 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _366_
timestamp 1694700623
transform 1 0 20944 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _367_
timestamp 1694700623
transform 1 0 7728 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _368_
timestamp 1694700623
transform 1 0 5712 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _369_
timestamp 1694700623
transform 1 0 1792 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _370_
timestamp 1694700623
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _371_
timestamp 1694700623
transform 1 0 5936 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _372_
timestamp 1694700623
transform 1 0 11088 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _373_
timestamp 1694700623
transform 1 0 8960 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _374_
timestamp 1694700623
transform 1 0 1568 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _375_
timestamp 1694700623
transform 1 0 1568 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _376_
timestamp 1694700623
transform 1 0 2688 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _377_
timestamp 1694700623
transform 1 0 5936 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _378_
timestamp 1694700623
transform -1 0 14448 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _379_
timestamp 1694700623
transform -1 0 15904 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _380_
timestamp 1694700623
transform 1 0 15344 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _381_
timestamp 1694700623
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _382_
timestamp 1694700623
transform 1 0 4816 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _383_
timestamp 1694700623
transform 1 0 3248 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _384_
timestamp 1694700623
transform 1 0 7168 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _385_
timestamp 1694700623
transform -1 0 17472 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _386_
timestamp 1694700623
transform -1 0 17024 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _387_
timestamp 1694700623
transform 1 0 11200 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _388_
timestamp 1694700623
transform 1 0 10752 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _389_
timestamp 1694700623
transform 1 0 12992 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _390_
timestamp 1694700623
transform 1 0 9744 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _391_
timestamp 1694700623
transform 1 0 4592 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__A1
timestamp 1694700623
transform -1 0 10192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__S
timestamp 1694700623
transform -1 0 7840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A2
timestamp 1694700623
transform 1 0 8512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1694700623
transform -1 0 12656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1694700623
transform -1 0 23520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1694700623
transform -1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1694700623
transform -1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1694700623
transform -1 0 23744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1694700623
transform -1 0 22960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1694700623
transform -1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1694700623
transform -1 0 22960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1694700623
transform -1 0 19040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1694700623
transform -1 0 24416 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1694700623
transform -1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1694700623
transform -1 0 22960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1694700623
transform -1 0 21728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1694700623
transform -1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 13328 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1694700623
transform -1 0 11760 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1694700623
transform -1 0 13104 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1694700623
transform 1 0 15344 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1694700623
transform 1 0 17248 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1694700623
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1694700623
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1694700623
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1694700623
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_188 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 22400 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1694700623
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1694700623
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1694700623
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_174
timestamp 1694700623
transform 1 0 20832 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_190
timestamp 1694700623
transform 1 0 22624 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1694700623
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1694700623
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1694700623
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1694700623
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1694700623
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1694700623
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_205
timestamp 1694700623
transform 1 0 24304 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_2
timestamp 1694700623
transform 1 0 1568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_10 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1694700623
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_117
timestamp 1694700623
transform 1 0 14448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_133
timestamp 1694700623
transform 1 0 16240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1694700623
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1694700623
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_142
timestamp 1694700623
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_158
timestamp 1694700623
transform 1 0 19040 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_166
timestamp 1694700623
transform 1 0 19936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_170
timestamp 1694700623
transform 1 0 20384 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_177
timestamp 1694700623
transform 1 0 21168 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_185
timestamp 1694700623
transform 1 0 22064 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_189
timestamp 1694700623
transform 1 0 22512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_205
timestamp 1694700623
transform 1 0 24304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_2
timestamp 1694700623
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_18
timestamp 1694700623
transform 1 0 3360 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_22
timestamp 1694700623
transform 1 0 3808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_30
timestamp 1694700623
transform 1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1694700623
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1694700623
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_53
timestamp 1694700623
transform 1 0 7280 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_55
timestamp 1694700623
transform 1 0 7504 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_62
timestamp 1694700623
transform 1 0 8288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_79
timestamp 1694700623
transform 1 0 10192 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_87
timestamp 1694700623
transform 1 0 11088 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_97
timestamp 1694700623
transform 1 0 12208 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_107
timestamp 1694700623
transform 1 0 13328 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_139
timestamp 1694700623
transform 1 0 16912 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_143
timestamp 1694700623
transform 1 0 17360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1694700623
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1694700623
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_12
timestamp 1694700623
transform 1 0 2688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_14
timestamp 1694700623
transform 1 0 2912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_30
timestamp 1694700623
transform 1 0 4704 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_34
timestamp 1694700623
transform 1 0 5152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_65
timestamp 1694700623
transform 1 0 8624 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1694700623
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1694700623
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1694700623
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_105
timestamp 1694700623
transform 1 0 13104 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_109
timestamp 1694700623
transform 1 0 13552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1694700623
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_146
timestamp 1694700623
transform 1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_167
timestamp 1694700623
transform 1 0 20048 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_175
timestamp 1694700623
transform 1 0 20944 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_184
timestamp 1694700623
transform 1 0 21952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_31
timestamp 1694700623
transform 1 0 4816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_52
timestamp 1694700623
transform 1 0 7168 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_68
timestamp 1694700623
transform 1 0 8960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_70
timestamp 1694700623
transform 1 0 9184 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_79
timestamp 1694700623
transform 1 0 10192 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_83
timestamp 1694700623
transform 1 0 10640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_85
timestamp 1694700623
transform 1 0 10864 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1694700623
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_115
timestamp 1694700623
transform 1 0 14224 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_123
timestamp 1694700623
transform 1 0 15120 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_132
timestamp 1694700623
transform 1 0 16128 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_148
timestamp 1694700623
transform 1 0 17920 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_155
timestamp 1694700623
transform 1 0 18704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_159
timestamp 1694700623
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_187
timestamp 1694700623
transform 1 0 22288 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_205
timestamp 1694700623
transform 1 0 24304 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1694700623
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_18
timestamp 1694700623
transform 1 0 3360 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_87
timestamp 1694700623
transform 1 0 11088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_95
timestamp 1694700623
transform 1 0 11984 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_99
timestamp 1694700623
transform 1 0 12432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1694700623
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_171
timestamp 1694700623
transform 1 0 20496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_186
timestamp 1694700623
transform 1 0 22176 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_190
timestamp 1694700623
transform 1 0 22624 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_203
timestamp 1694700623
transform 1 0 24080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_205
timestamp 1694700623
transform 1 0 24304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_31
timestamp 1694700623
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1694700623
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_45
timestamp 1694700623
transform 1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_47
timestamp 1694700623
transform 1 0 6608 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_54
timestamp 1694700623
transform 1 0 7392 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_97
timestamp 1694700623
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1694700623
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_115
timestamp 1694700623
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_127
timestamp 1694700623
transform 1 0 15568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_143
timestamp 1694700623
transform 1 0 17360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_147
timestamp 1694700623
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_155
timestamp 1694700623
transform 1 0 18704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_157
timestamp 1694700623
transform 1 0 18928 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2
timestamp 1694700623
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_12
timestamp 1694700623
transform 1 0 2688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_58
timestamp 1694700623
transform 1 0 7840 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1694700623
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1694700623
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1694700623
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_97
timestamp 1694700623
transform 1 0 12208 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_113
timestamp 1694700623
transform 1 0 14000 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_121
timestamp 1694700623
transform 1 0 14896 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1694700623
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_171
timestamp 1694700623
transform 1 0 20496 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_192
timestamp 1694700623
transform 1 0 22848 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_205
timestamp 1694700623
transform 1 0 24304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1694700623
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1694700623
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1694700623
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_41
timestamp 1694700623
transform 1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_93
timestamp 1694700623
transform 1 0 11760 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1694700623
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_122
timestamp 1694700623
transform 1 0 15008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_124
timestamp 1694700623
transform 1 0 15232 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_201
timestamp 1694700623
transform 1 0 23856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_203
timestamp 1694700623
transform 1 0 24080 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1694700623
transform 1 0 1568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_33
timestamp 1694700623
transform 1 0 5040 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_37
timestamp 1694700623
transform 1 0 5488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1694700623
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_116
timestamp 1694700623
transform 1 0 14336 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_120
timestamp 1694700623
transform 1 0 14784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_137
timestamp 1694700623
transform 1 0 16688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1694700623
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_146
timestamp 1694700623
transform 1 0 17696 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_150
timestamp 1694700623
transform 1 0 18144 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_2
timestamp 1694700623
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_10
timestamp 1694700623
transform 1 0 2464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_20
timestamp 1694700623
transform 1 0 3584 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_28
timestamp 1694700623
transform 1 0 4480 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1694700623
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_41
timestamp 1694700623
transform 1 0 5936 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_48
timestamp 1694700623
transform 1 0 6720 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_56
timestamp 1694700623
transform 1 0 7616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_86
timestamp 1694700623
transform 1 0 10976 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_94
timestamp 1694700623
transform 1 0 11872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1694700623
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1694700623
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_144
timestamp 1694700623
transform 1 0 17472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_152
timestamp 1694700623
transform 1 0 18368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_177
timestamp 1694700623
transform 1 0 21168 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1694700623
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_199
timestamp 1694700623
transform 1 0 23632 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_47
timestamp 1694700623
transform 1 0 6608 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_63
timestamp 1694700623
transform 1 0 8400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1694700623
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1694700623
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_78
timestamp 1694700623
transform 1 0 10080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_86
timestamp 1694700623
transform 1 0 10976 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_123
timestamp 1694700623
transform 1 0 15120 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_132
timestamp 1694700623
transform 1 0 16128 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1694700623
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1694700623
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_2
timestamp 1694700623
transform 1 0 1568 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_6
timestamp 1694700623
transform 1 0 2016 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_22
timestamp 1694700623
transform 1 0 3808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_24
timestamp 1694700623
transform 1 0 4032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_33
timestamp 1694700623
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1694700623
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_41
timestamp 1694700623
transform 1 0 5936 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_54
timestamp 1694700623
transform 1 0 7392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_56
timestamp 1694700623
transform 1 0 7616 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_65
timestamp 1694700623
transform 1 0 8624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_67
timestamp 1694700623
transform 1 0 8848 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_97
timestamp 1694700623
transform 1 0 12208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1694700623
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1694700623
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_67
timestamp 1694700623
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1694700623
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1694700623
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_88
timestamp 1694700623
transform 1 0 11200 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_96
timestamp 1694700623
transform 1 0 12096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_100
timestamp 1694700623
transform 1 0 12544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_102
timestamp 1694700623
transform 1 0 12768 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1694700623
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1694700623
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1694700623
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_160
timestamp 1694700623
transform 1 0 19264 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2
timestamp 1694700623
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_6
timestamp 1694700623
transform 1 0 2016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_33
timestamp 1694700623
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1694700623
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_46
timestamp 1694700623
transform 1 0 6496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_50
timestamp 1694700623
transform 1 0 6944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_81
timestamp 1694700623
transform 1 0 10416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_85
timestamp 1694700623
transform 1 0 10864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_93
timestamp 1694700623
transform 1 0 11760 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_99
timestamp 1694700623
transform 1 0 12432 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1694700623
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1694700623
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_115
timestamp 1694700623
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_160
timestamp 1694700623
transform 1 0 19264 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1694700623
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1694700623
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1694700623
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1694700623
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1694700623
transform 1 0 22288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1694700623
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_18
timestamp 1694700623
transform 1 0 3360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_26
timestamp 1694700623
transform 1 0 4256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_30
timestamp 1694700623
transform 1 0 4704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_32
timestamp 1694700623
transform 1 0 4928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_49
timestamp 1694700623
transform 1 0 6832 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_51
timestamp 1694700623
transform 1 0 7056 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_62
timestamp 1694700623
transform 1 0 8288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1694700623
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_82
timestamp 1694700623
transform 1 0 10528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_117
timestamp 1694700623
transform 1 0 14448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_125
timestamp 1694700623
transform 1 0 15344 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_129
timestamp 1694700623
transform 1 0 15792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_131
timestamp 1694700623
transform 1 0 16016 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1694700623
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_205
timestamp 1694700623
transform 1 0 24304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2
timestamp 1694700623
transform 1 0 1568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_24
timestamp 1694700623
transform 1 0 4032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_26
timestamp 1694700623
transform 1 0 4256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1694700623
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1694700623
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1694700623
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1694700623
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_118
timestamp 1694700623
transform 1 0 14560 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_126
timestamp 1694700623
transform 1 0 15456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_128
timestamp 1694700623
transform 1 0 15680 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1694700623
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_205
timestamp 1694700623
transform 1 0 24304 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1694700623
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_10
timestamp 1694700623
transform 1 0 2464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_14
timestamp 1694700623
transform 1 0 2912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_16
timestamp 1694700623
transform 1 0 3136 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_40
timestamp 1694700623
transform 1 0 5824 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_56
timestamp 1694700623
transform 1 0 7616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_58
timestamp 1694700623
transform 1 0 7840 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_99
timestamp 1694700623
transform 1 0 12432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_112
timestamp 1694700623
transform 1 0 13888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_130
timestamp 1694700623
transform 1 0 15904 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1694700623
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_154
timestamp 1694700623
transform 1 0 18592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_158
timestamp 1694700623
transform 1 0 19040 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_172
timestamp 1694700623
transform 1 0 20608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_203
timestamp 1694700623
transform 1 0 24080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_205
timestamp 1694700623
transform 1 0 24304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1694700623
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_53
timestamp 1694700623
transform 1 0 7280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_55
timestamp 1694700623
transform 1 0 7504 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_73
timestamp 1694700623
transform 1 0 9520 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_92
timestamp 1694700623
transform 1 0 11648 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1694700623
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1694700623
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1694700623
transform 1 0 13552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_134
timestamp 1694700623
transform 1 0 16352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1694700623
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1694700623
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1694700623
transform 1 0 21392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2
timestamp 1694700623
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_10
timestamp 1694700623
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_14
timestamp 1694700623
transform 1 0 2912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_16
timestamp 1694700623
transform 1 0 3136 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_46
timestamp 1694700623
transform 1 0 6496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1694700623
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_79
timestamp 1694700623
transform 1 0 10192 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_119
timestamp 1694700623
transform 1 0 14672 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_126
timestamp 1694700623
transform 1 0 15456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_147
timestamp 1694700623
transform 1 0 17808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_155
timestamp 1694700623
transform 1 0 18704 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_159
timestamp 1694700623
transform 1 0 19152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_172
timestamp 1694700623
transform 1 0 20608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_174
timestamp 1694700623
transform 1 0 20832 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_188
timestamp 1694700623
transform 1 0 22400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_190
timestamp 1694700623
transform 1 0 22624 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_205
timestamp 1694700623
transform 1 0 24304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1694700623
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1694700623
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_37
timestamp 1694700623
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_53
timestamp 1694700623
transform 1 0 7280 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_86
timestamp 1694700623
transform 1 0 10976 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1694700623
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1694700623
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1694700623
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1694700623
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_154
timestamp 1694700623
transform 1 0 18592 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_170
timestamp 1694700623
transform 1 0 20384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1694700623
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1694700623
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_181
timestamp 1694700623
transform 1 0 21616 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_2
timestamp 1694700623
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_18
timestamp 1694700623
transform 1 0 3360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_26
timestamp 1694700623
transform 1 0 4256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_30
timestamp 1694700623
transform 1 0 4704 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1694700623
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1694700623
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_74
timestamp 1694700623
transform 1 0 9632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_133
timestamp 1694700623
transform 1 0 16240 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1694700623
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1694700623
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1694700623
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_204
timestamp 1694700623
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1694700623
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_36
timestamp 1694700623
transform 1 0 5376 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_70
timestamp 1694700623
transform 1 0 9184 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_86
timestamp 1694700623
transform 1 0 10976 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_94
timestamp 1694700623
transform 1 0 11872 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_98
timestamp 1694700623
transform 1 0 12320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_110
timestamp 1694700623
transform 1 0 13664 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_126
timestamp 1694700623
transform 1 0 15456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_134
timestamp 1694700623
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_138
timestamp 1694700623
transform 1 0 16800 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_154
timestamp 1694700623
transform 1 0 18592 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1694700623
transform -1 0 24192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1694700623
transform 1 0 20608 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1694700623
transform 1 0 19712 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1694700623
transform -1 0 24416 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1694700623
transform 1 0 23072 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1694700623
transform 1 0 22400 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1694700623
transform -1 0 24416 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1694700623
transform -1 0 24416 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1694700623
transform -1 0 24416 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1694700623
transform -1 0 24416 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1694700623
transform -1 0 24416 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1694700623
transform 1 0 21728 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1694700623
transform 1 0 12992 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 21280 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_25 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 24640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_26
timestamp 1694700623
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_27
timestamp 1694700623
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 24640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_28
timestamp 1694700623
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_29
timestamp 1694700623
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_30
timestamp 1694700623
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_31
timestamp 1694700623
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 24640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_32
timestamp 1694700623
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_33
timestamp 1694700623
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 24640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_34
timestamp 1694700623
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_35
timestamp 1694700623
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 24640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_36
timestamp 1694700623
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_37
timestamp 1694700623
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 24640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_38
timestamp 1694700623
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_39
timestamp 1694700623
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_40
timestamp 1694700623
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_41
timestamp 1694700623
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 24640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_42
timestamp 1694700623
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_43
timestamp 1694700623
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 24640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_44
timestamp 1694700623
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_45
timestamp 1694700623
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_46
timestamp 1694700623
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_47
timestamp 1694700623
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_48
timestamp 1694700623
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_49
timestamp 1694700623
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 24640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_50 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_51
timestamp 1694700623
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_52
timestamp 1694700623
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_53
timestamp 1694700623
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_54
timestamp 1694700623
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_55
timestamp 1694700623
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_56
timestamp 1694700623
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_57
timestamp 1694700623
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1694700623
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1694700623
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_60
timestamp 1694700623
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1694700623
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1694700623
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_63
timestamp 1694700623
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_64
timestamp 1694700623
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_65
timestamp 1694700623
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_66
timestamp 1694700623
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_67
timestamp 1694700623
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_68
timestamp 1694700623
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_69
timestamp 1694700623
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_70
timestamp 1694700623
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_71
timestamp 1694700623
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_72
timestamp 1694700623
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_73
timestamp 1694700623
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_74
timestamp 1694700623
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_75
timestamp 1694700623
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_76
timestamp 1694700623
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_77
timestamp 1694700623
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_78
timestamp 1694700623
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_79
timestamp 1694700623
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_80
timestamp 1694700623
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_81
timestamp 1694700623
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_82
timestamp 1694700623
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_83
timestamp 1694700623
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_84
timestamp 1694700623
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_85
timestamp 1694700623
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_86
timestamp 1694700623
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_87
timestamp 1694700623
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_88
timestamp 1694700623
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_89
timestamp 1694700623
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_90
timestamp 1694700623
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_91
timestamp 1694700623
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_92
timestamp 1694700623
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_93
timestamp 1694700623
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_94
timestamp 1694700623
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_95
timestamp 1694700623
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_96
timestamp 1694700623
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_97
timestamp 1694700623
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_98
timestamp 1694700623
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_99
timestamp 1694700623
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_100
timestamp 1694700623
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_101
timestamp 1694700623
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_102
timestamp 1694700623
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_103
timestamp 1694700623
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_104
timestamp 1694700623
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_105
timestamp 1694700623
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_106
timestamp 1694700623
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_107
timestamp 1694700623
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_108
timestamp 1694700623
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_109
timestamp 1694700623
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_110
timestamp 1694700623
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_111
timestamp 1694700623
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_112
timestamp 1694700623
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_113
timestamp 1694700623
transform 1 0 5152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_114
timestamp 1694700623
transform 1 0 8960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_115
timestamp 1694700623
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_116
timestamp 1694700623
transform 1 0 16576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_117
timestamp 1694700623
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_118
timestamp 1694700623
transform 1 0 24192 0 1 21952
box -86 -86 310 870
<< labels >>
flabel metal3 s 25200 1792 26000 1904 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 25200 21952 26000 22064 0 FreeSans 448 0 0 0 custom_settings[10]
port 1 nsew signal input
flabel metal3 s 25200 23968 26000 24080 0 FreeSans 448 0 0 0 custom_settings[11]
port 2 nsew signal input
flabel metal3 s 25200 3808 26000 3920 0 FreeSans 448 0 0 0 custom_settings[1]
port 3 nsew signal input
flabel metal3 s 25200 5824 26000 5936 0 FreeSans 448 0 0 0 custom_settings[2]
port 4 nsew signal input
flabel metal3 s 25200 7840 26000 7952 0 FreeSans 448 0 0 0 custom_settings[3]
port 5 nsew signal input
flabel metal3 s 25200 9856 26000 9968 0 FreeSans 448 0 0 0 custom_settings[4]
port 6 nsew signal input
flabel metal3 s 25200 11872 26000 11984 0 FreeSans 448 0 0 0 custom_settings[5]
port 7 nsew signal input
flabel metal3 s 25200 13888 26000 14000 0 FreeSans 448 0 0 0 custom_settings[6]
port 8 nsew signal input
flabel metal3 s 25200 15904 26000 16016 0 FreeSans 448 0 0 0 custom_settings[7]
port 9 nsew signal input
flabel metal3 s 25200 17920 26000 18032 0 FreeSans 448 0 0 0 custom_settings[8]
port 10 nsew signal input
flabel metal3 s 25200 19936 26000 20048 0 FreeSans 448 0 0 0 custom_settings[9]
port 11 nsew signal input
flabel metal2 s 21280 25200 21392 26000 0 FreeSans 448 90 0 0 io_out
port 12 nsew signal tristate
flabel metal2 s 12768 25200 12880 26000 0 FreeSans 448 90 0 0 rst_n
port 13 nsew signal input
flabel metal4 s 4096 3076 4416 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 9920 3076 10240 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 15744 3076 16064 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 21568 3076 21888 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 7008 3076 7328 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 12832 3076 13152 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 18656 3076 18976 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 24480 3076 24800 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal2 s 4256 25200 4368 26000 0 FreeSans 448 90 0 0 wb_clk_i
port 16 nsew signal input
rlabel metal1 12992 22736 12992 22736 0 vdd
rlabel via1 13072 21952 13072 21952 0 vss
rlabel metal2 4424 13944 4424 13944 0 _000_
rlabel metal2 6664 12488 6664 12488 0 _001_
rlabel metal2 2744 12320 2744 12320 0 _002_
rlabel metal2 2464 13832 2464 13832 0 _003_
rlabel metal2 6888 9352 6888 9352 0 _004_
rlabel metal2 9912 14168 9912 14168 0 _005_
rlabel metal2 18200 8680 18200 8680 0 _006_
rlabel metal2 18536 6832 18536 6832 0 _007_
rlabel metal2 22064 6664 22064 6664 0 _008_
rlabel metal2 22120 10136 22120 10136 0 _009_
rlabel metal2 18200 14056 18200 14056 0 _010_
rlabel metal2 18200 10248 18200 10248 0 _011_
rlabel metal2 19432 13328 19432 13328 0 _012_
rlabel metal2 19544 15456 19544 15456 0 _013_
rlabel metal2 21896 18312 21896 18312 0 _014_
rlabel metal2 18200 18872 18200 18872 0 _015_
rlabel metal2 19488 19880 19488 19880 0 _016_
rlabel metal2 21336 20776 21336 20776 0 _017_
rlabel metal2 12040 12488 12040 12488 0 _018_
rlabel metal2 9352 9576 9352 9576 0 _019_
rlabel metal2 2520 10304 2520 10304 0 _020_
rlabel metal2 2520 7896 2520 7896 0 _021_
rlabel metal2 3640 6216 3640 6216 0 _022_
rlabel metal2 6888 6216 6888 6216 0 _023_
rlabel metal2 13496 6216 13496 6216 0 _024_
rlabel metal2 14952 9352 14952 9352 0 _025_
rlabel metal2 16464 19880 16464 19880 0 _026_
rlabel metal2 2968 18480 2968 18480 0 _027_
rlabel metal2 6104 13496 6104 13496 0 _028_
rlabel metal2 4984 19712 4984 19712 0 _029_
rlabel metal2 6552 14112 6552 14112 0 _030_
rlabel metal2 17416 12600 17416 12600 0 _031_
rlabel metal2 16072 7784 16072 7784 0 _032_
rlabel metal2 12600 15512 12600 15512 0 _033_
rlabel metal2 11928 16408 11928 16408 0 _034_
rlabel metal2 14056 20832 14056 20832 0 _035_
rlabel metal3 11480 19432 11480 19432 0 _036_
rlabel metal2 4760 12208 4760 12208 0 _037_
rlabel metal3 22568 16856 22568 16856 0 _038_
rlabel metal2 24136 17920 24136 17920 0 _039_
rlabel metal2 24136 11480 24136 11480 0 _040_
rlabel metal2 23184 10696 23184 10696 0 _041_
rlabel metal2 22568 16352 22568 16352 0 _042_
rlabel metal2 23464 16520 23464 16520 0 _043_
rlabel metal2 16184 18424 16184 18424 0 _044_
rlabel metal2 14616 16352 14616 16352 0 _045_
rlabel metal3 20944 15848 20944 15848 0 _046_
rlabel metal2 24024 16464 24024 16464 0 _047_
rlabel metal2 10808 18480 10808 18480 0 _048_
rlabel metal2 8792 20944 8792 20944 0 _049_
rlabel metal2 8792 18760 8792 18760 0 _050_
rlabel metal2 10136 17136 10136 17136 0 _051_
rlabel metal2 8008 20104 8008 20104 0 _052_
rlabel metal3 9296 20776 9296 20776 0 _053_
rlabel metal2 9240 20048 9240 20048 0 _054_
rlabel metal2 8456 18872 8456 18872 0 _055_
rlabel metal2 9800 18536 9800 18536 0 _056_
rlabel metal2 9856 16744 9856 16744 0 _057_
rlabel metal3 8792 16856 8792 16856 0 _058_
rlabel metal2 5320 15624 5320 15624 0 _059_
rlabel metal3 16044 17416 16044 17416 0 _060_
rlabel metal2 8680 19768 8680 19768 0 _061_
rlabel metal2 7952 14616 7952 14616 0 _062_
rlabel metal2 5936 18536 5936 18536 0 _063_
rlabel metal3 4872 17864 4872 17864 0 _064_
rlabel metal2 8680 18480 8680 18480 0 _065_
rlabel metal3 5376 18424 5376 18424 0 _066_
rlabel metal3 3080 17640 3080 17640 0 _067_
rlabel metal2 16632 18928 16632 18928 0 _068_
rlabel metal2 3640 14784 3640 14784 0 _069_
rlabel metal3 11256 18648 11256 18648 0 _070_
rlabel metal2 10248 20720 10248 20720 0 _071_
rlabel metal2 10024 20552 10024 20552 0 _072_
rlabel metal2 11256 19488 11256 19488 0 _073_
rlabel metal2 11368 18592 11368 18592 0 _074_
rlabel metal3 8736 17080 8736 17080 0 _075_
rlabel metal2 3192 16016 3192 16016 0 _076_
rlabel metal2 4088 14504 4088 14504 0 _077_
rlabel metal2 3304 16688 3304 16688 0 _078_
rlabel metal2 4984 14168 4984 14168 0 _079_
rlabel metal2 7896 15960 7896 15960 0 _080_
rlabel metal2 6328 15792 6328 15792 0 _081_
rlabel metal2 6664 16072 6664 16072 0 _082_
rlabel metal2 5208 13832 5208 13832 0 _083_
rlabel metal2 6216 13048 6216 13048 0 _084_
rlabel metal3 2520 16296 2520 16296 0 _085_
rlabel metal2 4984 13272 4984 13272 0 _086_
rlabel metal2 3080 13664 3080 13664 0 _087_
rlabel metal2 8120 14448 8120 14448 0 _088_
rlabel metal2 3080 14280 3080 14280 0 _089_
rlabel metal3 2968 14504 2968 14504 0 _090_
rlabel metal2 2240 14728 2240 14728 0 _091_
rlabel metal2 6328 15064 6328 15064 0 _092_
rlabel metal2 7336 9800 7336 9800 0 _093_
rlabel metal2 9576 13776 9576 13776 0 _094_
rlabel metal2 20552 8008 20552 8008 0 _095_
rlabel metal3 20496 15400 20496 15400 0 _096_
rlabel metal2 16296 16576 16296 16576 0 _097_
rlabel metal3 20944 18424 20944 18424 0 _098_
rlabel metal2 19152 15736 19152 15736 0 _099_
rlabel metal2 20104 7840 20104 7840 0 _100_
rlabel metal2 19376 7448 19376 7448 0 _101_
rlabel metal3 20496 18536 20496 18536 0 _102_
rlabel metal3 21560 8344 21560 8344 0 _103_
rlabel metal2 21336 7728 21336 7728 0 _104_
rlabel metal2 21336 10584 21336 10584 0 _105_
rlabel metal2 22568 10696 22568 10696 0 _106_
rlabel metal2 21896 12376 21896 12376 0 _107_
rlabel metal2 17416 18312 17416 18312 0 _108_
rlabel metal2 17640 15456 17640 15456 0 _109_
rlabel metal3 20216 12264 20216 12264 0 _110_
rlabel metal2 18480 12264 18480 12264 0 _111_
rlabel metal2 18200 14784 18200 14784 0 _112_
rlabel metal2 20272 9800 20272 9800 0 _113_
rlabel metal2 18872 9688 18872 9688 0 _114_
rlabel metal2 21336 12376 21336 12376 0 _115_
rlabel metal3 20440 11480 20440 11480 0 _116_
rlabel metal3 21504 15176 21504 15176 0 _117_
rlabel metal2 21336 16576 21336 16576 0 _118_
rlabel metal2 19992 14840 19992 14840 0 _119_
rlabel metal3 21616 16184 21616 16184 0 _120_
rlabel metal3 22008 17864 22008 17864 0 _121_
rlabel metal2 18424 18368 18424 18368 0 _122_
rlabel metal2 19320 19992 19320 19992 0 _123_
rlabel metal3 17304 18424 17304 18424 0 _124_
rlabel metal2 19880 20160 19880 20160 0 _125_
rlabel metal2 22120 20328 22120 20328 0 _126_
rlabel metal2 21560 20104 21560 20104 0 _127_
rlabel metal3 12656 8232 12656 8232 0 _128_
rlabel metal2 11368 11760 11368 11760 0 _129_
rlabel metal2 11928 11032 11928 11032 0 _130_
rlabel metal2 16184 12936 16184 12936 0 _131_
rlabel metal2 15680 12152 15680 12152 0 _132_
rlabel metal3 13104 11592 13104 11592 0 _133_
rlabel metal2 10696 10528 10696 10528 0 _134_
rlabel metal2 12824 7504 12824 7504 0 _135_
rlabel metal2 6328 7728 6328 7728 0 _136_
rlabel metal2 9688 9296 9688 9296 0 _137_
rlabel metal2 8232 7560 8232 7560 0 _138_
rlabel metal2 4536 9968 4536 9968 0 _139_
rlabel metal2 2296 10752 2296 10752 0 _140_
rlabel metal2 4424 7784 4424 7784 0 _141_
rlabel metal2 2520 7448 2520 7448 0 _142_
rlabel metal3 6888 7560 6888 7560 0 _143_
rlabel metal2 4536 6944 4536 6944 0 _144_
rlabel metal2 9800 6888 9800 6888 0 _145_
rlabel metal3 8456 6552 8456 6552 0 _146_
rlabel metal2 12600 7784 12600 7784 0 _147_
rlabel metal2 11760 6664 11760 6664 0 _148_
rlabel metal2 15064 9100 15064 9100 0 _149_
rlabel metal2 15400 11956 15400 11956 0 _150_
rlabel metal2 16520 19208 16520 19208 0 _151_
rlabel metal2 16800 19992 16800 19992 0 _152_
rlabel metal3 17136 20104 17136 20104 0 _153_
rlabel metal3 16520 12040 16520 12040 0 _154_
rlabel metal2 15848 8400 15848 8400 0 _155_
rlabel metal2 12936 14896 12936 14896 0 _156_
rlabel metal2 14728 14560 14728 14560 0 _157_
rlabel metal3 13832 15288 13832 15288 0 _158_
rlabel metal2 14168 15680 14168 15680 0 _159_
rlabel metal3 14168 19096 14168 19096 0 _160_
rlabel metal2 14336 17864 14336 17864 0 _161_
rlabel metal2 15456 18648 15456 18648 0 _162_
rlabel metal2 14392 19656 14392 19656 0 _163_
rlabel metal2 14728 18536 14728 18536 0 _164_
rlabel metal3 13664 18648 13664 18648 0 _165_
rlabel metal3 14000 19208 14000 19208 0 _166_
rlabel metal3 12600 15064 12600 15064 0 _167_
rlabel metal2 23128 5936 23128 5936 0 _168_
rlabel metal2 24136 15204 24136 15204 0 _169_
rlabel metal2 20440 16240 20440 16240 0 _170_
rlabel metal2 22456 14056 22456 14056 0 _171_
rlabel metal2 22904 16744 22904 16744 0 _172_
rlabel metal2 23128 5432 23128 5432 0 _173_
rlabel metal2 22232 12264 22232 12264 0 _174_
rlabel metal2 22904 10640 22904 10640 0 _175_
rlabel metal2 23688 11872 23688 11872 0 _176_
rlabel metal3 22232 9016 22232 9016 0 baud_delay\[0\]
rlabel metal2 22008 20160 22008 20160 0 baud_delay\[10\]
rlabel metal2 24024 21168 24024 21168 0 baud_delay\[11\]
rlabel metal2 21000 5544 21000 5544 0 baud_delay\[1\]
rlabel metal2 24248 6328 24248 6328 0 baud_delay\[2\]
rlabel metal2 21672 9240 21672 9240 0 baud_delay\[3\]
rlabel metal3 21840 12152 21840 12152 0 baud_delay\[4\]
rlabel metal2 20328 10416 20328 10416 0 baud_delay\[5\]
rlabel metal2 23464 13048 23464 13048 0 baud_delay\[6\]
rlabel metal3 22624 16072 22624 16072 0 baud_delay\[7\]
rlabel metal2 21896 17416 21896 17416 0 baud_delay\[8\]
rlabel metal2 22232 19768 22232 19768 0 baud_delay\[9\]
rlabel metal2 11536 10584 11536 10584 0 char_at\[0\]
rlabel metal3 9632 12040 9632 12040 0 char_at\[1\]
rlabel metal2 4872 10528 4872 10528 0 char_at\[2\]
rlabel metal2 6104 8372 6104 8372 0 char_at\[3\]
rlabel metal2 7560 7924 7560 7924 0 char_at\[4\]
rlabel metal3 9688 7448 9688 7448 0 char_at\[5\]
rlabel metal2 12040 8372 12040 8372 0 char_at\[6\]
rlabel metal2 8344 19264 8344 19264 0 char_pointer\[0\]
rlabel metal2 8344 21392 8344 21392 0 char_pointer\[1\]
rlabel metal2 6608 19880 6608 19880 0 char_pointer\[2\]
rlabel metal2 11032 17304 11032 17304 0 char_pointer\[3\]
rlabel metal2 17304 16744 17304 16744 0 clknet_0_wb_clk_i
rlabel metal2 2968 7140 2968 7140 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 9240 14112 9240 14112 0 clknet_2_1__leaf_wb_clk_i
rlabel via2 16856 6664 16856 6664 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 21000 17696 21000 17696 0 clknet_2_3__leaf_wb_clk_i
rlabel metal3 24626 1848 24626 1848 0 custom_settings[0]
rlabel metal2 20888 22288 20888 22288 0 custom_settings[10]
rlabel metal2 20160 22344 20160 22344 0 custom_settings[11]
rlabel metal2 24248 4088 24248 4088 0 custom_settings[1]
rlabel metal2 23352 6664 23352 6664 0 custom_settings[2]
rlabel metal2 22680 7560 22680 7560 0 custom_settings[3]
rlabel metal2 24304 7560 24304 7560 0 custom_settings[4]
rlabel metal3 21616 12824 21616 12824 0 custom_settings[5]
rlabel metal2 24248 13888 24248 13888 0 custom_settings[6]
rlabel metal3 24794 15960 24794 15960 0 custom_settings[7]
rlabel metal2 24248 18536 24248 18536 0 custom_settings[8]
rlabel metal2 22008 19488 22008 19488 0 custom_settings[9]
rlabel metal3 14616 13608 14616 13608 0 frame_counter\[0\]
rlabel metal2 14224 16968 14224 16968 0 frame_counter\[1\]
rlabel metal2 15176 18648 15176 18648 0 frame_counter\[2\]
rlabel metal2 15624 19320 15624 19320 0 frame_counter\[3\]
rlabel metal2 21336 23898 21336 23898 0 io_out
rlabel metal2 23632 3416 23632 3416 0 net1
rlabel metal2 23128 14448 23128 14448 0 net10
rlabel metal2 23800 18312 23800 18312 0 net11
rlabel metal2 22232 18928 22232 18928 0 net12
rlabel metal2 13384 19432 13384 19432 0 net13
rlabel metal2 18424 21616 18424 21616 0 net14
rlabel metal2 21112 22008 21112 22008 0 net2
rlabel metal3 21952 22120 21952 22120 0 net3
rlabel metal2 23856 5096 23856 5096 0 net4
rlabel metal2 23576 6720 23576 6720 0 net5
rlabel metal2 22960 7672 22960 7672 0 net6
rlabel metal2 23800 9128 23800 9128 0 net7
rlabel metal2 23128 12040 23128 12040 0 net8
rlabel metal2 23128 13384 23128 13384 0 net9
rlabel metal2 12768 22456 12768 22456 0 rst_n
rlabel metal2 14392 12712 14392 12712 0 uart_frame\[0\]
rlabel metal2 14168 12096 14168 12096 0 uart_frame\[1\]
rlabel metal2 11032 9856 11032 9856 0 uart_frame\[2\]
rlabel metal2 4648 10304 4648 10304 0 uart_frame\[3\]
rlabel metal3 5040 9128 5040 9128 0 uart_frame\[4\]
rlabel metal2 5880 7784 5880 7784 0 uart_frame\[5\]
rlabel metal2 9128 7224 9128 7224 0 uart_frame\[6\]
rlabel metal2 12040 7504 12040 7504 0 uart_frame\[7\]
rlabel metal2 11480 7728 11480 7728 0 uart_frame\[8\]
rlabel metal2 12824 8960 12824 8960 0 uart_frame\[9\]
rlabel metal3 6468 14280 6468 14280 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 26000 26000
<< end >>
