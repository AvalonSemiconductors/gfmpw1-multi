magic
tech gf180mcuD
magscale 1 10
timestamp 1753965954
<< metal1 >>
rect 1344 42362 44576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 44576 42362
rect 1344 42276 44576 42310
rect 5014 41970 5066 41982
rect 5014 41906 5066 41918
rect 5742 41970 5794 41982
rect 5742 41906 5794 41918
rect 8822 41970 8874 41982
rect 8822 41906 8874 41918
rect 9550 41970 9602 41982
rect 13458 41945 13470 41997
rect 13522 41945 13534 41997
rect 17266 41945 17278 41997
rect 17330 41945 17342 41997
rect 21074 41945 21086 41997
rect 21138 41945 21150 41997
rect 24882 41945 24894 41997
rect 24946 41945 24958 41997
rect 28690 41945 28702 41997
rect 28754 41945 28766 41997
rect 32498 41945 32510 41997
rect 32562 41945 32574 41997
rect 36306 41945 36318 41997
rect 36370 41945 36382 41997
rect 40114 41945 40126 41997
rect 40178 41945 40190 41997
rect 9550 41906 9602 41918
rect 14466 41806 14478 41858
rect 14530 41806 14542 41858
rect 18274 41806 18286 41858
rect 18338 41806 18350 41858
rect 22082 41806 22094 41858
rect 22146 41806 22158 41858
rect 25890 41806 25902 41858
rect 25954 41806 25966 41858
rect 29698 41806 29710 41858
rect 29762 41806 29774 41858
rect 33506 41806 33518 41858
rect 33570 41806 33582 41858
rect 37314 41806 37326 41858
rect 37378 41806 37390 41858
rect 41122 41806 41134 41858
rect 41186 41806 41198 41858
rect 6078 41746 6130 41758
rect 6078 41682 6130 41694
rect 9886 41746 9938 41758
rect 9886 41682 9938 41694
rect 1344 41578 44576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 44576 41578
rect 1344 41492 44576 41526
rect 43710 41186 43762 41198
rect 41794 41106 41806 41158
rect 41858 41106 41870 41158
rect 43710 41122 43762 41134
rect 32790 40962 32842 40974
rect 9314 40910 9326 40962
rect 9378 40959 9390 40962
rect 9874 40959 9886 40962
rect 9378 40913 9886 40959
rect 9378 40910 9390 40913
rect 9874 40910 9886 40913
rect 9938 40910 9950 40962
rect 32790 40898 32842 40910
rect 36374 40962 36426 40974
rect 36374 40898 36426 40910
rect 1344 40794 44576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 44576 40794
rect 1344 40708 44576 40742
rect 39678 40626 39730 40638
rect 39678 40562 39730 40574
rect 11790 40514 11842 40526
rect 11790 40450 11842 40462
rect 21086 40514 21138 40526
rect 21086 40450 21138 40462
rect 24558 40514 24610 40526
rect 24558 40450 24610 40462
rect 28702 40514 28754 40526
rect 28702 40450 28754 40462
rect 32398 40514 32450 40526
rect 32398 40450 32450 40462
rect 35982 40514 36034 40526
rect 35982 40450 36034 40462
rect 39006 40514 39058 40526
rect 39006 40450 39058 40462
rect 2158 40402 2210 40414
rect 2158 40338 2210 40350
rect 5462 40402 5514 40414
rect 5462 40338 5514 40350
rect 5742 40402 5794 40414
rect 5742 40338 5794 40350
rect 8430 40402 8482 40414
rect 8430 40338 8482 40350
rect 9046 40402 9098 40414
rect 9046 40338 9098 40350
rect 14478 40402 14530 40414
rect 14478 40338 14530 40350
rect 18398 40402 18450 40414
rect 18398 40338 18450 40350
rect 21870 40402 21922 40414
rect 21870 40338 21922 40350
rect 25398 40402 25450 40414
rect 25398 40338 25450 40350
rect 26014 40402 26066 40414
rect 26014 40338 26066 40350
rect 29318 40402 29370 40414
rect 29318 40338 29370 40350
rect 29710 40402 29762 40414
rect 29710 40338 29762 40350
rect 33294 40402 33346 40414
rect 39342 40402 39394 40414
rect 36362 40350 36374 40402
rect 36426 40350 36438 40402
rect 33294 40338 33346 40350
rect 39342 40338 39394 40350
rect 40406 40402 40458 40414
rect 40406 40338 40458 40350
rect 40798 40402 40850 40414
rect 40798 40338 40850 40350
rect 2930 40238 2942 40290
rect 2994 40238 3006 40290
rect 4834 40238 4846 40290
rect 4898 40238 4910 40290
rect 6514 40238 6526 40290
rect 6578 40238 6590 40290
rect 13682 40238 13694 40290
rect 13746 40238 13758 40290
rect 19170 40238 19182 40290
rect 19234 40238 19246 40290
rect 22642 40238 22654 40290
rect 22706 40238 22718 40290
rect 26786 40238 26798 40290
rect 26850 40238 26862 40290
rect 30482 40238 30494 40290
rect 30546 40238 30558 40290
rect 34066 40238 34078 40290
rect 34130 40238 34142 40290
rect 37090 40238 37102 40290
rect 37154 40238 37166 40290
rect 41570 40238 41582 40290
rect 41634 40238 41646 40290
rect 43474 40238 43486 40290
rect 43538 40238 43550 40290
rect 1344 40010 44576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 44576 40010
rect 1344 39924 44576 39958
rect 13918 39842 13970 39854
rect 13918 39778 13970 39790
rect 20190 39842 20242 39854
rect 20190 39778 20242 39790
rect 24446 39842 24498 39854
rect 23650 39734 23662 39786
rect 23714 39734 23726 39786
rect 24446 39778 24498 39790
rect 30270 39842 30322 39854
rect 30270 39778 30322 39790
rect 32846 39842 32898 39854
rect 32846 39778 32898 39790
rect 37214 39842 37266 39854
rect 37214 39778 37266 39790
rect 41022 39842 41074 39854
rect 41022 39778 41074 39790
rect 42590 39842 42642 39854
rect 42590 39778 42642 39790
rect 5058 39678 5070 39730
rect 5122 39678 5134 39730
rect 15810 39678 15822 39730
rect 15874 39678 15886 39730
rect 17714 39678 17726 39730
rect 17778 39678 17790 39730
rect 9886 39618 9938 39630
rect 13022 39618 13074 39630
rect 4610 39566 4622 39618
rect 4674 39566 4686 39618
rect 4946 39522 4958 39574
rect 5010 39522 5022 39574
rect 8997 39566 9009 39618
rect 9061 39566 9073 39618
rect 12226 39566 12238 39618
rect 12290 39566 12302 39618
rect 9886 39554 9938 39566
rect 13022 39554 13074 39566
rect 14254 39618 14306 39630
rect 14254 39554 14306 39566
rect 18510 39618 18562 39630
rect 18510 39554 18562 39566
rect 20526 39618 20578 39630
rect 24110 39618 24162 39630
rect 23538 39566 23550 39618
rect 23602 39566 23614 39618
rect 23762 39566 23774 39618
rect 23826 39566 23838 39618
rect 20526 39554 20578 39566
rect 24110 39554 24162 39566
rect 29038 39618 29090 39630
rect 29038 39554 29090 39566
rect 29262 39618 29314 39630
rect 29934 39618 29986 39630
rect 29530 39566 29542 39618
rect 29594 39566 29606 39618
rect 29262 39554 29314 39566
rect 29934 39554 29986 39566
rect 32510 39618 32562 39630
rect 32510 39554 32562 39566
rect 36878 39618 36930 39630
rect 36878 39554 36930 39566
rect 40686 39618 40738 39630
rect 40686 39554 40738 39566
rect 42926 39618 42978 39630
rect 42926 39554 42978 39566
rect 43318 39618 43370 39630
rect 43318 39554 43370 39566
rect 8766 39506 8818 39518
rect 8766 39442 8818 39454
rect 10334 39506 10386 39518
rect 10334 39442 10386 39454
rect 36150 39394 36202 39406
rect 36150 39330 36202 39342
rect 1344 39226 44576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 44576 39226
rect 1344 39140 44576 39174
rect 16046 39058 16098 39070
rect 16046 38994 16098 39006
rect 2830 38946 2882 38958
rect 2830 38882 2882 38894
rect 7758 38946 7810 38958
rect 3950 38872 4002 38884
rect 7758 38882 7810 38894
rect 2662 38834 2714 38846
rect 3042 38782 3054 38834
rect 3106 38782 3118 38834
rect 3266 38810 3278 38862
rect 3330 38810 3342 38862
rect 36392 38871 36444 38883
rect 4510 38834 4562 38846
rect 3950 38808 4002 38820
rect 4274 38782 4286 38834
rect 4338 38782 4350 38834
rect 5058 38797 5070 38849
rect 5122 38797 5134 38849
rect 8094 38834 8146 38846
rect 2662 38770 2714 38782
rect 4510 38770 4562 38782
rect 4678 38778 4730 38790
rect 5282 38782 5294 38834
rect 5346 38782 5358 38834
rect 8094 38770 8146 38782
rect 13470 38834 13522 38846
rect 13470 38770 13522 38782
rect 16382 38834 16434 38846
rect 16382 38770 16434 38782
rect 24168 38834 24220 38846
rect 24446 38834 24498 38846
rect 24322 38782 24334 38834
rect 24386 38782 24398 38834
rect 28354 38782 28366 38834
rect 28418 38782 28430 38834
rect 28690 38797 28702 38849
rect 28754 38797 28766 38849
rect 36094 38834 36146 38846
rect 36194 38782 36206 38834
rect 36258 38782 36270 38834
rect 36392 38807 36444 38819
rect 24168 38770 24220 38782
rect 24446 38770 24498 38782
rect 36094 38770 36146 38782
rect 4678 38714 4730 38726
rect 23774 38722 23826 38734
rect 35814 38722 35866 38734
rect 4946 38670 4958 38722
rect 5010 38670 5022 38722
rect 28802 38670 28814 38722
rect 28866 38670 28878 38722
rect 23774 38658 23826 38670
rect 35814 38658 35866 38670
rect 36766 38722 36818 38734
rect 36766 38658 36818 38670
rect 13806 38610 13858 38622
rect 13806 38546 13858 38558
rect 1344 38442 44576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 44576 38442
rect 1344 38356 44576 38390
rect 3950 38274 4002 38286
rect 3950 38210 4002 38222
rect 23438 38274 23490 38286
rect 23438 38210 23490 38222
rect 4622 38050 4674 38062
rect 4498 37998 4510 38050
rect 4562 37998 4574 38050
rect 4332 37942 4344 37994
rect 4396 37942 4408 37994
rect 4622 37986 4674 37998
rect 23832 38050 23884 38062
rect 24110 38050 24162 38062
rect 23986 37998 23998 38050
rect 24050 37998 24062 38050
rect 23832 37986 23884 37998
rect 24110 37986 24162 37998
rect 29038 38050 29090 38062
rect 29038 37986 29090 37998
rect 29262 38050 29314 38062
rect 29262 37986 29314 37998
rect 29822 38050 29874 38062
rect 29822 37986 29874 37998
rect 39678 38050 39730 38062
rect 40450 37998 40462 38050
rect 40514 37998 40526 38050
rect 39678 37986 39730 37998
rect 42366 37938 42418 37950
rect 29530 37886 29542 37938
rect 29594 37886 29606 37938
rect 42366 37874 42418 37886
rect 5126 37826 5178 37838
rect 30158 37826 30210 37838
rect 17490 37774 17502 37826
rect 17554 37823 17566 37826
rect 18386 37823 18398 37826
rect 17554 37777 18398 37823
rect 17554 37774 17566 37777
rect 18386 37774 18398 37777
rect 18450 37774 18462 37826
rect 5126 37762 5178 37774
rect 30158 37762 30210 37774
rect 39510 37826 39562 37838
rect 39510 37762 39562 37774
rect 1344 37658 44576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 44576 37658
rect 1344 37572 44576 37606
rect 9718 37490 9770 37502
rect 9718 37426 9770 37438
rect 21702 37490 21754 37502
rect 21702 37426 21754 37438
rect 26686 37378 26738 37390
rect 3938 37214 3950 37266
rect 4002 37214 4014 37266
rect 4678 37252 4690 37304
rect 4742 37252 4754 37304
rect 17648 37303 17700 37315
rect 5126 37266 5178 37278
rect 5126 37202 5178 37214
rect 17390 37266 17442 37278
rect 17490 37214 17502 37266
rect 17554 37214 17566 37266
rect 17648 37239 17700 37251
rect 21310 37266 21362 37278
rect 25442 37247 25454 37299
rect 25506 37247 25518 37299
rect 25890 37250 25902 37302
rect 25954 37250 25966 37302
rect 26338 37270 26350 37322
rect 26402 37270 26414 37322
rect 26686 37314 26738 37326
rect 26494 37247 26506 37299
rect 26558 37247 26570 37299
rect 27570 37214 27582 37266
rect 27634 37214 27646 37266
rect 27906 37214 27918 37266
rect 27970 37214 27982 37266
rect 41122 37214 41134 37266
rect 41186 37214 41198 37266
rect 17390 37202 17442 37214
rect 21310 37202 21362 37214
rect 18062 37154 18114 37166
rect 3838 37098 3890 37110
rect 18610 37102 18622 37154
rect 18674 37102 18686 37154
rect 20514 37102 20526 37154
rect 20578 37102 20590 37154
rect 18062 37090 18114 37102
rect 28030 37098 28082 37110
rect 3838 37034 3890 37046
rect 28030 37034 28082 37046
rect 40966 37042 41018 37054
rect 40966 36978 41018 36990
rect 1344 36874 44576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 44576 36874
rect 1344 36788 44576 36822
rect 19518 36706 19570 36718
rect 19518 36642 19570 36654
rect 25006 36594 25058 36606
rect 40126 36594 40178 36606
rect 32946 36542 32958 36594
rect 33010 36542 33022 36594
rect 25006 36530 25058 36542
rect 40126 36530 40178 36542
rect 6526 36482 6578 36494
rect 12798 36482 12850 36494
rect 7298 36430 7310 36482
rect 7362 36430 7374 36482
rect 12002 36430 12014 36482
rect 12066 36430 12078 36482
rect 6526 36418 6578 36430
rect 12798 36418 12850 36430
rect 19182 36482 19234 36494
rect 33742 36482 33794 36494
rect 40786 36486 40798 36538
rect 40850 36486 40862 36538
rect 19182 36418 19234 36430
rect 24838 36426 24890 36438
rect 25218 36430 25230 36482
rect 25282 36430 25294 36482
rect 25566 36444 25618 36456
rect 9214 36370 9266 36382
rect 9214 36306 9266 36318
rect 10110 36370 10162 36382
rect 33742 36418 33794 36430
rect 39958 36426 40010 36438
rect 25566 36380 25618 36392
rect 24838 36362 24890 36374
rect 31054 36370 31106 36382
rect 10110 36306 10162 36318
rect 40562 36374 40574 36426
rect 40626 36374 40638 36426
rect 39958 36362 40010 36374
rect 31054 36306 31106 36318
rect 18454 36258 18506 36270
rect 18454 36194 18506 36206
rect 34134 36258 34186 36270
rect 34134 36194 34186 36206
rect 37158 36258 37210 36270
rect 37158 36194 37210 36206
rect 41302 36258 41354 36270
rect 41302 36194 41354 36206
rect 1344 36090 44576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 44576 36090
rect 1344 36004 44576 36038
rect 6638 35922 6690 35934
rect 6638 35858 6690 35870
rect 11678 35922 11730 35934
rect 11678 35858 11730 35870
rect 6302 35698 6354 35710
rect 9893 35702 9905 35754
rect 9957 35702 9969 35754
rect 28960 35736 29012 35748
rect 6302 35634 6354 35646
rect 10782 35698 10834 35710
rect 10782 35634 10834 35646
rect 12014 35698 12066 35710
rect 12014 35634 12066 35646
rect 13358 35698 13410 35710
rect 14366 35698 14418 35710
rect 13906 35646 13918 35698
rect 13970 35646 13982 35698
rect 13358 35634 13410 35646
rect 14366 35634 14418 35646
rect 18398 35698 18450 35710
rect 18398 35634 18450 35646
rect 28702 35698 28754 35710
rect 28802 35646 28814 35698
rect 28866 35646 28878 35698
rect 33966 35698 34018 35710
rect 28960 35672 29012 35684
rect 29810 35646 29822 35698
rect 29874 35646 29886 35698
rect 30146 35646 30158 35698
rect 30210 35646 30222 35698
rect 28702 35634 28754 35646
rect 33966 35634 34018 35646
rect 36654 35698 36706 35710
rect 36654 35634 36706 35646
rect 37102 35698 37154 35710
rect 39118 35698 39170 35710
rect 39982 35702 39994 35754
rect 40046 35702 40058 35754
rect 37966 35646 37978 35698
rect 38030 35646 38042 35698
rect 37102 35634 37154 35646
rect 39118 35634 39170 35646
rect 41134 35698 41186 35710
rect 41134 35634 41186 35646
rect 29374 35586 29426 35598
rect 38838 35586 38890 35598
rect 34738 35534 34750 35586
rect 34802 35534 34814 35586
rect 41906 35534 41918 35586
rect 41970 35534 41982 35586
rect 43810 35534 43822 35586
rect 43874 35534 43886 35586
rect 9662 35474 9714 35486
rect 14130 35478 14142 35530
rect 14194 35478 14206 35530
rect 29374 35522 29426 35534
rect 9662 35410 9714 35422
rect 14702 35474 14754 35486
rect 14702 35410 14754 35422
rect 18734 35474 18786 35486
rect 29922 35478 29934 35530
rect 29986 35478 29998 35530
rect 38838 35522 38890 35534
rect 38222 35474 38274 35486
rect 25330 35422 25342 35474
rect 25394 35471 25406 35474
rect 26562 35471 26574 35474
rect 25394 35425 26574 35471
rect 25394 35422 25406 35425
rect 26562 35422 26574 35425
rect 26626 35422 26638 35474
rect 18734 35410 18786 35422
rect 38222 35410 38274 35422
rect 40238 35474 40290 35486
rect 40238 35410 40290 35422
rect 1344 35306 44576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 44576 35306
rect 1344 35220 44576 35254
rect 19238 35138 19290 35150
rect 19238 35074 19290 35086
rect 25230 35138 25282 35150
rect 25230 35074 25282 35086
rect 26854 35138 26906 35150
rect 26854 35074 26906 35086
rect 39174 35138 39226 35150
rect 39174 35074 39226 35086
rect 16942 35026 16994 35038
rect 37158 35026 37210 35038
rect 29250 34974 29262 35026
rect 29314 34974 29326 35026
rect 16942 34962 16994 34974
rect 37158 34962 37210 34974
rect 5854 34914 5906 34926
rect 7030 34914 7082 34926
rect 6402 34862 6414 34914
rect 6466 34862 6478 34914
rect 5854 34850 5906 34862
rect 6066 34806 6078 34858
rect 6130 34806 6142 34858
rect 7030 34850 7082 34862
rect 15262 34914 15314 34926
rect 17278 34914 17330 34926
rect 16594 34862 16606 34914
rect 16658 34862 16670 34914
rect 14142 34802 14194 34814
rect 14373 34806 14385 34858
rect 14437 34806 14449 34858
rect 15262 34850 15314 34862
rect 16930 34806 16942 34858
rect 16994 34806 17006 34858
rect 17278 34850 17330 34862
rect 17614 34914 17666 34926
rect 17614 34850 17666 34862
rect 18510 34914 18562 34926
rect 18510 34850 18562 34862
rect 18958 34914 19010 34926
rect 18666 34806 18678 34858
rect 18730 34806 18742 34858
rect 18958 34850 19010 34862
rect 24838 34914 24890 34926
rect 24838 34850 24890 34862
rect 25622 34914 25674 34926
rect 25902 34914 25954 34926
rect 27806 34914 27858 34926
rect 29822 34914 29874 34926
rect 25778 34862 25790 34914
rect 25842 34862 25854 34914
rect 26674 34862 26686 34914
rect 26738 34862 26750 34914
rect 27346 34862 27358 34914
rect 27410 34862 27422 34914
rect 28242 34862 28254 34914
rect 28306 34862 28318 34914
rect 28466 34862 28478 34914
rect 28530 34862 28542 34914
rect 29138 34862 29150 34914
rect 29202 34862 29214 34914
rect 25622 34850 25674 34862
rect 25902 34850 25954 34862
rect 27806 34850 27858 34862
rect 6290 34694 6302 34746
rect 6354 34694 6366 34746
rect 14142 34738 14194 34750
rect 18846 34802 18898 34814
rect 18846 34738 18898 34750
rect 27918 34802 27970 34814
rect 29586 34806 29598 34858
rect 29650 34806 29662 34858
rect 29822 34850 29874 34862
rect 30158 34914 30210 34926
rect 38446 34914 38498 34926
rect 36418 34862 36430 34914
rect 36482 34862 36494 34914
rect 30158 34850 30210 34862
rect 38446 34850 38498 34862
rect 38894 34914 38946 34926
rect 38602 34806 38614 34858
rect 38666 34806 38678 34858
rect 38894 34850 38946 34862
rect 39678 34914 39730 34926
rect 39678 34850 39730 34862
rect 40126 34914 40178 34926
rect 27918 34738 27970 34750
rect 38782 34802 38834 34814
rect 39834 34806 39846 34858
rect 39898 34806 39910 34858
rect 40126 34850 40178 34862
rect 40406 34914 40458 34926
rect 40406 34850 40458 34862
rect 40966 34914 41018 34926
rect 40966 34850 41018 34862
rect 41134 34914 41186 34926
rect 41346 34862 41358 34914
rect 41410 34862 41422 34914
rect 41134 34850 41186 34862
rect 41570 34834 41582 34886
rect 41634 34834 41646 34886
rect 42802 34862 42814 34914
rect 42866 34862 42878 34914
rect 38782 34738 38834 34750
rect 40014 34802 40066 34814
rect 40014 34738 40066 34750
rect 36262 34690 36314 34702
rect 36262 34626 36314 34638
rect 42646 34690 42698 34702
rect 42646 34626 42698 34638
rect 1344 34522 44576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 44576 34522
rect 1344 34436 44576 34470
rect 23662 34354 23714 34366
rect 23662 34290 23714 34302
rect 13862 34242 13914 34254
rect 17446 34242 17498 34254
rect 28354 34246 28366 34298
rect 28418 34246 28430 34298
rect 30158 34242 30210 34254
rect 13862 34178 13914 34190
rect 14310 34186 14362 34198
rect 14142 34158 14194 34170
rect 3266 34093 3278 34145
rect 3330 34093 3342 34145
rect 4734 34130 4786 34142
rect 3602 34078 3614 34130
rect 3666 34078 3678 34130
rect 4734 34066 4786 34078
rect 4958 34130 5010 34142
rect 5618 34078 5630 34130
rect 5682 34078 5694 34130
rect 5954 34093 5966 34145
rect 6018 34093 6030 34145
rect 14702 34186 14754 34198
rect 18890 34190 18902 34242
rect 18954 34190 18966 34242
rect 36094 34242 36146 34254
rect 14310 34122 14362 34134
rect 14590 34158 14642 34170
rect 14142 34094 14194 34106
rect 14702 34122 14754 34134
rect 16046 34130 16098 34142
rect 16202 34134 16214 34186
rect 16266 34134 16278 34186
rect 17446 34178 17498 34190
rect 28030 34169 28082 34181
rect 30158 34178 30210 34190
rect 30830 34186 30882 34198
rect 16494 34130 16546 34142
rect 14590 34094 14642 34106
rect 16370 34078 16382 34130
rect 16434 34078 16446 34130
rect 4958 34066 5010 34078
rect 16046 34066 16098 34078
rect 16494 34066 16546 34078
rect 16774 34130 16826 34142
rect 16774 34066 16826 34078
rect 17726 34130 17778 34142
rect 18174 34130 18226 34142
rect 17826 34078 17838 34130
rect 17890 34078 17902 34130
rect 17726 34066 17778 34078
rect 18006 34074 18058 34086
rect 15206 34018 15258 34030
rect 3154 33966 3166 34018
rect 3218 33966 3230 34018
rect 5226 33966 5238 34018
rect 5290 33966 5302 34018
rect 6066 33966 6078 34018
rect 6130 33966 6142 34018
rect 18174 34066 18226 34078
rect 18398 34130 18450 34142
rect 18398 34066 18450 34078
rect 18622 34130 18674 34142
rect 21982 34130 22034 34142
rect 23326 34130 23378 34142
rect 19394 34078 19406 34130
rect 19458 34078 19470 34130
rect 19618 34078 19630 34130
rect 19682 34078 19694 34130
rect 22306 34078 22318 34130
rect 22370 34078 22382 34130
rect 18622 34066 18674 34078
rect 21982 34066 22034 34078
rect 23326 34066 23378 34078
rect 27806 34130 27858 34142
rect 28030 34105 28082 34117
rect 28466 34078 28478 34130
rect 28530 34078 28542 34130
rect 30594 34106 30606 34158
rect 30658 34106 30670 34158
rect 36094 34178 36146 34190
rect 30830 34122 30882 34134
rect 35634 34106 35646 34158
rect 35698 34106 35710 34158
rect 27806 34066 27858 34078
rect 29990 34074 30042 34086
rect 35858 34078 35870 34130
rect 35922 34078 35934 34130
rect 18006 34010 18058 34022
rect 20246 34018 20298 34030
rect 15206 33954 15258 33966
rect 19294 33962 19346 33974
rect 20246 33954 20298 33966
rect 21254 34018 21306 34030
rect 21254 33954 21306 33966
rect 23046 34018 23098 34030
rect 23046 33954 23098 33966
rect 27302 34018 27354 34030
rect 29990 34010 30042 34022
rect 36262 34074 36314 34086
rect 36262 34010 36314 34022
rect 27302 33954 27354 33966
rect 19294 33898 19346 33910
rect 21646 33906 21698 33918
rect 21646 33842 21698 33854
rect 22486 33906 22538 33918
rect 22486 33842 22538 33854
rect 1344 33738 44576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 44576 33738
rect 1344 33652 44576 33686
rect 18846 33570 18898 33582
rect 6010 33518 6022 33570
rect 6074 33518 6086 33570
rect 6794 33518 6806 33570
rect 6858 33518 6870 33570
rect 18846 33506 18898 33518
rect 24558 33570 24610 33582
rect 24558 33506 24610 33518
rect 29374 33514 29426 33526
rect 5126 33458 5178 33470
rect 2594 33406 2606 33458
rect 2658 33406 2670 33458
rect 5126 33394 5178 33406
rect 22598 33458 22650 33470
rect 29374 33450 29426 33462
rect 22598 33394 22650 33406
rect 1822 33346 1874 33358
rect 1822 33282 1874 33294
rect 5630 33346 5682 33358
rect 5630 33282 5682 33294
rect 5742 33346 5794 33358
rect 5742 33282 5794 33294
rect 6302 33346 6354 33358
rect 6302 33282 6354 33294
rect 6526 33346 6578 33358
rect 6526 33282 6578 33294
rect 8766 33346 8818 33358
rect 8766 33282 8818 33294
rect 18174 33346 18226 33358
rect 18452 33346 18504 33358
rect 18274 33294 18286 33346
rect 18338 33294 18350 33346
rect 18174 33282 18226 33294
rect 18452 33282 18504 33294
rect 19462 33346 19514 33358
rect 19462 33282 19514 33294
rect 21646 33346 21698 33358
rect 21646 33282 21698 33294
rect 23438 33346 23490 33358
rect 23438 33282 23490 33294
rect 23662 33346 23714 33358
rect 24222 33346 24274 33358
rect 32510 33346 32562 33358
rect 23930 33294 23942 33346
rect 23994 33294 24006 33346
rect 29474 33294 29486 33346
rect 29538 33294 29550 33346
rect 29810 33294 29822 33346
rect 29874 33294 29886 33346
rect 23662 33282 23714 33294
rect 24222 33282 24274 33294
rect 32510 33282 32562 33294
rect 4510 33234 4562 33246
rect 4510 33170 4562 33182
rect 8430 33122 8482 33134
rect 8430 33058 8482 33070
rect 21982 33122 22034 33134
rect 21982 33058 22034 33070
rect 23270 33122 23322 33134
rect 23270 33058 23322 33070
rect 32846 33122 32898 33134
rect 32846 33058 32898 33070
rect 1344 32954 44576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 44576 32954
rect 1344 32868 44576 32902
rect 31278 32674 31330 32686
rect 6302 32601 6354 32613
rect 31278 32610 31330 32622
rect 36374 32674 36426 32686
rect 36374 32610 36426 32622
rect 36766 32674 36818 32686
rect 36766 32610 36818 32622
rect 41246 32674 41298 32686
rect 4622 32562 4674 32574
rect 4274 32510 4286 32562
rect 4338 32510 4350 32562
rect 4946 32510 4958 32562
rect 5010 32510 5022 32562
rect 5394 32510 5406 32562
rect 5458 32510 5470 32562
rect 5842 32510 5854 32562
rect 5906 32510 5918 32562
rect 6302 32537 6354 32549
rect 6526 32562 6578 32574
rect 4622 32498 4674 32510
rect 6526 32498 6578 32510
rect 21870 32562 21922 32574
rect 28590 32562 28642 32574
rect 36654 32562 36706 32574
rect 22642 32510 22654 32562
rect 22706 32510 22718 32562
rect 29362 32510 29374 32562
rect 29426 32510 29438 32562
rect 37102 32562 37154 32574
rect 21870 32498 21922 32510
rect 28590 32498 28642 32510
rect 36654 32498 36706 32510
rect 36934 32506 36986 32518
rect 4062 32450 4114 32462
rect 4062 32386 4114 32398
rect 6190 32450 6242 32462
rect 6190 32386 6242 32398
rect 7254 32450 7306 32462
rect 7254 32386 7306 32398
rect 16214 32450 16266 32462
rect 25398 32450 25450 32462
rect 24546 32398 24558 32450
rect 24610 32398 24622 32450
rect 16214 32386 16266 32398
rect 25398 32386 25450 32398
rect 31894 32450 31946 32462
rect 37102 32498 37154 32510
rect 37326 32562 37378 32574
rect 37326 32498 37378 32510
rect 37662 32562 37714 32574
rect 37662 32498 37714 32510
rect 40910 32562 40962 32574
rect 41066 32566 41078 32618
rect 41130 32566 41142 32618
rect 41246 32610 41298 32622
rect 40910 32498 40962 32510
rect 41358 32562 41410 32574
rect 41358 32498 41410 32510
rect 36934 32442 36986 32454
rect 31894 32386 31946 32398
rect 41638 32338 41690 32350
rect 41638 32274 41690 32286
rect 1344 32170 44576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 44576 32170
rect 1344 32084 44576 32118
rect 30494 32002 30546 32014
rect 30494 31938 30546 31950
rect 23382 31890 23434 31902
rect 16650 31838 16662 31890
rect 16714 31838 16726 31890
rect 23382 31826 23434 31838
rect 27750 31890 27802 31902
rect 27750 31826 27802 31838
rect 33462 31890 33514 31902
rect 33462 31826 33514 31838
rect 42086 31834 42138 31846
rect 7758 31778 7810 31790
rect 12574 31778 12626 31790
rect 6869 31726 6881 31778
rect 6933 31726 6945 31778
rect 11778 31726 11790 31778
rect 11842 31726 11854 31778
rect 16158 31778 16210 31790
rect 7758 31714 7810 31726
rect 12574 31714 12626 31726
rect 13794 31698 13806 31750
rect 13858 31698 13870 31750
rect 16158 31714 16210 31726
rect 16382 31778 16434 31790
rect 16382 31714 16434 31726
rect 17166 31778 17218 31790
rect 17166 31714 17218 31726
rect 22430 31778 22482 31790
rect 33630 31778 33682 31790
rect 36318 31778 36370 31790
rect 25778 31726 25790 31778
rect 25842 31726 25854 31778
rect 28354 31726 28366 31778
rect 28418 31726 28430 31778
rect 22430 31714 22482 31726
rect 29138 31698 29150 31750
rect 29202 31698 29214 31750
rect 34402 31726 34414 31778
rect 34466 31726 34478 31778
rect 36866 31726 36878 31778
rect 36930 31726 36942 31778
rect 33630 31714 33682 31726
rect 36318 31714 36370 31726
rect 41458 31698 41470 31750
rect 41522 31698 41534 31750
rect 41682 31726 41694 31778
rect 41746 31726 41758 31778
rect 42086 31770 42138 31782
rect 6638 31666 6690 31678
rect 6638 31602 6690 31614
rect 9886 31666 9938 31678
rect 9886 31602 9938 31614
rect 41918 31666 41970 31678
rect 41918 31602 41970 31614
rect 5910 31554 5962 31566
rect 5910 31490 5962 31502
rect 14814 31554 14866 31566
rect 14814 31490 14866 31502
rect 17502 31554 17554 31566
rect 17502 31490 17554 31502
rect 22766 31554 22818 31566
rect 22766 31490 22818 31502
rect 25958 31554 26010 31566
rect 25958 31490 26010 31502
rect 28198 31554 28250 31566
rect 28198 31490 28250 31502
rect 37046 31554 37098 31566
rect 40966 31554 41018 31566
rect 39330 31502 39342 31554
rect 39394 31551 39406 31554
rect 40282 31551 40294 31554
rect 39394 31505 40294 31551
rect 39394 31502 39406 31505
rect 40282 31502 40294 31505
rect 40346 31502 40358 31554
rect 37046 31490 37098 31502
rect 40966 31490 41018 31502
rect 1344 31386 44576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 44576 31386
rect 1344 31300 44576 31334
rect 32566 31218 32618 31230
rect 5618 31166 5630 31218
rect 5682 31215 5694 31218
rect 5898 31215 5910 31218
rect 5682 31169 5910 31215
rect 5682 31166 5694 31169
rect 5898 31166 5910 31169
rect 5962 31166 5974 31218
rect 32566 31154 32618 31166
rect 40294 31218 40346 31230
rect 40294 31154 40346 31166
rect 27134 31106 27186 31118
rect 9982 30980 9994 31032
rect 10046 30980 10058 31032
rect 11678 30994 11730 31006
rect 10658 30942 10670 30994
rect 10722 30942 10734 30994
rect 12226 30942 12238 30994
rect 12290 30942 12302 30994
rect 14914 30969 14926 31021
rect 14978 30969 14990 31021
rect 17950 30994 18002 31006
rect 16258 30942 16270 30994
rect 16322 30942 16334 30994
rect 16594 30942 16606 30994
rect 16658 30942 16670 30994
rect 18834 30986 18846 31038
rect 18898 30986 18910 31038
rect 26450 30998 26462 31050
rect 26514 30998 26526 31050
rect 27134 31042 27186 31054
rect 35982 31106 36034 31118
rect 28130 30998 28142 31050
rect 28194 30998 28206 31050
rect 28466 30998 28478 31050
rect 28530 30998 28542 31050
rect 35982 31042 36034 31054
rect 19170 30942 19182 30994
rect 19234 30942 19246 30994
rect 27570 30942 27582 30994
rect 27634 30942 27646 30994
rect 33058 30969 33070 31021
rect 33122 30969 33134 31021
rect 11678 30930 11730 30942
rect 17950 30930 18002 30942
rect 35814 30938 35866 30950
rect 36194 30942 36206 30994
rect 36258 30942 36270 30994
rect 36418 30970 36430 31022
rect 36482 30970 36494 31022
rect 41134 30994 41186 31006
rect 41906 30942 41918 30994
rect 41970 30942 41982 30994
rect 17558 30882 17610 30894
rect 41134 30930 41186 30942
rect 10782 30826 10834 30838
rect 16158 30826 16210 30838
rect 12450 30774 12462 30826
rect 12514 30774 12526 30826
rect 18722 30830 18734 30882
rect 18786 30830 18798 30882
rect 34066 30830 34078 30882
rect 34130 30830 34142 30882
rect 35814 30874 35866 30886
rect 43810 30830 43822 30882
rect 43874 30830 43886 30882
rect 17558 30818 17610 30830
rect 10782 30762 10834 30774
rect 16158 30762 16210 30774
rect 18286 30770 18338 30782
rect 18286 30706 18338 30718
rect 1344 30602 44576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 44576 30602
rect 1344 30516 44576 30550
rect 12126 30434 12178 30446
rect 12126 30370 12178 30382
rect 39902 30434 39954 30446
rect 39902 30370 39954 30382
rect 41974 30434 42026 30446
rect 41974 30370 42026 30382
rect 17110 30266 17162 30278
rect 19954 30270 19966 30322
rect 20018 30270 20030 30322
rect 8150 30210 8202 30222
rect 12462 30210 12514 30222
rect 8306 30158 8318 30210
rect 8370 30158 8382 30210
rect 9426 30158 9438 30210
rect 9490 30158 9502 30210
rect 8150 30146 8202 30158
rect 11666 30130 11678 30182
rect 11730 30130 11742 30182
rect 12462 30146 12514 30158
rect 12854 30210 12906 30222
rect 15598 30210 15650 30222
rect 14914 30158 14926 30210
rect 14978 30158 14990 30210
rect 16706 30158 16718 30210
rect 16770 30158 16782 30210
rect 17110 30202 17162 30214
rect 27414 30210 27466 30222
rect 12854 30146 12906 30158
rect 15362 30102 15374 30154
rect 15426 30102 15438 30154
rect 15598 30146 15650 30158
rect 16482 30102 16494 30154
rect 16546 30102 16558 30154
rect 20066 30114 20078 30166
rect 20130 30114 20142 30166
rect 20402 30158 20414 30210
rect 20466 30158 20478 30210
rect 26506 30142 26518 30194
rect 26570 30142 26582 30194
rect 27134 30182 27186 30194
rect 16942 30098 16994 30110
rect 15138 29990 15150 30042
rect 15202 29990 15214 30042
rect 16942 30034 16994 30046
rect 17558 30098 17610 30110
rect 17558 30034 17610 30046
rect 21478 30098 21530 30110
rect 26674 30102 26686 30154
rect 26738 30102 26750 30154
rect 26898 30102 26910 30154
rect 26962 30102 26974 30154
rect 27414 30146 27466 30158
rect 39230 30210 39282 30222
rect 40350 30210 40402 30222
rect 39330 30158 39342 30210
rect 39394 30158 39406 30210
rect 41214 30158 41226 30210
rect 41278 30158 41290 30210
rect 42130 30158 42142 30210
rect 42194 30158 42206 30210
rect 39230 30146 39282 30158
rect 27134 30118 27186 30130
rect 39498 30102 39510 30154
rect 39562 30102 39574 30154
rect 40350 30146 40402 30158
rect 21478 30034 21530 30046
rect 41470 30098 41522 30110
rect 41470 30034 41522 30046
rect 29250 29934 29262 29986
rect 29314 29983 29326 29986
rect 29810 29983 29822 29986
rect 29314 29937 29822 29983
rect 29314 29934 29326 29937
rect 29810 29934 29822 29937
rect 29874 29934 29886 29986
rect 1344 29818 44576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 44576 29818
rect 1344 29732 44576 29766
rect 22038 29650 22090 29662
rect 22038 29586 22090 29598
rect 3714 29389 3726 29441
rect 3778 29389 3790 29441
rect 6346 29430 6358 29482
rect 6410 29430 6422 29482
rect 6750 29426 6802 29438
rect 4050 29374 4062 29426
rect 4114 29374 4126 29426
rect 6066 29374 6078 29426
rect 6130 29374 6142 29426
rect 6750 29362 6802 29374
rect 6974 29426 7026 29438
rect 10094 29412 10106 29464
rect 10158 29412 10170 29464
rect 15542 29455 15594 29467
rect 11566 29426 11618 29438
rect 10770 29374 10782 29426
rect 10834 29374 10846 29426
rect 6974 29362 7026 29374
rect 11566 29362 11618 29374
rect 11902 29426 11954 29438
rect 15250 29374 15262 29426
rect 15314 29374 15326 29426
rect 21048 29464 21100 29476
rect 15542 29391 15594 29403
rect 20750 29426 20802 29438
rect 20850 29374 20862 29426
rect 20914 29374 20926 29426
rect 21048 29400 21100 29412
rect 26910 29426 26962 29438
rect 11902 29362 11954 29374
rect 20750 29362 20802 29374
rect 26910 29362 26962 29374
rect 33630 29426 33682 29438
rect 33630 29362 33682 29374
rect 16214 29314 16266 29326
rect 3602 29262 3614 29314
rect 3666 29262 3678 29314
rect 6514 29262 6526 29314
rect 6578 29262 6590 29314
rect 15698 29262 15710 29314
rect 15762 29262 15774 29314
rect 10546 29206 10558 29258
rect 10610 29206 10622 29258
rect 16214 29250 16266 29262
rect 20470 29314 20522 29326
rect 20470 29250 20522 29262
rect 40070 29314 40122 29326
rect 40070 29250 40122 29262
rect 21422 29202 21474 29214
rect 7242 29150 7254 29202
rect 7306 29150 7318 29202
rect 21422 29138 21474 29150
rect 27246 29202 27298 29214
rect 33294 29202 33346 29214
rect 27794 29150 27806 29202
rect 27858 29199 27870 29202
rect 29026 29199 29038 29202
rect 27858 29153 29038 29199
rect 27858 29150 27870 29153
rect 29026 29150 29038 29153
rect 29090 29150 29102 29202
rect 33954 29150 33966 29202
rect 34018 29199 34030 29202
rect 34402 29199 34414 29202
rect 34018 29153 34414 29199
rect 34018 29150 34030 29153
rect 34402 29150 34414 29153
rect 34466 29150 34478 29202
rect 27246 29138 27298 29150
rect 33294 29138 33346 29150
rect 1344 29034 44576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 44576 29034
rect 1344 28948 44576 28982
rect 20638 28866 20690 28878
rect 8206 28810 8258 28822
rect 20638 28802 20690 28814
rect 29878 28866 29930 28878
rect 2594 28702 2606 28754
rect 2658 28702 2670 28754
rect 8206 28746 8258 28758
rect 10222 28754 10274 28766
rect 25062 28754 25114 28766
rect 27234 28758 27246 28810
rect 27298 28758 27310 28810
rect 29878 28802 29930 28814
rect 34414 28866 34466 28878
rect 39218 28814 39230 28866
rect 39282 28863 39294 28866
rect 39666 28863 39678 28866
rect 39282 28817 39678 28863
rect 39282 28814 39294 28817
rect 39666 28814 39678 28817
rect 39730 28814 39742 28866
rect 34414 28802 34466 28814
rect 10994 28702 11006 28754
rect 11058 28702 11070 28754
rect 19506 28702 19518 28754
rect 19570 28702 19582 28754
rect 33282 28702 33294 28754
rect 33346 28702 33358 28754
rect 10222 28690 10274 28702
rect 25062 28690 25114 28702
rect 1822 28642 1874 28654
rect 1822 28578 1874 28590
rect 4510 28642 4562 28654
rect 4510 28578 4562 28590
rect 5126 28642 5178 28654
rect 9886 28642 9938 28654
rect 11566 28642 11618 28654
rect 20302 28642 20354 28654
rect 7746 28590 7758 28642
rect 7810 28590 7822 28642
rect 8082 28590 8094 28642
rect 8146 28590 8158 28642
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 10882 28590 10894 28642
rect 10946 28590 10958 28642
rect 19058 28590 19070 28642
rect 19122 28590 19134 28642
rect 5126 28578 5178 28590
rect 9886 28578 9938 28590
rect 10266 28534 10278 28586
rect 10330 28534 10342 28586
rect 11162 28534 11174 28586
rect 11226 28534 11238 28586
rect 11566 28578 11618 28590
rect 19394 28546 19406 28598
rect 19458 28546 19470 28598
rect 20302 28578 20354 28590
rect 21982 28642 22034 28654
rect 24670 28642 24722 28654
rect 23874 28590 23886 28642
rect 23938 28590 23950 28642
rect 21982 28578 22034 28590
rect 24670 28578 24722 28590
rect 26462 28642 26514 28654
rect 29150 28642 29202 28654
rect 27010 28590 27022 28642
rect 27074 28590 27086 28642
rect 26462 28578 26514 28590
rect 29150 28578 29202 28590
rect 29598 28642 29650 28654
rect 29306 28534 29318 28586
rect 29370 28534 29382 28586
rect 29598 28578 29650 28590
rect 31390 28642 31442 28654
rect 31390 28578 31442 28590
rect 34078 28642 34130 28654
rect 34078 28578 34130 28590
rect 34808 28642 34860 28654
rect 35086 28642 35138 28654
rect 34962 28590 34974 28642
rect 35026 28590 35038 28642
rect 34808 28578 34860 28590
rect 35086 28578 35138 28590
rect 35422 28642 35474 28654
rect 35422 28578 35474 28590
rect 35870 28642 35922 28654
rect 29486 28530 29538 28542
rect 35578 28534 35590 28586
rect 35642 28534 35654 28586
rect 35870 28578 35922 28590
rect 29486 28466 29538 28478
rect 35758 28530 35810 28542
rect 35758 28466 35810 28478
rect 36150 28530 36202 28542
rect 36150 28466 36202 28478
rect 39442 28366 39454 28418
rect 39506 28415 39518 28418
rect 40114 28415 40126 28418
rect 39506 28369 40126 28415
rect 39506 28366 39518 28369
rect 40114 28366 40126 28369
rect 40178 28366 40190 28418
rect 40674 28366 40686 28418
rect 40738 28415 40750 28418
rect 41570 28415 41582 28418
rect 40738 28369 41582 28415
rect 40738 28366 40750 28369
rect 41570 28366 41582 28369
rect 41634 28366 41646 28418
rect 1344 28250 44576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 44576 28250
rect 1344 28164 44576 28198
rect 6134 28082 6186 28094
rect 6134 28018 6186 28030
rect 18790 28082 18842 28094
rect 4622 27970 4674 27982
rect 4622 27906 4674 27918
rect 5686 27970 5738 27982
rect 10098 27974 10110 28026
rect 10162 27974 10174 28026
rect 17490 27974 17502 28026
rect 17554 27974 17566 28026
rect 18790 28018 18842 28030
rect 34246 28082 34298 28094
rect 34246 28018 34298 28030
rect 35142 28082 35194 28094
rect 35142 28018 35194 28030
rect 37102 28082 37154 28094
rect 37102 28018 37154 28030
rect 39118 28082 39170 28094
rect 39118 28018 39170 28030
rect 5686 27906 5738 27918
rect 37942 27970 37994 27982
rect 10322 27862 10334 27914
rect 10386 27862 10398 27914
rect 10670 27858 10722 27870
rect 4050 27806 4062 27858
rect 4114 27806 4126 27858
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 4834 27806 4846 27858
rect 4898 27806 4910 27858
rect 5058 27806 5070 27858
rect 5122 27806 5134 27858
rect 9986 27806 9998 27858
rect 10050 27806 10062 27858
rect 13682 27806 13694 27858
rect 13746 27806 13758 27858
rect 14018 27833 14030 27885
rect 14082 27833 14094 27885
rect 14366 27858 14418 27870
rect 10670 27794 10722 27806
rect 14366 27794 14418 27806
rect 14702 27858 14754 27870
rect 17826 27862 17838 27914
rect 17890 27862 17902 27914
rect 37942 27906 37994 27918
rect 41246 27970 41298 27982
rect 41246 27906 41298 27918
rect 18062 27858 18114 27870
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 25554 27806 25566 27858
rect 25618 27806 25630 27858
rect 25890 27833 25902 27885
rect 25954 27833 25966 27885
rect 26238 27858 26290 27870
rect 14702 27794 14754 27806
rect 18062 27794 18114 27806
rect 26238 27794 26290 27806
rect 26574 27858 26626 27870
rect 36766 27858 36818 27870
rect 28914 27806 28926 27858
rect 28978 27806 28990 27858
rect 29250 27806 29262 27858
rect 29314 27806 29326 27858
rect 29810 27806 29822 27858
rect 29874 27806 29886 27858
rect 30034 27806 30046 27858
rect 30098 27806 30110 27858
rect 26574 27794 26626 27806
rect 36766 27794 36818 27806
rect 38110 27858 38162 27870
rect 38110 27794 38162 27806
rect 38446 27858 38498 27870
rect 38446 27794 38498 27806
rect 39454 27858 39506 27870
rect 39454 27794 39506 27806
rect 40910 27858 40962 27870
rect 41358 27858 41410 27870
rect 40910 27794 40962 27806
rect 41078 27802 41130 27814
rect 24726 27746 24778 27758
rect 36598 27746 36650 27758
rect 13906 27694 13918 27746
rect 13970 27694 13982 27746
rect 25666 27694 25678 27746
rect 25730 27694 25742 27746
rect 24726 27682 24778 27694
rect 29710 27690 29762 27702
rect 29026 27638 29038 27690
rect 29090 27638 29102 27690
rect 41358 27794 41410 27806
rect 41078 27738 41130 27750
rect 36598 27682 36650 27694
rect 29710 27626 29762 27638
rect 41638 27634 41690 27646
rect 41638 27570 41690 27582
rect 1344 27466 44576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 44576 27466
rect 1344 27380 44576 27414
rect 6302 27298 6354 27310
rect 35926 27298 35978 27310
rect 6302 27234 6354 27246
rect 28142 27242 28194 27254
rect 22598 27186 22650 27198
rect 14802 27134 14814 27186
rect 14866 27134 14878 27186
rect 22598 27122 22650 27134
rect 23550 27186 23602 27198
rect 35926 27234 35978 27246
rect 37214 27298 37266 27310
rect 37214 27234 37266 27246
rect 37886 27298 37938 27310
rect 37886 27234 37938 27246
rect 39846 27298 39898 27310
rect 39846 27234 39898 27246
rect 40462 27298 40514 27310
rect 40462 27234 40514 27246
rect 28142 27178 28194 27190
rect 29934 27186 29986 27198
rect 23550 27122 23602 27134
rect 29934 27122 29986 27134
rect 39286 27130 39338 27142
rect 7422 27074 7474 27086
rect 21758 27074 21810 27086
rect 29598 27074 29650 27086
rect 35198 27074 35250 27086
rect 35646 27074 35698 27086
rect 14354 27022 14366 27074
rect 14418 27022 14430 27074
rect 6533 26966 6545 27018
rect 6597 26966 6609 27018
rect 7422 27010 7474 27022
rect 14690 26978 14702 27030
rect 14754 26978 14766 27030
rect 22990 27036 23042 27048
rect 21758 27010 21810 27022
rect 22878 27018 22930 27030
rect 15318 26962 15370 26974
rect 15318 26898 15370 26910
rect 18902 26962 18954 26974
rect 18902 26898 18954 26910
rect 21422 26962 21474 26974
rect 22990 26972 23042 26984
rect 23718 27018 23770 27030
rect 28242 27022 28254 27074
rect 28306 27022 28318 27074
rect 28578 27022 28590 27074
rect 28642 27022 28654 27074
rect 30258 27022 30270 27074
rect 30322 27022 30334 27074
rect 35522 27022 35534 27074
rect 35586 27022 35598 27074
rect 22878 26954 22930 26966
rect 29598 27010 29650 27022
rect 29922 26966 29934 27018
rect 29986 26966 29998 27018
rect 35198 27010 35250 27022
rect 35354 26966 35366 27018
rect 35418 26966 35430 27018
rect 35646 27010 35698 27022
rect 36878 27074 36930 27086
rect 36878 27010 36930 27022
rect 37550 27074 37602 27086
rect 37550 27010 37602 27022
rect 39118 27074 39170 27086
rect 41974 27130 42026 27142
rect 39286 27066 39338 27078
rect 39566 27074 39618 27086
rect 39442 27022 39454 27074
rect 39506 27022 39518 27074
rect 39118 27010 39170 27022
rect 39566 27010 39618 27022
rect 40126 27074 40178 27086
rect 41570 27022 41582 27074
rect 41634 27022 41646 27074
rect 41974 27066 42026 27078
rect 40126 27010 40178 27022
rect 23718 26954 23770 26966
rect 36486 26962 36538 26974
rect 41402 26966 41414 27018
rect 41466 26966 41478 27018
rect 21422 26898 21474 26910
rect 36486 26898 36538 26910
rect 41806 26962 41858 26974
rect 41806 26898 41858 26910
rect 34918 26850 34970 26862
rect 34918 26786 34970 26798
rect 1344 26682 44576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 44576 26682
rect 1344 26596 44576 26630
rect 22710 26514 22762 26526
rect 15362 26406 15374 26458
rect 15426 26406 15438 26458
rect 22710 26450 22762 26462
rect 36542 26514 36594 26526
rect 36542 26450 36594 26462
rect 30606 26402 30658 26414
rect 18218 26350 18230 26402
rect 18282 26350 18294 26402
rect 9534 26276 9546 26328
rect 9598 26276 9610 26328
rect 10210 26238 10222 26290
rect 10274 26238 10286 26290
rect 13570 26238 13582 26290
rect 13634 26238 13646 26290
rect 13906 26253 13918 26305
rect 13970 26253 13982 26305
rect 14590 26290 14642 26302
rect 18510 26290 18562 26302
rect 15138 26238 15150 26290
rect 15202 26238 15214 26290
rect 14590 26226 14642 26238
rect 18510 26226 18562 26238
rect 18622 26290 18674 26302
rect 18622 26226 18674 26238
rect 18958 26290 19010 26302
rect 19114 26294 19126 26346
rect 19178 26294 19190 26346
rect 30606 26338 30658 26350
rect 19406 26290 19458 26302
rect 19282 26238 19294 26290
rect 19346 26238 19358 26290
rect 22530 26238 22542 26290
rect 22594 26238 22606 26290
rect 28242 26238 28254 26290
rect 28306 26238 28318 26290
rect 28578 26265 28590 26317
rect 28642 26265 28654 26317
rect 28926 26290 28978 26302
rect 18958 26226 19010 26238
rect 19406 26226 19458 26238
rect 28926 26226 28978 26238
rect 29486 26290 29538 26302
rect 33966 26290 34018 26302
rect 30350 26238 30362 26290
rect 30414 26238 30426 26290
rect 29486 26226 29538 26238
rect 33966 26226 34018 26238
rect 36878 26290 36930 26302
rect 36878 26226 36930 26238
rect 37102 26290 37154 26302
rect 37102 26226 37154 26238
rect 40406 26290 40458 26302
rect 40406 26226 40458 26238
rect 41134 26290 41186 26302
rect 41906 26238 41918 26290
rect 41970 26238 41982 26290
rect 41134 26226 41186 26238
rect 24278 26178 24330 26190
rect 31222 26178 31274 26190
rect 10334 26122 10386 26134
rect 14018 26126 14030 26178
rect 14082 26126 14094 26178
rect 28354 26126 28366 26178
rect 28418 26126 28430 26178
rect 43810 26126 43822 26178
rect 43874 26126 43886 26178
rect 24278 26114 24330 26126
rect 31222 26114 31274 26126
rect 10334 26058 10386 26070
rect 19686 26066 19738 26078
rect 19686 26002 19738 26014
rect 34302 26066 34354 26078
rect 34302 26002 34354 26014
rect 37438 26066 37490 26078
rect 37438 26002 37490 26014
rect 1344 25898 44576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 44576 25898
rect 1344 25812 44576 25846
rect 10670 25730 10722 25742
rect 30830 25730 30882 25742
rect 18666 25678 18678 25730
rect 18730 25678 18742 25730
rect 9314 25622 9326 25674
rect 9378 25622 9390 25674
rect 10670 25666 10722 25678
rect 30830 25666 30882 25678
rect 24110 25618 24162 25630
rect 19282 25566 19294 25618
rect 19346 25566 19358 25618
rect 24110 25554 24162 25566
rect 25174 25562 25226 25574
rect 10334 25506 10386 25518
rect 9314 25454 9326 25506
rect 9378 25454 9390 25506
rect 9990 25416 10002 25468
rect 10054 25416 10066 25468
rect 10334 25442 10386 25454
rect 13806 25506 13858 25518
rect 18174 25506 18226 25518
rect 14670 25454 14682 25506
rect 14734 25454 14746 25506
rect 13806 25442 13858 25454
rect 18174 25442 18226 25454
rect 18398 25506 18450 25518
rect 19854 25506 19906 25518
rect 19170 25454 19182 25506
rect 19234 25454 19246 25506
rect 18398 25442 18450 25454
rect 14926 25394 14978 25406
rect 19618 25398 19630 25450
rect 19682 25398 19694 25450
rect 19854 25442 19906 25454
rect 22990 25506 23042 25518
rect 22990 25442 23042 25454
rect 24894 25506 24946 25518
rect 24994 25454 25006 25506
rect 25058 25454 25070 25506
rect 25174 25498 25226 25510
rect 25342 25506 25394 25518
rect 23854 25398 23866 25450
rect 23918 25398 23930 25450
rect 24894 25442 24946 25454
rect 25342 25442 25394 25454
rect 29710 25506 29762 25518
rect 30574 25454 30586 25506
rect 30638 25454 30650 25506
rect 42802 25454 42814 25506
rect 42866 25454 42878 25506
rect 29710 25442 29762 25454
rect 14926 25330 14978 25342
rect 24614 25394 24666 25406
rect 24614 25330 24666 25342
rect 25846 25394 25898 25406
rect 25846 25330 25898 25342
rect 42646 25282 42698 25294
rect 42646 25218 42698 25230
rect 1344 25114 44576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 44576 25114
rect 1344 25028 44576 25062
rect 6750 24946 6802 24958
rect 6750 24882 6802 24894
rect 15094 24946 15146 24958
rect 15094 24882 15146 24894
rect 23438 24946 23490 24958
rect 23438 24882 23490 24894
rect 13974 24778 14026 24790
rect 14590 24778 14642 24790
rect 1934 24722 1986 24734
rect 1934 24658 1986 24670
rect 4622 24722 4674 24734
rect 5954 24714 5966 24766
rect 6018 24714 6030 24766
rect 7086 24722 7138 24734
rect 6290 24670 6302 24722
rect 6354 24670 6366 24722
rect 14242 24726 14254 24778
rect 14306 24726 14318 24778
rect 14478 24750 14530 24762
rect 13974 24714 14026 24726
rect 14590 24714 14642 24726
rect 19892 24760 19944 24772
rect 14478 24686 14530 24698
rect 20190 24722 20242 24734
rect 19892 24696 19944 24708
rect 20066 24670 20078 24722
rect 20130 24670 20142 24722
rect 4622 24658 4674 24670
rect 7086 24658 7138 24670
rect 20190 24658 20242 24670
rect 22934 24722 22986 24734
rect 22934 24658 22986 24670
rect 23102 24722 23154 24734
rect 34750 24722 34802 24734
rect 23762 24670 23774 24722
rect 23826 24670 23838 24722
rect 23102 24658 23154 24670
rect 34750 24658 34802 24670
rect 5238 24610 5290 24622
rect 19518 24610 19570 24622
rect 2706 24558 2718 24610
rect 2770 24558 2782 24610
rect 5842 24558 5854 24610
rect 5906 24558 5918 24610
rect 5238 24546 5290 24558
rect 19518 24546 19570 24558
rect 13750 24498 13802 24510
rect 13750 24434 13802 24446
rect 23942 24498 23994 24510
rect 23942 24434 23994 24446
rect 34414 24498 34466 24510
rect 35802 24446 35814 24498
rect 35866 24495 35878 24498
rect 36306 24495 36318 24498
rect 35866 24449 36318 24495
rect 35866 24446 35878 24449
rect 36306 24446 36318 24449
rect 36370 24446 36382 24498
rect 34414 24434 34466 24446
rect 1344 24330 44576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 44576 24330
rect 1344 24244 44576 24278
rect 3166 24162 3218 24174
rect 3166 24098 3218 24110
rect 11902 24162 11954 24174
rect 35802 24110 35814 24162
rect 35866 24110 35878 24162
rect 11902 24098 11954 24110
rect 4902 24050 4954 24062
rect 4902 23986 4954 23998
rect 15094 24050 15146 24062
rect 15094 23986 15146 23998
rect 22934 24050 22986 24062
rect 25286 24050 25338 24062
rect 37090 24054 37102 24106
rect 37154 24054 37166 24106
rect 22934 23986 22986 23998
rect 24838 23994 24890 24006
rect 3502 23938 3554 23950
rect 3502 23874 3554 23886
rect 10110 23938 10162 23950
rect 10110 23874 10162 23886
rect 11566 23938 11618 23950
rect 11566 23874 11618 23886
rect 15262 23938 15314 23950
rect 15262 23874 15314 23886
rect 23550 23938 23602 23950
rect 23550 23874 23602 23886
rect 23774 23938 23826 23950
rect 23986 23942 23998 23994
rect 24050 23942 24062 23994
rect 25286 23986 25338 23998
rect 24838 23930 24890 23942
rect 36094 23938 36146 23950
rect 23774 23874 23826 23886
rect 24110 23900 24162 23912
rect 36094 23874 36146 23886
rect 36318 23938 36370 23950
rect 37662 23938 37714 23950
rect 40406 23938 40458 23950
rect 36978 23886 36990 23938
rect 37042 23886 37054 23938
rect 37314 23886 37326 23938
rect 37378 23886 37390 23938
rect 40002 23886 40014 23938
rect 40066 23886 40078 23938
rect 36318 23874 36370 23886
rect 37662 23874 37714 23886
rect 40406 23874 40458 23886
rect 24110 23836 24162 23848
rect 24670 23826 24722 23838
rect 23258 23774 23270 23826
rect 23322 23774 23334 23826
rect 24670 23762 24722 23774
rect 9774 23714 9826 23726
rect 9774 23650 9826 23662
rect 15598 23714 15650 23726
rect 15598 23650 15650 23662
rect 35478 23714 35530 23726
rect 35478 23650 35530 23662
rect 37998 23714 38050 23726
rect 37998 23650 38050 23662
rect 39846 23714 39898 23726
rect 39846 23650 39898 23662
rect 1344 23546 44576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 44576 23546
rect 1344 23460 44576 23494
rect 15878 23378 15930 23390
rect 3826 23270 3838 23322
rect 3890 23270 3902 23322
rect 15878 23314 15930 23326
rect 16606 23378 16658 23390
rect 16606 23314 16658 23326
rect 14702 23266 14754 23278
rect 21366 23266 21418 23278
rect 18554 23214 18566 23266
rect 18618 23214 18630 23266
rect 3950 23154 4002 23166
rect 4274 23158 4286 23210
rect 4338 23158 4350 23210
rect 5730 23158 5742 23210
rect 5794 23158 5806 23210
rect 14702 23202 14754 23214
rect 21366 23202 21418 23214
rect 30382 23266 30434 23278
rect 30382 23202 30434 23214
rect 5966 23154 6018 23166
rect 4610 23102 4622 23154
rect 4674 23102 4686 23154
rect 5394 23102 5406 23154
rect 5458 23102 5470 23154
rect 3950 23090 4002 23102
rect 5966 23090 6018 23102
rect 6302 23154 6354 23166
rect 6302 23090 6354 23102
rect 15038 23154 15090 23166
rect 16270 23154 16322 23166
rect 15474 23102 15486 23154
rect 15538 23102 15550 23154
rect 15038 23090 15090 23102
rect 16270 23090 16322 23102
rect 18062 23154 18114 23166
rect 18062 23090 18114 23102
rect 18286 23154 18338 23166
rect 21634 23129 21646 23181
rect 21698 23129 21710 23181
rect 29262 23154 29314 23166
rect 18286 23090 18338 23102
rect 30126 23102 30138 23154
rect 30190 23102 30202 23154
rect 39554 23102 39566 23154
rect 39618 23151 39630 23154
rect 39778 23151 39790 23154
rect 39618 23105 39790 23151
rect 39618 23102 39630 23105
rect 39778 23102 39790 23105
rect 39842 23102 39854 23154
rect 29262 23090 29314 23102
rect 5630 23042 5682 23054
rect 5630 22978 5682 22990
rect 36710 23042 36762 23054
rect 36710 22978 36762 22990
rect 15318 22930 15370 22942
rect 15318 22866 15370 22878
rect 22654 22930 22706 22942
rect 22654 22866 22706 22878
rect 1344 22762 44576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 44576 22762
rect 1344 22676 44576 22710
rect 28478 22594 28530 22606
rect 5674 22542 5686 22594
rect 5738 22542 5750 22594
rect 13682 22486 13694 22538
rect 13746 22486 13758 22538
rect 28478 22530 28530 22542
rect 30494 22594 30546 22606
rect 30494 22530 30546 22542
rect 31950 22594 32002 22606
rect 31950 22530 32002 22542
rect 15598 22482 15650 22494
rect 16998 22482 17050 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 8754 22430 8766 22482
rect 8818 22430 8830 22482
rect 10658 22430 10670 22482
rect 10722 22430 10734 22482
rect 16594 22430 16606 22482
rect 16658 22479 16670 22482
rect 16818 22479 16830 22482
rect 16658 22433 16830 22479
rect 16658 22430 16670 22433
rect 16818 22430 16830 22433
rect 16882 22430 16894 22482
rect 15598 22418 15650 22430
rect 16998 22418 17050 22430
rect 18958 22482 19010 22494
rect 18958 22418 19010 22430
rect 34526 22482 34578 22494
rect 34526 22418 34578 22430
rect 39622 22426 39674 22438
rect 5966 22370 6018 22382
rect 5058 22318 5070 22370
rect 5122 22318 5134 22370
rect 4778 22262 4790 22314
rect 4842 22262 4854 22314
rect 5966 22306 6018 22318
rect 6078 22370 6130 22382
rect 6078 22306 6130 22318
rect 7982 22370 8034 22382
rect 7982 22306 8034 22318
rect 11286 22370 11338 22382
rect 14926 22370 14978 22382
rect 16382 22370 16434 22382
rect 13570 22318 13582 22370
rect 13634 22318 13646 22370
rect 13906 22318 13918 22370
rect 13970 22318 13982 22370
rect 15026 22318 15038 22370
rect 15090 22318 15102 22370
rect 11286 22306 11338 22318
rect 14926 22306 14978 22318
rect 15192 22262 15204 22314
rect 15256 22262 15268 22314
rect 16382 22306 16434 22318
rect 16606 22370 16658 22382
rect 16606 22306 16658 22318
rect 17726 22370 17778 22382
rect 17726 22306 17778 22318
rect 17950 22370 18002 22382
rect 19294 22370 19346 22382
rect 18610 22318 18622 22370
rect 18674 22318 18686 22370
rect 17950 22306 18002 22318
rect 17558 22258 17610 22270
rect 18946 22262 18958 22314
rect 19010 22262 19022 22314
rect 19294 22306 19346 22318
rect 19630 22370 19682 22382
rect 19630 22306 19682 22318
rect 23774 22370 23826 22382
rect 23774 22306 23826 22318
rect 23998 22370 24050 22382
rect 23998 22306 24050 22318
rect 27358 22370 27410 22382
rect 27358 22306 27410 22318
rect 29374 22370 29426 22382
rect 33070 22370 33122 22382
rect 30238 22318 30250 22370
rect 30302 22318 30314 22370
rect 28222 22262 28234 22314
rect 28286 22262 28298 22314
rect 29374 22306 29426 22318
rect 32181 22262 32193 22314
rect 32245 22262 32257 22314
rect 33070 22306 33122 22318
rect 33406 22370 33458 22382
rect 36374 22370 36426 22382
rect 34270 22318 34282 22370
rect 34334 22318 34346 22370
rect 34850 22318 34862 22370
rect 34914 22318 34926 22370
rect 33406 22306 33458 22318
rect 35646 22314 35698 22326
rect 35970 22318 35982 22370
rect 36034 22318 36046 22370
rect 36374 22306 36426 22318
rect 39062 22370 39114 22382
rect 39062 22306 39114 22318
rect 39342 22370 39394 22382
rect 39622 22362 39674 22374
rect 39790 22370 39842 22382
rect 39342 22306 39394 22318
rect 39790 22306 39842 22318
rect 40910 22370 40962 22382
rect 41682 22318 41694 22370
rect 41746 22318 41758 22370
rect 40910 22306 40962 22318
rect 16090 22206 16102 22258
rect 16154 22206 16166 22258
rect 18218 22206 18230 22258
rect 18282 22206 18294 22258
rect 24266 22206 24278 22258
rect 24330 22206 24342 22258
rect 35646 22250 35698 22262
rect 36206 22258 36258 22270
rect 17558 22194 17610 22206
rect 35030 22202 35082 22214
rect 36206 22194 36258 22206
rect 39454 22258 39506 22270
rect 39454 22194 39506 22206
rect 43598 22258 43650 22270
rect 43598 22194 43650 22206
rect 35030 22138 35082 22150
rect 40742 22146 40794 22158
rect 40742 22082 40794 22094
rect 1344 21978 44576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 44576 21978
rect 1344 21892 44576 21926
rect 19462 21810 19514 21822
rect 19462 21746 19514 21758
rect 34190 21810 34242 21822
rect 34190 21746 34242 21758
rect 29486 21698 29538 21710
rect 12014 21642 12066 21654
rect 10005 21590 10017 21642
rect 10069 21590 10081 21642
rect 11902 21624 11954 21636
rect 10894 21586 10946 21598
rect 12014 21578 12066 21590
rect 12518 21586 12570 21598
rect 11902 21560 11954 21572
rect 10894 21522 10946 21534
rect 11174 21530 11226 21542
rect 12518 21522 12570 21534
rect 15934 21586 15986 21598
rect 15934 21522 15986 21534
rect 16158 21586 16210 21598
rect 20078 21586 20130 21598
rect 16482 21534 16494 21586
rect 16546 21534 16558 21586
rect 16818 21534 16830 21586
rect 16882 21534 16894 21586
rect 16158 21522 16210 21534
rect 20078 21522 20130 21534
rect 20302 21586 20354 21598
rect 20302 21522 20354 21534
rect 23774 21586 23826 21598
rect 28802 21590 28814 21642
rect 28866 21590 28878 21642
rect 29486 21634 29538 21646
rect 34862 21698 34914 21710
rect 34862 21634 34914 21646
rect 41246 21698 41298 21710
rect 29026 21564 29038 21616
rect 29090 21564 29102 21616
rect 34526 21586 34578 21598
rect 37550 21586 37602 21598
rect 23774 21522 23826 21534
rect 36754 21534 36766 21586
rect 36818 21534 36830 21586
rect 11174 21466 11226 21478
rect 11342 21474 11394 21486
rect 29194 21478 29206 21530
rect 29258 21478 29270 21530
rect 34526 21522 34578 21534
rect 37550 21522 37602 21534
rect 39566 21586 39618 21598
rect 40014 21586 40066 21598
rect 39566 21522 39618 21534
rect 39734 21530 39786 21542
rect 39890 21534 39902 21586
rect 39954 21534 39966 21586
rect 37942 21474 37994 21486
rect 19786 21422 19798 21474
rect 19850 21422 19862 21474
rect 40014 21522 40066 21534
rect 40910 21586 40962 21598
rect 41066 21590 41078 21642
rect 41130 21590 41142 21642
rect 41246 21634 41298 21646
rect 40910 21522 40962 21534
rect 41358 21586 41410 21598
rect 42802 21534 42814 21586
rect 42866 21534 42878 21586
rect 41358 21522 41410 21534
rect 39734 21466 39786 21478
rect 11342 21410 11394 21422
rect 9774 21362 9826 21374
rect 16594 21366 16606 21418
rect 16658 21366 16670 21418
rect 37942 21410 37994 21422
rect 23438 21362 23490 21374
rect 15642 21310 15654 21362
rect 15706 21310 15718 21362
rect 9774 21298 9826 21310
rect 23438 21298 23490 21310
rect 40294 21362 40346 21374
rect 40294 21298 40346 21310
rect 41638 21362 41690 21374
rect 41638 21298 41690 21310
rect 42646 21362 42698 21374
rect 42646 21298 42698 21310
rect 1344 21194 44576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 44576 21194
rect 1344 21108 44576 21142
rect 12014 20970 12066 20982
rect 29530 20974 29542 21026
rect 29594 20974 29606 21026
rect 5618 20862 5630 20914
rect 5682 20862 5694 20914
rect 12014 20906 12066 20918
rect 41470 20914 41522 20926
rect 13906 20862 13918 20914
rect 13970 20862 13982 20914
rect 21858 20862 21870 20914
rect 21922 20862 21934 20914
rect 23762 20862 23774 20914
rect 23826 20862 23838 20914
rect 41470 20850 41522 20862
rect 41638 20858 41690 20870
rect 24558 20802 24610 20814
rect 5730 20706 5742 20758
rect 5794 20706 5806 20758
rect 5954 20750 5966 20802
rect 6018 20750 6030 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 11890 20750 11902 20802
rect 11954 20750 11966 20802
rect 13458 20750 13470 20802
rect 13522 20750 13534 20802
rect 13738 20694 13750 20746
rect 13802 20694 13814 20746
rect 24558 20738 24610 20750
rect 29038 20802 29090 20814
rect 29038 20738 29090 20750
rect 29262 20802 29314 20814
rect 29262 20738 29314 20750
rect 40910 20746 40962 20758
rect 41234 20750 41246 20802
rect 41298 20750 41310 20802
rect 41638 20794 41690 20806
rect 40910 20682 40962 20694
rect 24950 20578 25002 20590
rect 24950 20514 25002 20526
rect 1344 20410 44576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 44576 20410
rect 1344 20324 44576 20358
rect 33126 20186 33178 20198
rect 4274 20134 4286 20186
rect 4338 20134 4350 20186
rect 11006 20130 11058 20142
rect 3502 20018 3554 20030
rect 4610 20022 4622 20074
rect 4674 20022 4686 20074
rect 11006 20066 11058 20078
rect 12630 20130 12682 20142
rect 12630 20066 12682 20078
rect 27806 20130 27858 20142
rect 33126 20122 33178 20134
rect 35366 20130 35418 20142
rect 27806 20066 27858 20078
rect 35366 20066 35418 20078
rect 35982 20130 36034 20142
rect 4846 20018 4898 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 3502 19954 3554 19966
rect 4846 19954 4898 19966
rect 5574 20018 5626 20030
rect 5574 19954 5626 19966
rect 6190 20018 6242 20030
rect 6190 19954 6242 19966
rect 6302 20018 6354 20030
rect 12126 20018 12178 20030
rect 11237 19966 11249 20018
rect 11301 19966 11313 20018
rect 6302 19954 6354 19966
rect 12126 19954 12178 19966
rect 25118 20018 25170 20030
rect 25118 19954 25170 19966
rect 28702 20018 28754 20030
rect 28702 19954 28754 19966
rect 29094 20018 29146 20030
rect 35646 20018 35698 20030
rect 35802 20022 35814 20074
rect 35866 20022 35878 20074
rect 35982 20066 36034 20078
rect 32050 19966 32062 20018
rect 32114 19966 32126 20018
rect 33282 19966 33294 20018
rect 33346 19966 33358 20018
rect 29094 19954 29146 19966
rect 35646 19954 35698 19966
rect 36094 20018 36146 20030
rect 36094 19954 36146 19966
rect 25890 19854 25902 19906
rect 25954 19854 25966 19906
rect 3166 19794 3218 19806
rect 28366 19794 28418 19806
rect 5898 19742 5910 19794
rect 5962 19742 5974 19794
rect 3166 19730 3218 19742
rect 28366 19730 28418 19742
rect 32230 19794 32282 19806
rect 32230 19730 32282 19742
rect 36374 19794 36426 19806
rect 36374 19730 36426 19742
rect 1344 19626 44576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 44576 19626
rect 1344 19540 44576 19574
rect 11006 19458 11058 19470
rect 5898 19406 5910 19458
rect 5962 19406 5974 19458
rect 11006 19394 11058 19406
rect 25902 19458 25954 19470
rect 25902 19394 25954 19406
rect 39566 19458 39618 19470
rect 39566 19394 39618 19406
rect 2594 19294 2606 19346
rect 2658 19294 2670 19346
rect 4498 19294 4510 19346
rect 4562 19294 4574 19346
rect 18162 19294 18174 19346
rect 18226 19294 18238 19346
rect 35814 19290 35866 19302
rect 1822 19234 1874 19246
rect 1822 19170 1874 19182
rect 5126 19234 5178 19246
rect 5126 19170 5178 19182
rect 6190 19234 6242 19246
rect 6190 19170 6242 19182
rect 6414 19234 6466 19246
rect 6974 19234 7026 19246
rect 6682 19182 6694 19234
rect 6746 19182 6758 19234
rect 6414 19170 6466 19182
rect 6974 19170 7026 19182
rect 7198 19234 7250 19246
rect 7198 19170 7250 19182
rect 9438 19234 9490 19246
rect 10670 19234 10722 19246
rect 9438 19170 9490 19182
rect 9762 19155 9774 19207
rect 9826 19155 9838 19207
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 10670 19170 10722 19182
rect 17782 19234 17834 19246
rect 20862 19234 20914 19246
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 17782 19170 17834 19182
rect 20862 19170 20914 19182
rect 26238 19234 26290 19246
rect 34962 19238 34974 19290
rect 35026 19238 35038 19290
rect 40742 19290 40794 19302
rect 35814 19226 35866 19238
rect 39230 19234 39282 19246
rect 26238 19170 26290 19182
rect 40742 19226 40794 19238
rect 41122 19182 41134 19234
rect 41186 19182 41198 19234
rect 35242 19126 35254 19178
rect 35306 19126 35318 19178
rect 39230 19170 39282 19182
rect 41346 19154 41358 19206
rect 41410 19154 41422 19206
rect 35646 19122 35698 19134
rect 9986 19014 9998 19066
rect 10050 19014 10062 19066
rect 35646 19058 35698 19070
rect 40910 19122 40962 19134
rect 40910 19058 40962 19070
rect 1344 18842 44576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 44576 18842
rect 1344 18756 44576 18790
rect 41190 18674 41242 18686
rect 10390 18562 10442 18574
rect 10390 18498 10442 18510
rect 15598 18562 15650 18574
rect 26562 18566 26574 18618
rect 26626 18566 26638 18618
rect 41190 18610 41242 18622
rect 15598 18498 15650 18510
rect 33406 18562 33458 18574
rect 9998 18450 10050 18462
rect 9998 18386 10050 18398
rect 14702 18450 14754 18462
rect 14702 18386 14754 18398
rect 14814 18450 14866 18462
rect 14814 18386 14866 18398
rect 15206 18450 15258 18462
rect 15206 18386 15258 18398
rect 15486 18450 15538 18462
rect 15934 18450 15986 18462
rect 16606 18450 16658 18462
rect 15486 18386 15538 18398
rect 15766 18394 15818 18406
rect 14086 18338 14138 18350
rect 16314 18398 16326 18450
rect 16378 18398 16390 18450
rect 15934 18386 15986 18398
rect 16606 18386 16658 18398
rect 16718 18450 16770 18462
rect 16718 18386 16770 18398
rect 17838 18450 17890 18462
rect 17838 18386 17890 18398
rect 19966 18450 20018 18462
rect 19966 18386 20018 18398
rect 20078 18450 20130 18462
rect 20638 18450 20690 18462
rect 26898 18454 26910 18506
rect 26962 18454 26974 18506
rect 27134 18450 27186 18462
rect 20346 18398 20358 18450
rect 20410 18398 20422 18450
rect 26450 18398 26462 18450
rect 26514 18398 26526 18450
rect 27794 18413 27806 18465
rect 27858 18413 27870 18465
rect 28758 18450 28810 18462
rect 28130 18398 28142 18450
rect 28194 18398 28206 18450
rect 20078 18386 20130 18398
rect 20638 18386 20690 18398
rect 27134 18386 27186 18398
rect 28758 18386 28810 18398
rect 28926 18450 28978 18462
rect 28926 18386 28978 18398
rect 29150 18450 29202 18462
rect 29150 18386 29202 18398
rect 30158 18450 30210 18462
rect 31022 18454 31034 18506
rect 31086 18454 31098 18506
rect 33406 18498 33458 18510
rect 30158 18386 30210 18398
rect 31278 18450 31330 18462
rect 36094 18450 36146 18462
rect 35298 18398 35310 18450
rect 35362 18398 35374 18450
rect 31278 18386 31330 18398
rect 36094 18386 36146 18398
rect 36486 18450 36538 18462
rect 36486 18386 36538 18398
rect 38670 18450 38722 18462
rect 38670 18386 38722 18398
rect 39006 18450 39058 18462
rect 39006 18386 39058 18398
rect 39118 18450 39170 18462
rect 39118 18386 39170 18398
rect 39454 18450 39506 18462
rect 41010 18398 41022 18450
rect 41074 18398 41086 18450
rect 39454 18386 39506 18398
rect 15766 18330 15818 18342
rect 21590 18338 21642 18350
rect 14086 18274 14138 18286
rect 21590 18274 21642 18286
rect 26182 18338 26234 18350
rect 27682 18286 27694 18338
rect 27746 18286 27758 18338
rect 29418 18286 29430 18338
rect 29482 18286 29494 18338
rect 26182 18274 26234 18286
rect 9662 18226 9714 18238
rect 17502 18226 17554 18238
rect 14410 18174 14422 18226
rect 14474 18174 14486 18226
rect 9662 18162 9714 18174
rect 17502 18162 17554 18174
rect 20974 18226 21026 18238
rect 20974 18162 21026 18174
rect 1344 18058 44576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 44576 18058
rect 1344 17972 44576 18006
rect 37326 17890 37378 17902
rect 21354 17838 21366 17890
rect 21418 17838 21430 17890
rect 37326 17826 37378 17838
rect 37998 17890 38050 17902
rect 38546 17838 38558 17890
rect 38610 17887 38622 17890
rect 39106 17887 39118 17890
rect 38610 17841 39118 17887
rect 38610 17838 38622 17841
rect 39106 17838 39118 17841
rect 39170 17887 39182 17890
rect 39442 17887 39454 17890
rect 39170 17841 39454 17887
rect 39170 17838 39182 17841
rect 39442 17838 39454 17841
rect 39506 17838 39518 17890
rect 37998 17826 38050 17838
rect 14198 17778 14250 17790
rect 8754 17726 8766 17778
rect 8818 17726 8830 17778
rect 10658 17726 10670 17778
rect 10722 17726 10734 17778
rect 14198 17714 14250 17726
rect 15374 17778 15426 17790
rect 15374 17714 15426 17726
rect 40742 17778 40794 17790
rect 41682 17726 41694 17778
rect 41746 17726 41758 17778
rect 43586 17726 43598 17778
rect 43650 17726 43662 17778
rect 40742 17714 40794 17726
rect 7982 17666 8034 17678
rect 7982 17602 8034 17614
rect 14702 17666 14754 17678
rect 14702 17602 14754 17614
rect 15038 17666 15090 17678
rect 17390 17666 17442 17678
rect 15698 17614 15710 17666
rect 15762 17614 15774 17666
rect 15038 17602 15090 17614
rect 15418 17558 15430 17610
rect 15482 17558 15494 17610
rect 17390 17602 17442 17614
rect 21646 17666 21698 17678
rect 21646 17602 21698 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 22262 17666 22314 17678
rect 36990 17666 37042 17678
rect 22262 17602 22314 17614
rect 33394 17586 33406 17638
rect 33458 17586 33470 17638
rect 35634 17614 35646 17666
rect 35698 17614 35710 17666
rect 36990 17602 37042 17614
rect 37662 17666 37714 17678
rect 37662 17602 37714 17614
rect 40910 17666 40962 17678
rect 40910 17602 40962 17614
rect 11286 17442 11338 17454
rect 11286 17378 11338 17390
rect 17726 17442 17778 17454
rect 17726 17378 17778 17390
rect 27414 17442 27466 17454
rect 27414 17378 27466 17390
rect 33126 17442 33178 17454
rect 33126 17378 33178 17390
rect 1344 17274 44576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 44576 17274
rect 1344 17188 44576 17222
rect 21702 17106 21754 17118
rect 21702 17042 21754 17054
rect 22206 17106 22258 17118
rect 22206 17042 22258 17054
rect 33686 17106 33738 17118
rect 33686 17042 33738 17054
rect 34190 17106 34242 17118
rect 34190 17042 34242 17054
rect 37494 16994 37546 17006
rect 14478 16882 14530 16894
rect 14478 16818 14530 16830
rect 14702 16882 14754 16894
rect 14702 16818 14754 16830
rect 20750 16882 20802 16894
rect 21018 16886 21030 16938
rect 21082 16886 21094 16938
rect 37494 16930 37546 16942
rect 21198 16882 21250 16894
rect 20850 16830 20862 16882
rect 20914 16830 20926 16882
rect 20750 16818 20802 16830
rect 21198 16818 21250 16830
rect 21870 16882 21922 16894
rect 21870 16818 21922 16830
rect 28030 16882 28082 16894
rect 28030 16818 28082 16830
rect 28366 16882 28418 16894
rect 29150 16882 29202 16894
rect 28858 16830 28870 16882
rect 28922 16830 28934 16882
rect 28366 16818 28418 16830
rect 29150 16818 29202 16830
rect 29262 16882 29314 16894
rect 29262 16818 29314 16830
rect 33854 16882 33906 16894
rect 33854 16818 33906 16830
rect 39006 16882 39058 16894
rect 39162 16886 39174 16938
rect 39226 16886 39238 16938
rect 39454 16882 39506 16894
rect 39330 16830 39342 16882
rect 39394 16830 39406 16882
rect 39006 16818 39058 16830
rect 39454 16818 39506 16830
rect 20470 16658 20522 16670
rect 14970 16606 14982 16658
rect 15034 16606 15046 16658
rect 20470 16594 20522 16606
rect 39734 16658 39786 16670
rect 39734 16594 39786 16606
rect 1344 16490 44576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 44576 16490
rect 1344 16404 44576 16438
rect 30158 16322 30210 16334
rect 30158 16258 30210 16270
rect 24950 16210 25002 16222
rect 24950 16146 25002 16158
rect 27862 16210 27914 16222
rect 27862 16146 27914 16158
rect 14926 16098 14978 16110
rect 14926 16034 14978 16046
rect 21478 16098 21530 16110
rect 21478 16034 21530 16046
rect 23046 16098 23098 16110
rect 23046 16034 23098 16046
rect 23214 16098 23266 16110
rect 23214 16034 23266 16046
rect 28142 16098 28194 16110
rect 28142 16034 28194 16046
rect 28254 16098 28306 16110
rect 39566 16098 39618 16110
rect 28254 16034 28306 16046
rect 29138 16018 29150 16070
rect 29202 16018 29214 16070
rect 39566 16034 39618 16046
rect 28522 15934 28534 15986
rect 28586 15934 28598 15986
rect 15262 15874 15314 15886
rect 15262 15810 15314 15822
rect 23550 15874 23602 15886
rect 23550 15810 23602 15822
rect 39230 15874 39282 15886
rect 39230 15810 39282 15822
rect 1344 15706 44576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 44576 15706
rect 1344 15620 44576 15654
rect 17558 15538 17610 15550
rect 17558 15474 17610 15486
rect 23886 15538 23938 15550
rect 23886 15474 23938 15486
rect 32566 15538 32618 15550
rect 32566 15474 32618 15486
rect 27806 15426 27858 15438
rect 27806 15362 27858 15374
rect 30046 15426 30098 15438
rect 4510 15314 4562 15326
rect 4510 15250 4562 15262
rect 7814 15314 7866 15326
rect 9426 15262 9438 15314
rect 9490 15262 9502 15314
rect 10322 15289 10334 15341
rect 10386 15289 10398 15341
rect 14030 15314 14082 15326
rect 23550 15314 23602 15326
rect 14802 15262 14814 15314
rect 14866 15262 14878 15314
rect 7814 15250 7866 15262
rect 14030 15250 14082 15262
rect 23550 15250 23602 15262
rect 24782 15314 24834 15326
rect 24782 15250 24834 15262
rect 25118 15314 25170 15326
rect 29710 15314 29762 15326
rect 29866 15318 29878 15370
rect 29930 15318 29942 15370
rect 30046 15362 30098 15374
rect 38334 15426 38386 15438
rect 38334 15362 38386 15374
rect 28354 15262 28366 15314
rect 28418 15262 28430 15314
rect 28578 15262 28590 15314
rect 28642 15262 28654 15314
rect 29026 15262 29038 15314
rect 29090 15262 29102 15314
rect 25118 15250 25170 15262
rect 29710 15250 29762 15262
rect 30158 15314 30210 15326
rect 30158 15250 30210 15262
rect 30438 15314 30490 15326
rect 30930 15262 30942 15314
rect 30994 15262 31006 15314
rect 31154 15306 31166 15358
rect 31218 15306 31230 15358
rect 31602 15262 31614 15314
rect 31666 15262 31678 15314
rect 31938 15277 31950 15329
rect 32002 15277 32014 15329
rect 34626 15306 34638 15358
rect 34690 15306 34702 15358
rect 39824 15351 39876 15363
rect 37998 15314 38050 15326
rect 34962 15262 34974 15314
rect 35026 15262 35038 15314
rect 30438 15250 30490 15262
rect 37998 15250 38050 15262
rect 38166 15314 38218 15326
rect 38166 15250 38218 15262
rect 38446 15314 38498 15326
rect 38446 15250 38498 15262
rect 38726 15314 38778 15326
rect 38726 15250 38778 15262
rect 39566 15314 39618 15326
rect 39666 15262 39678 15314
rect 39730 15262 39742 15314
rect 39824 15287 39876 15299
rect 39566 15250 39618 15262
rect 12966 15202 13018 15214
rect 5282 15150 5294 15202
rect 5346 15150 5358 15202
rect 7186 15150 7198 15202
rect 7250 15150 7262 15202
rect 10994 15150 11006 15202
rect 11058 15150 11070 15202
rect 12966 15138 13018 15150
rect 13862 15202 13914 15214
rect 24446 15202 24498 15214
rect 34246 15202 34298 15214
rect 16706 15150 16718 15202
rect 16770 15150 16782 15202
rect 25890 15150 25902 15202
rect 25954 15150 25966 15202
rect 31266 15150 31278 15202
rect 31330 15150 31342 15202
rect 32050 15150 32062 15202
rect 32114 15150 32126 15202
rect 34514 15150 34526 15202
rect 34578 15150 34590 15202
rect 13862 15138 13914 15150
rect 24446 15138 24498 15150
rect 28354 15094 28366 15146
rect 28418 15094 28430 15146
rect 34246 15138 34298 15150
rect 40238 15090 40290 15102
rect 41010 15038 41022 15090
rect 41074 15087 41086 15090
rect 41906 15087 41918 15090
rect 41074 15041 41918 15087
rect 41074 15038 41086 15041
rect 41906 15038 41918 15041
rect 41970 15038 41982 15090
rect 40238 15026 40290 15038
rect 1344 14922 44576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 44576 14922
rect 1344 14836 44576 14870
rect 15374 14754 15426 14766
rect 15374 14690 15426 14702
rect 40798 14754 40850 14766
rect 40798 14690 40850 14702
rect 17334 14642 17386 14654
rect 5842 14590 5854 14642
rect 5906 14590 5918 14642
rect 17334 14578 17386 14590
rect 25622 14642 25674 14654
rect 28198 14642 28250 14654
rect 27010 14590 27022 14642
rect 27074 14590 27086 14642
rect 25622 14578 25674 14590
rect 28198 14578 28250 14590
rect 29542 14642 29594 14654
rect 33126 14642 33178 14654
rect 30034 14590 30046 14642
rect 30098 14590 30110 14642
rect 31938 14590 31950 14642
rect 32002 14590 32014 14642
rect 29542 14578 29594 14590
rect 33126 14578 33178 14590
rect 40294 14642 40346 14654
rect 41906 14590 41918 14642
rect 41970 14590 41982 14642
rect 43810 14590 43822 14642
rect 43874 14590 43886 14642
rect 40294 14578 40346 14590
rect 6750 14530 6802 14542
rect 5954 14463 5966 14515
rect 6018 14463 6030 14515
rect 6290 14478 6302 14530
rect 6354 14478 6366 14530
rect 6750 14466 6802 14478
rect 7870 14530 7922 14542
rect 25230 14530 25282 14542
rect 32734 14530 32786 14542
rect 6981 14422 6993 14474
rect 7045 14422 7057 14474
rect 7870 14466 7922 14478
rect 12114 14434 12126 14486
rect 12178 14434 12190 14486
rect 12450 14478 12462 14530
rect 12514 14478 12526 14530
rect 14130 14478 14142 14530
rect 14194 14478 14206 14530
rect 14690 14450 14702 14502
rect 14754 14450 14766 14502
rect 25230 14466 25282 14478
rect 27122 14434 27134 14486
rect 27186 14434 27198 14486
rect 27458 14478 27470 14530
rect 27522 14478 27534 14530
rect 32734 14466 32786 14478
rect 33798 14530 33850 14542
rect 34750 14530 34802 14542
rect 34066 14478 34078 14530
rect 34130 14478 34142 14530
rect 33798 14466 33850 14478
rect 34402 14451 34414 14503
rect 34466 14451 34478 14503
rect 34750 14466 34802 14478
rect 38894 14530 38946 14542
rect 39342 14530 39394 14542
rect 38994 14478 39006 14530
rect 39058 14478 39070 14530
rect 38894 14466 38946 14478
rect 9942 14418 9994 14430
rect 9942 14354 9994 14366
rect 38614 14418 38666 14430
rect 39162 14422 39174 14474
rect 39226 14422 39238 14474
rect 39342 14466 39394 14478
rect 40462 14530 40514 14542
rect 40462 14466 40514 14478
rect 41134 14530 41186 14542
rect 41134 14466 41186 14478
rect 12338 14310 12350 14362
rect 12402 14310 12414 14362
rect 20358 14306 20410 14318
rect 20358 14242 20410 14254
rect 24894 14306 24946 14318
rect 34290 14310 34302 14362
rect 34354 14310 34366 14362
rect 38614 14354 38666 14366
rect 24894 14242 24946 14254
rect 1344 14138 44576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 44576 14138
rect 1344 14052 44576 14086
rect 15654 13970 15706 13982
rect 36934 13970 36986 13982
rect 7186 13918 7198 13970
rect 7250 13967 7262 13970
rect 7858 13967 7870 13970
rect 7250 13921 7870 13967
rect 7250 13918 7262 13921
rect 7858 13918 7870 13921
rect 7922 13918 7934 13970
rect 27122 13918 27134 13970
rect 27186 13967 27198 13970
rect 28354 13967 28366 13970
rect 27186 13921 28366 13967
rect 27186 13918 27198 13921
rect 28354 13918 28366 13921
rect 28418 13918 28430 13970
rect 14802 13862 14814 13914
rect 14866 13862 14878 13914
rect 15654 13906 15706 13918
rect 36934 13906 36986 13918
rect 36318 13858 36370 13870
rect 36318 13794 36370 13806
rect 10446 13746 10498 13758
rect 10446 13682 10498 13694
rect 13134 13746 13186 13758
rect 13134 13682 13186 13694
rect 13582 13746 13634 13758
rect 13862 13746 13914 13758
rect 13682 13694 13694 13746
rect 13746 13694 13758 13746
rect 14690 13694 14702 13746
rect 14754 13694 14766 13746
rect 15026 13738 15038 13790
rect 15090 13738 15102 13790
rect 19730 13738 19742 13790
rect 19794 13738 19806 13790
rect 20302 13746 20354 13758
rect 20066 13694 20078 13746
rect 20130 13694 20142 13746
rect 13582 13682 13634 13694
rect 13862 13682 13914 13694
rect 20302 13682 20354 13694
rect 20526 13746 20578 13758
rect 20526 13682 20578 13694
rect 21086 13746 21138 13758
rect 21086 13682 21138 13694
rect 21310 13746 21362 13758
rect 21310 13682 21362 13694
rect 33630 13746 33682 13758
rect 33630 13682 33682 13694
rect 11218 13582 11230 13634
rect 11282 13582 11294 13634
rect 19618 13582 19630 13634
rect 19682 13582 19694 13634
rect 34402 13582 34414 13634
rect 34466 13582 34478 13634
rect 14254 13522 14306 13534
rect 20794 13470 20806 13522
rect 20858 13470 20870 13522
rect 21578 13470 21590 13522
rect 21642 13470 21654 13522
rect 27458 13470 27470 13522
rect 27522 13519 27534 13522
rect 28130 13519 28142 13522
rect 27522 13473 28142 13519
rect 27522 13470 27534 13473
rect 28130 13470 28142 13473
rect 28194 13470 28206 13522
rect 14254 13458 14306 13470
rect 1344 13354 44576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 44576 13354
rect 1344 13268 44576 13302
rect 13526 13186 13578 13198
rect 8654 13130 8706 13142
rect 13526 13122 13578 13134
rect 34638 13186 34690 13198
rect 34638 13122 34690 13134
rect 8654 13066 8706 13078
rect 17558 13074 17610 13086
rect 40574 13074 40626 13086
rect 9426 13022 9438 13074
rect 9490 13022 9502 13074
rect 11218 13022 11230 13074
rect 11282 13022 11294 13074
rect 18498 13022 18510 13074
rect 18562 13022 18574 13074
rect 20402 13022 20414 13074
rect 20466 13022 20478 13074
rect 38210 13022 38222 13074
rect 38274 13022 38286 13074
rect 17558 13010 17610 13022
rect 40574 13010 40626 13022
rect 12238 12962 12290 12974
rect 17726 12962 17778 12974
rect 21982 12962 22034 12974
rect 7030 12906 7082 12918
rect 7410 12910 7422 12962
rect 7474 12910 7486 12962
rect 7634 12882 7646 12934
rect 7698 12882 7710 12934
rect 8194 12910 8206 12962
rect 8258 12910 8270 12962
rect 8530 12910 8542 12962
rect 8594 12910 8606 12962
rect 8978 12910 8990 12962
rect 9042 12910 9054 12962
rect 9314 12895 9326 12947
rect 9378 12895 9390 12947
rect 11330 12895 11342 12947
rect 11394 12895 11406 12947
rect 11554 12910 11566 12962
rect 11618 12910 11630 12962
rect 12238 12898 12290 12910
rect 12562 12883 12574 12935
rect 12626 12883 12638 12935
rect 12898 12910 12910 12962
rect 12962 12910 12974 12962
rect 13682 12910 13694 12962
rect 13746 12910 13758 12962
rect 21298 12910 21310 12962
rect 21362 12910 21374 12962
rect 17726 12898 17778 12910
rect 7030 12842 7082 12854
rect 7198 12850 7250 12862
rect 21746 12854 21758 12906
rect 21810 12854 21822 12906
rect 21982 12898 22034 12910
rect 34302 12962 34354 12974
rect 39902 12962 39954 12974
rect 40180 12962 40232 12974
rect 34302 12898 34354 12910
rect 38322 12866 38334 12918
rect 38386 12866 38398 12918
rect 38658 12910 38670 12962
rect 38722 12910 38734 12962
rect 40002 12910 40014 12962
rect 40066 12910 40078 12962
rect 39902 12898 39954 12910
rect 40180 12898 40232 12910
rect 7198 12786 7250 12798
rect 12574 12794 12626 12806
rect 21646 12794 21698 12806
rect 12574 12730 12626 12742
rect 14086 12738 14138 12750
rect 21646 12730 21698 12742
rect 14086 12674 14138 12686
rect 1344 12570 44576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 44576 12570
rect 1344 12484 44576 12518
rect 4958 12290 5010 12302
rect 4958 12226 5010 12238
rect 20078 12290 20130 12302
rect 20078 12226 20130 12238
rect 39156 12216 39208 12228
rect 2270 12178 2322 12190
rect 2270 12114 2322 12126
rect 5574 12178 5626 12190
rect 12562 12126 12574 12178
rect 12626 12126 12638 12178
rect 12898 12153 12910 12205
rect 12962 12153 12974 12205
rect 13246 12178 13298 12190
rect 5574 12114 5626 12126
rect 13246 12114 13298 12126
rect 13582 12178 13634 12190
rect 13582 12114 13634 12126
rect 16886 12178 16938 12190
rect 16886 12114 16938 12126
rect 17390 12178 17442 12190
rect 20626 12126 20638 12178
rect 20690 12126 20702 12178
rect 20962 12126 20974 12178
rect 21026 12126 21038 12178
rect 39454 12178 39506 12190
rect 39156 12152 39208 12164
rect 39330 12126 39342 12178
rect 39394 12126 39406 12178
rect 17390 12114 17442 12126
rect 39454 12114 39506 12126
rect 41134 12178 41186 12190
rect 41134 12114 41186 12126
rect 21478 12066 21530 12078
rect 3042 12014 3054 12066
rect 3106 12014 3118 12066
rect 12786 12014 12798 12066
rect 12850 12014 12862 12066
rect 18162 12014 18174 12066
rect 18226 12014 18238 12066
rect 20526 12010 20578 12022
rect 21478 12002 21530 12014
rect 20526 11946 20578 11958
rect 38782 11954 38834 11966
rect 38782 11890 38834 11902
rect 41470 11954 41522 11966
rect 41470 11890 41522 11902
rect 1344 11786 44576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 44576 11786
rect 1344 11700 44576 11734
rect 3726 11618 3778 11630
rect 3726 11554 3778 11566
rect 40854 11506 40906 11518
rect 19730 11454 19742 11506
rect 19794 11454 19806 11506
rect 41794 11454 41806 11506
rect 41858 11454 41870 11506
rect 43698 11454 43710 11506
rect 43762 11454 43774 11506
rect 40854 11442 40906 11454
rect 4062 11394 4114 11406
rect 7422 11394 7474 11406
rect 27918 11394 27970 11406
rect 6738 11342 6750 11394
rect 6802 11342 6814 11394
rect 7198 11355 7250 11367
rect 4062 11330 4114 11342
rect 7422 11330 7474 11342
rect 19842 11327 19854 11379
rect 19906 11327 19918 11379
rect 20178 11342 20190 11394
rect 20242 11342 20254 11394
rect 27918 11330 27970 11342
rect 38894 11394 38946 11406
rect 38894 11330 38946 11342
rect 41022 11394 41074 11406
rect 41022 11330 41074 11342
rect 7198 11291 7250 11303
rect 6850 11174 6862 11226
rect 6914 11174 6926 11226
rect 28254 11170 28306 11182
rect 28254 11106 28306 11118
rect 38558 11170 38610 11182
rect 38558 11106 38610 11118
rect 1344 11002 44576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 44576 11002
rect 1344 10916 44576 10950
rect 12966 10834 13018 10846
rect 26518 10834 26570 10846
rect 12966 10770 13018 10782
rect 24614 10778 24666 10790
rect 26518 10770 26570 10782
rect 36710 10834 36762 10846
rect 36710 10770 36762 10782
rect 22474 10670 22486 10722
rect 22538 10670 22550 10722
rect 24614 10714 24666 10726
rect 39566 10722 39618 10734
rect 25756 10648 25808 10660
rect 39566 10658 39618 10670
rect 9998 10610 10050 10622
rect 9998 10546 10050 10558
rect 12686 10610 12738 10622
rect 21982 10610 22034 10622
rect 13122 10558 13134 10610
rect 13186 10558 13198 10610
rect 12686 10546 12738 10558
rect 21982 10546 22034 10558
rect 22206 10610 22258 10622
rect 24434 10558 24446 10610
rect 24498 10558 24510 10610
rect 26014 10610 26066 10622
rect 25756 10584 25808 10596
rect 25890 10558 25902 10610
rect 25954 10558 25966 10610
rect 22206 10546 22258 10558
rect 26014 10546 26066 10558
rect 27470 10610 27522 10622
rect 30606 10610 30658 10622
rect 32958 10610 33010 10622
rect 28242 10558 28254 10610
rect 28306 10558 28318 10610
rect 31470 10558 31482 10610
rect 31534 10558 31546 10610
rect 27470 10546 27522 10558
rect 30606 10546 30658 10558
rect 32958 10546 33010 10558
rect 33182 10610 33234 10622
rect 33182 10546 33234 10558
rect 36878 10610 36930 10622
rect 37650 10558 37662 10610
rect 37714 10558 37726 10610
rect 36878 10546 36930 10558
rect 10390 10498 10442 10510
rect 30146 10446 30158 10498
rect 30210 10446 30222 10498
rect 10390 10434 10442 10446
rect 9662 10386 9714 10398
rect 9662 10322 9714 10334
rect 12350 10386 12402 10398
rect 12350 10322 12402 10334
rect 25342 10386 25394 10398
rect 25342 10322 25394 10334
rect 31726 10386 31778 10398
rect 33450 10334 33462 10386
rect 33514 10334 33526 10386
rect 31726 10322 31778 10334
rect 1344 10218 44576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 44576 10218
rect 1344 10132 44576 10166
rect 28074 9998 28086 10050
rect 28138 9998 28150 10050
rect 32554 9998 32566 10050
rect 32618 9998 32630 10050
rect 5798 9938 5850 9950
rect 11510 9938 11562 9950
rect 30550 9938 30602 9950
rect 4946 9886 4958 9938
rect 5010 9886 5022 9938
rect 7858 9886 7870 9938
rect 7922 9886 7934 9938
rect 23762 9886 23774 9938
rect 23826 9886 23838 9938
rect 27122 9886 27134 9938
rect 27186 9886 27198 9938
rect 5798 9874 5850 9886
rect 11510 9874 11562 9886
rect 30550 9874 30602 9886
rect 37158 9938 37210 9950
rect 37158 9874 37210 9886
rect 2270 9826 2322 9838
rect 7086 9826 7138 9838
rect 3042 9774 3054 9826
rect 3106 9774 3118 9826
rect 2270 9762 2322 9774
rect 7086 9762 7138 9774
rect 7422 9826 7474 9838
rect 8990 9826 9042 9838
rect 7422 9762 7474 9774
rect 7970 9759 7982 9811
rect 8034 9759 8046 9811
rect 8194 9774 8206 9826
rect 8258 9774 8270 9826
rect 8990 9762 9042 9774
rect 9102 9826 9154 9838
rect 26462 9826 26514 9838
rect 27582 9826 27634 9838
rect 25666 9774 25678 9826
rect 25730 9774 25742 9826
rect 26674 9774 26686 9826
rect 26738 9774 26750 9826
rect 9102 9762 9154 9774
rect 26462 9762 26514 9774
rect 27010 9759 27022 9811
rect 27074 9759 27086 9811
rect 27582 9762 27634 9774
rect 27806 9826 27858 9838
rect 31614 9826 31666 9838
rect 30930 9774 30942 9826
rect 30994 9774 31006 9826
rect 27806 9762 27858 9774
rect 31378 9718 31390 9770
rect 31442 9718 31454 9770
rect 31614 9762 31666 9774
rect 32062 9826 32114 9838
rect 32062 9762 32114 9774
rect 32286 9826 32338 9838
rect 36206 9826 36258 9838
rect 35410 9774 35422 9826
rect 35474 9774 35486 9826
rect 32286 9762 32338 9774
rect 36206 9762 36258 9774
rect 33518 9714 33570 9726
rect 8698 9662 8710 9714
rect 8762 9662 8774 9714
rect 31714 9606 31726 9658
rect 31778 9606 31790 9658
rect 33518 9650 33570 9662
rect 1344 9434 44576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 44576 9434
rect 1344 9348 44576 9382
rect 4174 9266 4226 9278
rect 4174 9202 4226 9214
rect 27414 9266 27466 9278
rect 7298 9158 7310 9210
rect 7362 9158 7374 9210
rect 10782 9154 10834 9166
rect 4510 9042 4562 9054
rect 7634 9046 7646 9098
rect 7698 9046 7710 9098
rect 10782 9090 10834 9102
rect 13470 9154 13522 9166
rect 25554 9158 25566 9210
rect 25618 9158 25630 9210
rect 27414 9202 27466 9214
rect 34078 9266 34130 9278
rect 34078 9202 34130 9214
rect 33114 9102 33126 9154
rect 33178 9102 33190 9154
rect 7870 9042 7922 9054
rect 7186 8990 7198 9042
rect 7250 8990 7262 9042
rect 9762 9034 9774 9086
rect 9826 9034 9838 9086
rect 10446 9042 10498 9054
rect 10098 8990 10110 9042
rect 10162 8990 10174 9042
rect 4510 8978 4562 8990
rect 7870 8978 7922 8990
rect 10446 8978 10498 8990
rect 10614 9042 10666 9054
rect 10614 8978 10666 8990
rect 10894 9042 10946 9054
rect 10894 8978 10946 8990
rect 11790 9042 11842 9054
rect 11790 8978 11842 8990
rect 12126 9042 12178 9054
rect 12338 9046 12350 9098
rect 12402 9046 12414 9098
rect 13134 9042 13186 9054
rect 13290 9046 13302 9098
rect 13354 9046 13366 9098
rect 13470 9090 13522 9102
rect 12786 8990 12798 9042
rect 12850 8990 12862 9042
rect 12126 8978 12178 8990
rect 13134 8978 13186 8990
rect 13582 9042 13634 9054
rect 19730 8990 19742 9042
rect 19794 8990 19806 9042
rect 19954 9034 19966 9086
rect 20018 9034 20030 9086
rect 25386 9046 25398 9098
rect 25450 9046 25462 9098
rect 33406 9042 33458 9054
rect 25666 8990 25678 9042
rect 25730 8990 25742 9042
rect 32162 8990 32174 9042
rect 32226 8990 32238 9042
rect 32386 8990 32398 9042
rect 32450 8990 32462 9042
rect 13582 8978 13634 8990
rect 33406 8978 33458 8990
rect 33518 9042 33570 9054
rect 33518 8978 33570 8990
rect 33742 9042 33794 9054
rect 33742 8978 33794 8990
rect 20806 8930 20858 8942
rect 9650 8878 9662 8930
rect 9714 8878 9726 8930
rect 12562 8878 12574 8930
rect 12626 8878 12638 8930
rect 20066 8878 20078 8930
rect 20130 8878 20142 8930
rect 20806 8866 20858 8878
rect 26630 8930 26682 8942
rect 26630 8866 26682 8878
rect 11174 8818 11226 8830
rect 11174 8754 11226 8766
rect 13862 8818 13914 8830
rect 32274 8822 32286 8874
rect 32338 8822 32350 8874
rect 13862 8754 13914 8766
rect 1344 8650 44576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 44576 8650
rect 1344 8564 44576 8598
rect 7522 8430 7534 8482
rect 7586 8479 7598 8482
rect 8194 8479 8206 8482
rect 7586 8433 8206 8479
rect 7586 8430 7598 8433
rect 8194 8430 8206 8433
rect 8258 8430 8270 8482
rect 16326 8370 16378 8382
rect 21646 8370 21698 8382
rect 19170 8318 19182 8370
rect 19234 8318 19246 8370
rect 16326 8306 16378 8318
rect 21646 8306 21698 8318
rect 13470 8258 13522 8270
rect 14758 8258 14810 8270
rect 10658 8206 10670 8258
rect 10722 8206 10734 8258
rect 10994 8191 11006 8243
rect 11058 8191 11070 8243
rect 14130 8206 14142 8258
rect 14194 8206 14206 8258
rect 13470 8194 13522 8206
rect 14758 8194 14810 8206
rect 16494 8258 16546 8270
rect 20302 8258 20354 8270
rect 21982 8258 22034 8270
rect 17266 8206 17278 8258
rect 17330 8206 17342 8258
rect 19730 8206 19742 8258
rect 19794 8206 19806 8258
rect 20078 8219 20130 8231
rect 16494 8194 16546 8206
rect 21298 8206 21310 8258
rect 21362 8206 21374 8258
rect 21758 8219 21810 8231
rect 20302 8194 20354 8206
rect 20078 8155 20130 8167
rect 21982 8194 22034 8206
rect 22318 8258 22370 8270
rect 22318 8194 22370 8206
rect 24222 8258 24274 8270
rect 24222 8194 24274 8206
rect 24446 8258 24498 8270
rect 24446 8194 24498 8206
rect 21758 8155 21810 8167
rect 23930 8094 23942 8146
rect 23994 8094 24006 8146
rect 10882 8038 10894 8090
rect 10946 8038 10958 8090
rect 14242 8038 14254 8090
rect 14306 8038 14318 8090
rect 19730 8038 19742 8090
rect 19794 8038 19806 8090
rect 1344 7866 44576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 44576 7866
rect 1344 7780 44576 7814
rect 18062 7698 18114 7710
rect 18062 7634 18114 7646
rect 20570 7534 20582 7586
rect 20634 7534 20646 7586
rect 22138 7534 22150 7586
rect 22202 7534 22214 7586
rect 14142 7474 14194 7486
rect 14142 7410 14194 7422
rect 14366 7474 14418 7486
rect 14366 7410 14418 7422
rect 18398 7474 18450 7486
rect 18398 7410 18450 7422
rect 20190 7474 20242 7486
rect 20190 7410 20242 7422
rect 20302 7474 20354 7486
rect 20302 7410 20354 7422
rect 21646 7474 21698 7486
rect 21646 7410 21698 7422
rect 21870 7474 21922 7486
rect 21870 7410 21922 7422
rect 14634 7198 14646 7250
rect 14698 7198 14710 7250
rect 1344 7082 44576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 44576 7082
rect 1344 6996 44576 7030
rect 21858 6862 21870 6914
rect 21922 6911 21934 6914
rect 22418 6911 22430 6914
rect 21922 6865 22430 6911
rect 21922 6862 21934 6865
rect 22418 6862 22430 6865
rect 22482 6862 22494 6914
rect 8374 6746 8426 6758
rect 7646 6652 7698 6664
rect 7970 6638 7982 6690
rect 8034 6638 8046 6690
rect 8374 6682 8426 6694
rect 12686 6690 12738 6702
rect 12686 6626 12738 6638
rect 13022 6690 13074 6702
rect 30830 6690 30882 6702
rect 14130 6638 14142 6690
rect 14194 6687 14206 6690
rect 14634 6687 14646 6690
rect 14194 6641 14646 6687
rect 14194 6638 14206 6641
rect 14634 6638 14646 6641
rect 14698 6638 14710 6690
rect 13022 6626 13074 6638
rect 30830 6626 30882 6638
rect 30942 6690 30994 6702
rect 31502 6690 31554 6702
rect 31210 6638 31222 6690
rect 31274 6638 31286 6690
rect 30942 6626 30994 6638
rect 31502 6626 31554 6638
rect 31726 6690 31778 6702
rect 31994 6638 32006 6690
rect 32058 6638 32070 6690
rect 31726 6626 31778 6638
rect 7646 6588 7698 6600
rect 8206 6578 8258 6590
rect 8206 6514 8258 6526
rect 20358 6466 20410 6478
rect 20358 6402 20410 6414
rect 1344 6298 44576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 44576 6298
rect 1344 6212 44576 6246
rect 27190 6130 27242 6142
rect 12114 6022 12126 6074
rect 12178 6022 12190 6074
rect 27190 6066 27242 6078
rect 30774 6130 30826 6142
rect 28466 6022 28478 6074
rect 28530 6022 28542 6074
rect 30774 6066 30826 6078
rect 31826 6022 31838 6074
rect 31890 6022 31902 6074
rect 12462 5945 12514 5957
rect 7758 5906 7810 5918
rect 7758 5842 7810 5854
rect 7870 5906 7922 5918
rect 8430 5906 8482 5918
rect 8138 5854 8150 5906
rect 8202 5854 8214 5906
rect 7870 5842 7922 5854
rect 8430 5842 8482 5854
rect 8654 5906 8706 5918
rect 9762 5854 9774 5906
rect 9826 5854 9838 5906
rect 12002 5854 12014 5906
rect 12066 5854 12078 5906
rect 12462 5881 12514 5893
rect 12686 5906 12738 5918
rect 8654 5842 8706 5854
rect 12686 5842 12738 5854
rect 14142 5906 14194 5918
rect 20750 5906 20802 5918
rect 19730 5854 19742 5906
rect 19794 5854 19806 5906
rect 19954 5854 19966 5906
rect 20018 5854 20030 5906
rect 20458 5854 20470 5906
rect 20522 5854 20534 5906
rect 14142 5842 14194 5854
rect 20750 5842 20802 5854
rect 20862 5906 20914 5918
rect 20862 5842 20914 5854
rect 21086 5906 21138 5918
rect 21086 5842 21138 5854
rect 21310 5906 21362 5918
rect 21310 5842 21362 5854
rect 22430 5906 22482 5918
rect 22430 5842 22482 5854
rect 22542 5906 22594 5918
rect 23550 5906 23602 5918
rect 22810 5854 22822 5906
rect 22874 5854 22886 5906
rect 22542 5842 22594 5854
rect 23550 5842 23602 5854
rect 23774 5906 23826 5918
rect 27570 5898 27582 5950
rect 27634 5898 27646 5950
rect 31502 5945 31554 5957
rect 27906 5854 27918 5906
rect 27970 5854 27982 5906
rect 28242 5854 28254 5906
rect 28306 5854 28318 5906
rect 28578 5881 28590 5933
rect 28642 5881 28654 5933
rect 28926 5906 28978 5918
rect 23774 5842 23826 5854
rect 28926 5842 28978 5854
rect 29486 5906 29538 5918
rect 29486 5842 29538 5854
rect 29598 5906 29650 5918
rect 31042 5854 31054 5906
rect 31106 5854 31118 5906
rect 31502 5881 31554 5893
rect 31726 5906 31778 5918
rect 29598 5842 29650 5854
rect 31726 5842 31778 5854
rect 32958 5906 33010 5918
rect 32958 5842 33010 5854
rect 9606 5738 9658 5750
rect 20078 5738 20130 5750
rect 27458 5742 27470 5794
rect 27522 5742 27534 5794
rect 29866 5742 29878 5794
rect 29930 5742 29942 5794
rect 8922 5630 8934 5682
rect 8986 5630 8998 5682
rect 9606 5674 9658 5686
rect 13806 5682 13858 5694
rect 20078 5674 20130 5686
rect 33294 5682 33346 5694
rect 21578 5630 21590 5682
rect 21642 5630 21654 5682
rect 24042 5630 24054 5682
rect 24106 5630 24118 5682
rect 13806 5618 13858 5630
rect 33294 5618 33346 5630
rect 1344 5514 44576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 44576 5514
rect 1344 5428 44576 5462
rect 9830 5234 9882 5246
rect 13638 5234 13690 5246
rect 17446 5234 17498 5246
rect 35254 5234 35306 5246
rect 9202 5182 9214 5234
rect 9266 5182 9278 5234
rect 10882 5182 10894 5234
rect 10946 5182 10958 5234
rect 12786 5182 12798 5234
rect 12850 5182 12862 5234
rect 14018 5182 14030 5234
rect 14082 5182 14094 5234
rect 15922 5182 15934 5234
rect 15986 5182 15998 5234
rect 20290 5182 20302 5234
rect 20354 5182 20366 5234
rect 23202 5182 23214 5234
rect 23266 5182 23278 5234
rect 31602 5182 31614 5234
rect 31666 5182 31678 5234
rect 34066 5182 34078 5234
rect 34130 5182 34142 5234
rect 9830 5170 9882 5182
rect 13638 5170 13690 5182
rect 17446 5170 17498 5182
rect 35254 5170 35306 5182
rect 6526 5122 6578 5134
rect 10110 5122 10162 5134
rect 7298 5070 7310 5122
rect 7362 5070 7374 5122
rect 6526 5058 6578 5070
rect 10110 5058 10162 5070
rect 16718 5122 16770 5134
rect 16718 5058 16770 5070
rect 17614 5122 17666 5134
rect 25902 5122 25954 5134
rect 18386 5070 18398 5122
rect 18450 5070 18462 5122
rect 25106 5070 25118 5122
rect 25170 5070 25182 5122
rect 17614 5058 17666 5070
rect 25902 5058 25954 5070
rect 26294 5122 26346 5134
rect 26294 5058 26346 5070
rect 28478 5122 28530 5134
rect 32174 5122 32226 5134
rect 31266 5070 31278 5122
rect 31330 5070 31342 5122
rect 31558 5092 31610 5104
rect 28478 5058 28530 5070
rect 32174 5058 32226 5070
rect 34862 5122 34914 5134
rect 34862 5058 34914 5070
rect 31558 5028 31610 5040
rect 28142 4898 28194 4910
rect 28142 4834 28194 4846
rect 1344 4730 44576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 44576 4730
rect 1344 4644 44576 4678
rect 7534 4562 7586 4574
rect 7534 4498 7586 4510
rect 16886 4562 16938 4574
rect 16886 4498 16938 4510
rect 24222 4562 24274 4574
rect 24222 4498 24274 4510
rect 29598 4450 29650 4462
rect 29598 4386 29650 4398
rect 7870 4338 7922 4350
rect 20066 4330 20078 4382
rect 20130 4330 20142 4382
rect 23886 4338 23938 4350
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 7870 4274 7922 4286
rect 23886 4274 23938 4286
rect 26910 4338 26962 4350
rect 30214 4338 30266 4350
rect 27682 4286 27694 4338
rect 27746 4286 27758 4338
rect 26910 4274 26962 4286
rect 30214 4274 30266 4286
rect 19954 4174 19966 4226
rect 20018 4174 20030 4226
rect 1344 3946 44576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 44576 3946
rect 1344 3860 44576 3894
rect 1344 3162 44576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 44576 3162
rect 1344 3076 44576 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 5014 41918 5066 41970
rect 5742 41918 5794 41970
rect 8822 41918 8874 41970
rect 9550 41918 9602 41970
rect 13470 41945 13522 41997
rect 17278 41945 17330 41997
rect 21086 41945 21138 41997
rect 24894 41945 24946 41997
rect 28702 41945 28754 41997
rect 32510 41945 32562 41997
rect 36318 41945 36370 41997
rect 40126 41945 40178 41997
rect 14478 41806 14530 41858
rect 18286 41806 18338 41858
rect 22094 41806 22146 41858
rect 25902 41806 25954 41858
rect 29710 41806 29762 41858
rect 33518 41806 33570 41858
rect 37326 41806 37378 41858
rect 41134 41806 41186 41858
rect 6078 41694 6130 41746
rect 9886 41694 9938 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 41806 41106 41858 41158
rect 43710 41134 43762 41186
rect 9326 40910 9378 40962
rect 9886 40910 9938 40962
rect 32790 40910 32842 40962
rect 36374 40910 36426 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 39678 40574 39730 40626
rect 11790 40462 11842 40514
rect 21086 40462 21138 40514
rect 24558 40462 24610 40514
rect 28702 40462 28754 40514
rect 32398 40462 32450 40514
rect 35982 40462 36034 40514
rect 39006 40462 39058 40514
rect 2158 40350 2210 40402
rect 5462 40350 5514 40402
rect 5742 40350 5794 40402
rect 8430 40350 8482 40402
rect 9046 40350 9098 40402
rect 14478 40350 14530 40402
rect 18398 40350 18450 40402
rect 21870 40350 21922 40402
rect 25398 40350 25450 40402
rect 26014 40350 26066 40402
rect 29318 40350 29370 40402
rect 29710 40350 29762 40402
rect 33294 40350 33346 40402
rect 36374 40350 36426 40402
rect 39342 40350 39394 40402
rect 40406 40350 40458 40402
rect 40798 40350 40850 40402
rect 2942 40238 2994 40290
rect 4846 40238 4898 40290
rect 6526 40238 6578 40290
rect 13694 40238 13746 40290
rect 19182 40238 19234 40290
rect 22654 40238 22706 40290
rect 26798 40238 26850 40290
rect 30494 40238 30546 40290
rect 34078 40238 34130 40290
rect 37102 40238 37154 40290
rect 41582 40238 41634 40290
rect 43486 40238 43538 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 13918 39790 13970 39842
rect 20190 39790 20242 39842
rect 24446 39790 24498 39842
rect 23662 39734 23714 39786
rect 30270 39790 30322 39842
rect 32846 39790 32898 39842
rect 37214 39790 37266 39842
rect 41022 39790 41074 39842
rect 42590 39790 42642 39842
rect 5070 39678 5122 39730
rect 15822 39678 15874 39730
rect 17726 39678 17778 39730
rect 4622 39566 4674 39618
rect 4958 39522 5010 39574
rect 9009 39566 9061 39618
rect 9886 39566 9938 39618
rect 12238 39566 12290 39618
rect 13022 39566 13074 39618
rect 14254 39566 14306 39618
rect 18510 39566 18562 39618
rect 20526 39566 20578 39618
rect 23550 39566 23602 39618
rect 23774 39566 23826 39618
rect 24110 39566 24162 39618
rect 29038 39566 29090 39618
rect 29262 39566 29314 39618
rect 29542 39566 29594 39618
rect 29934 39566 29986 39618
rect 32510 39566 32562 39618
rect 36878 39566 36930 39618
rect 40686 39566 40738 39618
rect 42926 39566 42978 39618
rect 43318 39566 43370 39618
rect 8766 39454 8818 39506
rect 10334 39454 10386 39506
rect 36150 39342 36202 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 16046 39006 16098 39058
rect 2830 38894 2882 38946
rect 7758 38894 7810 38946
rect 2662 38782 2714 38834
rect 3054 38782 3106 38834
rect 3278 38810 3330 38862
rect 3950 38820 4002 38872
rect 4286 38782 4338 38834
rect 4510 38782 4562 38834
rect 5070 38797 5122 38849
rect 5294 38782 5346 38834
rect 8094 38782 8146 38834
rect 4678 38726 4730 38778
rect 13470 38782 13522 38834
rect 16382 38782 16434 38834
rect 24168 38782 24220 38834
rect 24334 38782 24386 38834
rect 24446 38782 24498 38834
rect 28366 38782 28418 38834
rect 28702 38797 28754 38849
rect 36094 38782 36146 38834
rect 36206 38782 36258 38834
rect 36392 38819 36444 38871
rect 4958 38670 5010 38722
rect 23774 38670 23826 38722
rect 28814 38670 28866 38722
rect 35814 38670 35866 38722
rect 36766 38670 36818 38722
rect 13806 38558 13858 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 3950 38222 4002 38274
rect 23438 38222 23490 38274
rect 4510 37998 4562 38050
rect 4622 37998 4674 38050
rect 4344 37942 4396 37994
rect 23832 37998 23884 38050
rect 23998 37998 24050 38050
rect 24110 37998 24162 38050
rect 29038 37998 29090 38050
rect 29262 37998 29314 38050
rect 29822 37998 29874 38050
rect 39678 37998 39730 38050
rect 40462 37998 40514 38050
rect 29542 37886 29594 37938
rect 42366 37886 42418 37938
rect 5126 37774 5178 37826
rect 17502 37774 17554 37826
rect 18398 37774 18450 37826
rect 30158 37774 30210 37826
rect 39510 37774 39562 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 9718 37438 9770 37490
rect 21702 37438 21754 37490
rect 26686 37326 26738 37378
rect 3950 37214 4002 37266
rect 4690 37252 4742 37304
rect 5126 37214 5178 37266
rect 17390 37214 17442 37266
rect 17502 37214 17554 37266
rect 17648 37251 17700 37303
rect 21310 37214 21362 37266
rect 25454 37247 25506 37299
rect 25902 37250 25954 37302
rect 26350 37270 26402 37322
rect 26506 37247 26558 37299
rect 27582 37214 27634 37266
rect 27918 37214 27970 37266
rect 41134 37214 41186 37266
rect 3838 37046 3890 37098
rect 18062 37102 18114 37154
rect 18622 37102 18674 37154
rect 20526 37102 20578 37154
rect 28030 37046 28082 37098
rect 40966 36990 41018 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19518 36654 19570 36706
rect 25006 36542 25058 36594
rect 32958 36542 33010 36594
rect 40126 36542 40178 36594
rect 6526 36430 6578 36482
rect 7310 36430 7362 36482
rect 12014 36430 12066 36482
rect 12798 36430 12850 36482
rect 40798 36486 40850 36538
rect 19182 36430 19234 36482
rect 25230 36430 25282 36482
rect 9214 36318 9266 36370
rect 10110 36318 10162 36370
rect 24838 36374 24890 36426
rect 25566 36392 25618 36444
rect 33742 36430 33794 36482
rect 31054 36318 31106 36370
rect 39958 36374 40010 36426
rect 40574 36374 40626 36426
rect 18454 36206 18506 36258
rect 34134 36206 34186 36258
rect 37158 36206 37210 36258
rect 41302 36206 41354 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 6638 35870 6690 35922
rect 11678 35870 11730 35922
rect 9905 35702 9957 35754
rect 6302 35646 6354 35698
rect 10782 35646 10834 35698
rect 12014 35646 12066 35698
rect 13358 35646 13410 35698
rect 13918 35646 13970 35698
rect 14366 35646 14418 35698
rect 18398 35646 18450 35698
rect 28702 35646 28754 35698
rect 28814 35646 28866 35698
rect 28960 35684 29012 35736
rect 29822 35646 29874 35698
rect 30158 35646 30210 35698
rect 33966 35646 34018 35698
rect 36654 35646 36706 35698
rect 39994 35702 40046 35754
rect 37102 35646 37154 35698
rect 37978 35646 38030 35698
rect 39118 35646 39170 35698
rect 41134 35646 41186 35698
rect 29374 35534 29426 35586
rect 34750 35534 34802 35586
rect 38838 35534 38890 35586
rect 41918 35534 41970 35586
rect 43822 35534 43874 35586
rect 14142 35478 14194 35530
rect 9662 35422 9714 35474
rect 14702 35422 14754 35474
rect 29934 35478 29986 35530
rect 18734 35422 18786 35474
rect 25342 35422 25394 35474
rect 26574 35422 26626 35474
rect 38222 35422 38274 35474
rect 40238 35422 40290 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19238 35086 19290 35138
rect 25230 35086 25282 35138
rect 26854 35086 26906 35138
rect 39174 35086 39226 35138
rect 16942 34974 16994 35026
rect 29262 34974 29314 35026
rect 37158 34974 37210 35026
rect 5854 34862 5906 34914
rect 6414 34862 6466 34914
rect 7030 34862 7082 34914
rect 6078 34806 6130 34858
rect 15262 34862 15314 34914
rect 16606 34862 16658 34914
rect 17278 34862 17330 34914
rect 14385 34806 14437 34858
rect 16942 34806 16994 34858
rect 17614 34862 17666 34914
rect 18510 34862 18562 34914
rect 18958 34862 19010 34914
rect 18678 34806 18730 34858
rect 24838 34862 24890 34914
rect 25622 34862 25674 34914
rect 25790 34862 25842 34914
rect 25902 34862 25954 34914
rect 26686 34862 26738 34914
rect 27358 34862 27410 34914
rect 27806 34862 27858 34914
rect 28254 34862 28306 34914
rect 28478 34862 28530 34914
rect 29150 34862 29202 34914
rect 29822 34862 29874 34914
rect 14142 34750 14194 34802
rect 6302 34694 6354 34746
rect 18846 34750 18898 34802
rect 29598 34806 29650 34858
rect 30158 34862 30210 34914
rect 36430 34862 36482 34914
rect 38446 34862 38498 34914
rect 38894 34862 38946 34914
rect 38614 34806 38666 34858
rect 39678 34862 39730 34914
rect 40126 34862 40178 34914
rect 27918 34750 27970 34802
rect 39846 34806 39898 34858
rect 40406 34862 40458 34914
rect 40966 34862 41018 34914
rect 41134 34862 41186 34914
rect 41358 34862 41410 34914
rect 41582 34834 41634 34886
rect 42814 34862 42866 34914
rect 38782 34750 38834 34802
rect 40014 34750 40066 34802
rect 36262 34638 36314 34690
rect 42646 34638 42698 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 23662 34302 23714 34354
rect 13862 34190 13914 34242
rect 28366 34246 28418 34298
rect 3278 34093 3330 34145
rect 3614 34078 3666 34130
rect 4734 34078 4786 34130
rect 4958 34078 5010 34130
rect 5630 34078 5682 34130
rect 5966 34093 6018 34145
rect 14142 34106 14194 34158
rect 14310 34134 14362 34186
rect 17446 34190 17498 34242
rect 18902 34190 18954 34242
rect 30158 34190 30210 34242
rect 14590 34106 14642 34158
rect 14702 34134 14754 34186
rect 16214 34134 16266 34186
rect 16046 34078 16098 34130
rect 16382 34078 16434 34130
rect 16494 34078 16546 34130
rect 16774 34078 16826 34130
rect 17726 34078 17778 34130
rect 17838 34078 17890 34130
rect 3166 33966 3218 34018
rect 5238 33966 5290 34018
rect 6078 33966 6130 34018
rect 15206 33966 15258 34018
rect 18006 34022 18058 34074
rect 18174 34078 18226 34130
rect 18398 34078 18450 34130
rect 18622 34078 18674 34130
rect 19406 34078 19458 34130
rect 19630 34078 19682 34130
rect 21982 34078 22034 34130
rect 22318 34078 22370 34130
rect 23326 34078 23378 34130
rect 27806 34078 27858 34130
rect 28030 34117 28082 34169
rect 28478 34078 28530 34130
rect 30606 34106 30658 34158
rect 30830 34134 30882 34186
rect 36094 34190 36146 34242
rect 35646 34106 35698 34158
rect 35870 34078 35922 34130
rect 19294 33910 19346 33962
rect 20246 33966 20298 34018
rect 21254 33966 21306 34018
rect 23046 33966 23098 34018
rect 27302 33966 27354 34018
rect 29990 34022 30042 34074
rect 36262 34022 36314 34074
rect 21646 33854 21698 33906
rect 22486 33854 22538 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 6022 33518 6074 33570
rect 6806 33518 6858 33570
rect 18846 33518 18898 33570
rect 24558 33518 24610 33570
rect 2606 33406 2658 33458
rect 5126 33406 5178 33458
rect 22598 33406 22650 33458
rect 29374 33462 29426 33514
rect 1822 33294 1874 33346
rect 5630 33294 5682 33346
rect 5742 33294 5794 33346
rect 6302 33294 6354 33346
rect 6526 33294 6578 33346
rect 8766 33294 8818 33346
rect 18174 33294 18226 33346
rect 18286 33294 18338 33346
rect 18452 33294 18504 33346
rect 19462 33294 19514 33346
rect 21646 33294 21698 33346
rect 23438 33294 23490 33346
rect 23662 33294 23714 33346
rect 23942 33294 23994 33346
rect 24222 33294 24274 33346
rect 29486 33294 29538 33346
rect 29822 33294 29874 33346
rect 32510 33294 32562 33346
rect 4510 33182 4562 33234
rect 8430 33070 8482 33122
rect 21982 33070 22034 33122
rect 23270 33070 23322 33122
rect 32846 33070 32898 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 31278 32622 31330 32674
rect 36374 32622 36426 32674
rect 36766 32622 36818 32674
rect 41246 32622 41298 32674
rect 4286 32510 4338 32562
rect 4622 32510 4674 32562
rect 4958 32510 5010 32562
rect 5406 32510 5458 32562
rect 5854 32510 5906 32562
rect 6302 32549 6354 32601
rect 6526 32510 6578 32562
rect 21870 32510 21922 32562
rect 22654 32510 22706 32562
rect 28590 32510 28642 32562
rect 29374 32510 29426 32562
rect 36654 32510 36706 32562
rect 4062 32398 4114 32450
rect 6190 32398 6242 32450
rect 7254 32398 7306 32450
rect 16214 32398 16266 32450
rect 24558 32398 24610 32450
rect 25398 32398 25450 32450
rect 31894 32398 31946 32450
rect 36934 32454 36986 32506
rect 37102 32510 37154 32562
rect 37326 32510 37378 32562
rect 37662 32510 37714 32562
rect 41078 32566 41130 32618
rect 40910 32510 40962 32562
rect 41358 32510 41410 32562
rect 41638 32286 41690 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 30494 31950 30546 32002
rect 16662 31838 16714 31890
rect 23382 31838 23434 31890
rect 27750 31838 27802 31890
rect 33462 31838 33514 31890
rect 6881 31726 6933 31778
rect 7758 31726 7810 31778
rect 11790 31726 11842 31778
rect 12574 31726 12626 31778
rect 13806 31698 13858 31750
rect 16158 31726 16210 31778
rect 16382 31726 16434 31778
rect 17166 31726 17218 31778
rect 42086 31782 42138 31834
rect 22430 31726 22482 31778
rect 25790 31726 25842 31778
rect 28366 31726 28418 31778
rect 29150 31698 29202 31750
rect 33630 31726 33682 31778
rect 34414 31726 34466 31778
rect 36318 31726 36370 31778
rect 36878 31726 36930 31778
rect 41470 31698 41522 31750
rect 41694 31726 41746 31778
rect 6638 31614 6690 31666
rect 9886 31614 9938 31666
rect 41918 31614 41970 31666
rect 5910 31502 5962 31554
rect 14814 31502 14866 31554
rect 17502 31502 17554 31554
rect 22766 31502 22818 31554
rect 25958 31502 26010 31554
rect 28198 31502 28250 31554
rect 37046 31502 37098 31554
rect 39342 31502 39394 31554
rect 40294 31502 40346 31554
rect 40966 31502 41018 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 5630 31166 5682 31218
rect 5910 31166 5962 31218
rect 32566 31166 32618 31218
rect 40294 31166 40346 31218
rect 27134 31054 27186 31106
rect 9994 30980 10046 31032
rect 10670 30942 10722 30994
rect 11678 30942 11730 30994
rect 12238 30942 12290 30994
rect 14926 30969 14978 31021
rect 16270 30942 16322 30994
rect 16606 30942 16658 30994
rect 17950 30942 18002 30994
rect 18846 30986 18898 31038
rect 26462 30998 26514 31050
rect 35982 31054 36034 31106
rect 28142 30998 28194 31050
rect 28478 30998 28530 31050
rect 19182 30942 19234 30994
rect 27582 30942 27634 30994
rect 33070 30969 33122 31021
rect 36206 30942 36258 30994
rect 36430 30970 36482 31022
rect 41134 30942 41186 30994
rect 41918 30942 41970 30994
rect 35814 30886 35866 30938
rect 10782 30774 10834 30826
rect 12462 30774 12514 30826
rect 16158 30774 16210 30826
rect 17558 30830 17610 30882
rect 18734 30830 18786 30882
rect 34078 30830 34130 30882
rect 43822 30830 43874 30882
rect 18286 30718 18338 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 12126 30382 12178 30434
rect 39902 30382 39954 30434
rect 41974 30382 42026 30434
rect 19966 30270 20018 30322
rect 8150 30158 8202 30210
rect 8318 30158 8370 30210
rect 9438 30158 9490 30210
rect 11678 30130 11730 30182
rect 12462 30158 12514 30210
rect 17110 30214 17162 30266
rect 12854 30158 12906 30210
rect 14926 30158 14978 30210
rect 15598 30158 15650 30210
rect 16718 30158 16770 30210
rect 15374 30102 15426 30154
rect 16494 30102 16546 30154
rect 20078 30114 20130 30166
rect 20414 30158 20466 30210
rect 26518 30142 26570 30194
rect 16942 30046 16994 30098
rect 15150 29990 15202 30042
rect 17558 30046 17610 30098
rect 26686 30102 26738 30154
rect 26910 30102 26962 30154
rect 27134 30130 27186 30182
rect 27414 30158 27466 30210
rect 39230 30158 39282 30210
rect 39342 30158 39394 30210
rect 40350 30158 40402 30210
rect 41226 30158 41278 30210
rect 42142 30158 42194 30210
rect 39510 30102 39562 30154
rect 21478 30046 21530 30098
rect 41470 30046 41522 30098
rect 29262 29934 29314 29986
rect 29822 29934 29874 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 22038 29598 22090 29650
rect 3726 29389 3778 29441
rect 6358 29430 6410 29482
rect 4062 29374 4114 29426
rect 6078 29374 6130 29426
rect 6750 29374 6802 29426
rect 6974 29374 7026 29426
rect 10106 29412 10158 29464
rect 10782 29374 10834 29426
rect 11566 29374 11618 29426
rect 11902 29374 11954 29426
rect 15262 29374 15314 29426
rect 15542 29403 15594 29455
rect 20750 29374 20802 29426
rect 20862 29374 20914 29426
rect 21048 29412 21100 29464
rect 26910 29374 26962 29426
rect 33630 29374 33682 29426
rect 3614 29262 3666 29314
rect 6526 29262 6578 29314
rect 15710 29262 15762 29314
rect 16214 29262 16266 29314
rect 10558 29206 10610 29258
rect 20470 29262 20522 29314
rect 40070 29262 40122 29314
rect 7254 29150 7306 29202
rect 21422 29150 21474 29202
rect 27246 29150 27298 29202
rect 27806 29150 27858 29202
rect 29038 29150 29090 29202
rect 33294 29150 33346 29202
rect 33966 29150 34018 29202
rect 34414 29150 34466 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 8206 28758 8258 28810
rect 20638 28814 20690 28866
rect 29878 28814 29930 28866
rect 2606 28702 2658 28754
rect 27246 28758 27298 28810
rect 34414 28814 34466 28866
rect 39230 28814 39282 28866
rect 39678 28814 39730 28866
rect 10222 28702 10274 28754
rect 11006 28702 11058 28754
rect 19518 28702 19570 28754
rect 25062 28702 25114 28754
rect 33294 28702 33346 28754
rect 1822 28590 1874 28642
rect 4510 28590 4562 28642
rect 5126 28590 5178 28642
rect 7758 28590 7810 28642
rect 8094 28590 8146 28642
rect 9886 28590 9938 28642
rect 10446 28590 10498 28642
rect 10894 28590 10946 28642
rect 11566 28590 11618 28642
rect 19070 28590 19122 28642
rect 10278 28534 10330 28586
rect 11174 28534 11226 28586
rect 19406 28546 19458 28598
rect 20302 28590 20354 28642
rect 21982 28590 22034 28642
rect 23886 28590 23938 28642
rect 24670 28590 24722 28642
rect 26462 28590 26514 28642
rect 27022 28590 27074 28642
rect 29150 28590 29202 28642
rect 29598 28590 29650 28642
rect 29318 28534 29370 28586
rect 31390 28590 31442 28642
rect 34078 28590 34130 28642
rect 34808 28590 34860 28642
rect 34974 28590 35026 28642
rect 35086 28590 35138 28642
rect 35422 28590 35474 28642
rect 35870 28590 35922 28642
rect 35590 28534 35642 28586
rect 29486 28478 29538 28530
rect 35758 28478 35810 28530
rect 36150 28478 36202 28530
rect 39454 28366 39506 28418
rect 40126 28366 40178 28418
rect 40686 28366 40738 28418
rect 41582 28366 41634 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 6134 28030 6186 28082
rect 18790 28030 18842 28082
rect 4622 27918 4674 27970
rect 10110 27974 10162 28026
rect 17502 27974 17554 28026
rect 34246 28030 34298 28082
rect 35142 28030 35194 28082
rect 37102 28030 37154 28082
rect 39118 28030 39170 28082
rect 5686 27918 5738 27970
rect 37942 27918 37994 27970
rect 10334 27862 10386 27914
rect 4062 27806 4114 27858
rect 4286 27806 4338 27858
rect 4846 27806 4898 27858
rect 5070 27806 5122 27858
rect 9998 27806 10050 27858
rect 10670 27806 10722 27858
rect 13694 27806 13746 27858
rect 14030 27833 14082 27885
rect 14366 27806 14418 27858
rect 17838 27862 17890 27914
rect 41246 27918 41298 27970
rect 14702 27806 14754 27858
rect 17390 27806 17442 27858
rect 18062 27806 18114 27858
rect 25566 27806 25618 27858
rect 25902 27833 25954 27885
rect 26238 27806 26290 27858
rect 26574 27806 26626 27858
rect 28926 27806 28978 27858
rect 29262 27806 29314 27858
rect 29822 27806 29874 27858
rect 30046 27806 30098 27858
rect 36766 27806 36818 27858
rect 38110 27806 38162 27858
rect 38446 27806 38498 27858
rect 39454 27806 39506 27858
rect 40910 27806 40962 27858
rect 13918 27694 13970 27746
rect 24726 27694 24778 27746
rect 25678 27694 25730 27746
rect 29038 27638 29090 27690
rect 29710 27638 29762 27690
rect 36598 27694 36650 27746
rect 41078 27750 41130 27802
rect 41358 27806 41410 27858
rect 41638 27582 41690 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 6302 27246 6354 27298
rect 14814 27134 14866 27186
rect 22598 27134 22650 27186
rect 23550 27134 23602 27186
rect 28142 27190 28194 27242
rect 35926 27246 35978 27298
rect 37214 27246 37266 27298
rect 37886 27246 37938 27298
rect 39846 27246 39898 27298
rect 40462 27246 40514 27298
rect 29934 27134 29986 27186
rect 7422 27022 7474 27074
rect 14366 27022 14418 27074
rect 6545 26966 6597 27018
rect 14702 26978 14754 27030
rect 21758 27022 21810 27074
rect 15318 26910 15370 26962
rect 18902 26910 18954 26962
rect 21422 26910 21474 26962
rect 22878 26966 22930 27018
rect 22990 26984 23042 27036
rect 28254 27022 28306 27074
rect 28590 27022 28642 27074
rect 29598 27022 29650 27074
rect 30270 27022 30322 27074
rect 35198 27022 35250 27074
rect 35534 27022 35586 27074
rect 35646 27022 35698 27074
rect 23718 26966 23770 27018
rect 29934 26966 29986 27018
rect 35366 26966 35418 27018
rect 36878 27022 36930 27074
rect 37550 27022 37602 27074
rect 39118 27022 39170 27074
rect 39286 27078 39338 27130
rect 39454 27022 39506 27074
rect 39566 27022 39618 27074
rect 41974 27078 42026 27130
rect 40126 27022 40178 27074
rect 41582 27022 41634 27074
rect 41414 26966 41466 27018
rect 36486 26910 36538 26962
rect 41806 26910 41858 26962
rect 34918 26798 34970 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 22710 26462 22762 26514
rect 15374 26406 15426 26458
rect 36542 26462 36594 26514
rect 18230 26350 18282 26402
rect 30606 26350 30658 26402
rect 9546 26276 9598 26328
rect 10222 26238 10274 26290
rect 13582 26238 13634 26290
rect 13918 26253 13970 26305
rect 14590 26238 14642 26290
rect 15150 26238 15202 26290
rect 18510 26238 18562 26290
rect 18622 26238 18674 26290
rect 19126 26294 19178 26346
rect 18958 26238 19010 26290
rect 19294 26238 19346 26290
rect 19406 26238 19458 26290
rect 22542 26238 22594 26290
rect 28254 26238 28306 26290
rect 28590 26265 28642 26317
rect 28926 26238 28978 26290
rect 29486 26238 29538 26290
rect 30362 26238 30414 26290
rect 33966 26238 34018 26290
rect 36878 26238 36930 26290
rect 37102 26238 37154 26290
rect 40406 26238 40458 26290
rect 41134 26238 41186 26290
rect 41918 26238 41970 26290
rect 14030 26126 14082 26178
rect 24278 26126 24330 26178
rect 28366 26126 28418 26178
rect 31222 26126 31274 26178
rect 43822 26126 43874 26178
rect 10334 26070 10386 26122
rect 19686 26014 19738 26066
rect 34302 26014 34354 26066
rect 37438 26014 37490 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 10670 25678 10722 25730
rect 18678 25678 18730 25730
rect 30830 25678 30882 25730
rect 9326 25622 9378 25674
rect 19294 25566 19346 25618
rect 24110 25566 24162 25618
rect 9326 25454 9378 25506
rect 10002 25416 10054 25468
rect 10334 25454 10386 25506
rect 13806 25454 13858 25506
rect 14682 25454 14734 25506
rect 18174 25454 18226 25506
rect 18398 25454 18450 25506
rect 19182 25454 19234 25506
rect 19854 25454 19906 25506
rect 19630 25398 19682 25450
rect 22990 25454 23042 25506
rect 25174 25510 25226 25562
rect 24894 25454 24946 25506
rect 25006 25454 25058 25506
rect 25342 25454 25394 25506
rect 23866 25398 23918 25450
rect 29710 25454 29762 25506
rect 30586 25454 30638 25506
rect 42814 25454 42866 25506
rect 14926 25342 14978 25394
rect 24614 25342 24666 25394
rect 25846 25342 25898 25394
rect 42646 25230 42698 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 6750 24894 6802 24946
rect 15094 24894 15146 24946
rect 23438 24894 23490 24946
rect 1934 24670 1986 24722
rect 4622 24670 4674 24722
rect 5966 24714 6018 24766
rect 6302 24670 6354 24722
rect 7086 24670 7138 24722
rect 13974 24726 14026 24778
rect 14254 24726 14306 24778
rect 14478 24698 14530 24750
rect 14590 24726 14642 24778
rect 19892 24708 19944 24760
rect 20078 24670 20130 24722
rect 20190 24670 20242 24722
rect 22934 24670 22986 24722
rect 23102 24670 23154 24722
rect 23774 24670 23826 24722
rect 34750 24670 34802 24722
rect 2718 24558 2770 24610
rect 5238 24558 5290 24610
rect 5854 24558 5906 24610
rect 19518 24558 19570 24610
rect 13750 24446 13802 24498
rect 23942 24446 23994 24498
rect 34414 24446 34466 24498
rect 35814 24446 35866 24498
rect 36318 24446 36370 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3166 24110 3218 24162
rect 11902 24110 11954 24162
rect 35814 24110 35866 24162
rect 4902 23998 4954 24050
rect 15094 23998 15146 24050
rect 22934 23998 22986 24050
rect 37102 24054 37154 24106
rect 3502 23886 3554 23938
rect 10110 23886 10162 23938
rect 11566 23886 11618 23938
rect 15262 23886 15314 23938
rect 23550 23886 23602 23938
rect 23998 23942 24050 23994
rect 24838 23942 24890 23994
rect 25286 23998 25338 24050
rect 23774 23886 23826 23938
rect 24110 23848 24162 23900
rect 36094 23886 36146 23938
rect 36318 23886 36370 23938
rect 36990 23886 37042 23938
rect 37326 23886 37378 23938
rect 37662 23886 37714 23938
rect 40014 23886 40066 23938
rect 40406 23886 40458 23938
rect 23270 23774 23322 23826
rect 24670 23774 24722 23826
rect 9774 23662 9826 23714
rect 15598 23662 15650 23714
rect 35478 23662 35530 23714
rect 37998 23662 38050 23714
rect 39846 23662 39898 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15878 23326 15930 23378
rect 3838 23270 3890 23322
rect 16606 23326 16658 23378
rect 14702 23214 14754 23266
rect 18566 23214 18618 23266
rect 21366 23214 21418 23266
rect 4286 23158 4338 23210
rect 5742 23158 5794 23210
rect 30382 23214 30434 23266
rect 3950 23102 4002 23154
rect 4622 23102 4674 23154
rect 5406 23102 5458 23154
rect 5966 23102 6018 23154
rect 6302 23102 6354 23154
rect 15038 23102 15090 23154
rect 15486 23102 15538 23154
rect 16270 23102 16322 23154
rect 18062 23102 18114 23154
rect 18286 23102 18338 23154
rect 21646 23129 21698 23181
rect 29262 23102 29314 23154
rect 30138 23102 30190 23154
rect 39566 23102 39618 23154
rect 39790 23102 39842 23154
rect 5630 22990 5682 23042
rect 36710 22990 36762 23042
rect 15318 22878 15370 22930
rect 22654 22878 22706 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 5686 22542 5738 22594
rect 28478 22542 28530 22594
rect 13694 22486 13746 22538
rect 30494 22542 30546 22594
rect 31950 22542 32002 22594
rect 4622 22430 4674 22482
rect 8766 22430 8818 22482
rect 10670 22430 10722 22482
rect 15598 22430 15650 22482
rect 16606 22430 16658 22482
rect 16830 22430 16882 22482
rect 16998 22430 17050 22482
rect 18958 22430 19010 22482
rect 34526 22430 34578 22482
rect 5070 22318 5122 22370
rect 5966 22318 6018 22370
rect 4790 22262 4842 22314
rect 6078 22318 6130 22370
rect 7982 22318 8034 22370
rect 11286 22318 11338 22370
rect 13582 22318 13634 22370
rect 13918 22318 13970 22370
rect 14926 22318 14978 22370
rect 15038 22318 15090 22370
rect 16382 22318 16434 22370
rect 15204 22262 15256 22314
rect 16606 22318 16658 22370
rect 17726 22318 17778 22370
rect 17950 22318 18002 22370
rect 18622 22318 18674 22370
rect 19294 22318 19346 22370
rect 18958 22262 19010 22314
rect 19630 22318 19682 22370
rect 23774 22318 23826 22370
rect 23998 22318 24050 22370
rect 27358 22318 27410 22370
rect 29374 22318 29426 22370
rect 30250 22318 30302 22370
rect 33070 22318 33122 22370
rect 28234 22262 28286 22314
rect 32193 22262 32245 22314
rect 33406 22318 33458 22370
rect 34282 22318 34334 22370
rect 34862 22318 34914 22370
rect 35982 22318 36034 22370
rect 36374 22318 36426 22370
rect 35646 22262 35698 22314
rect 39062 22318 39114 22370
rect 39342 22318 39394 22370
rect 39622 22374 39674 22426
rect 39790 22318 39842 22370
rect 40910 22318 40962 22370
rect 41694 22318 41746 22370
rect 16102 22206 16154 22258
rect 17558 22206 17610 22258
rect 18230 22206 18282 22258
rect 24278 22206 24330 22258
rect 35030 22150 35082 22202
rect 36206 22206 36258 22258
rect 39454 22206 39506 22258
rect 43598 22206 43650 22258
rect 40742 22094 40794 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 19462 21758 19514 21810
rect 34190 21758 34242 21810
rect 29486 21646 29538 21698
rect 10017 21590 10069 21642
rect 10894 21534 10946 21586
rect 11902 21572 11954 21624
rect 12014 21590 12066 21642
rect 11174 21478 11226 21530
rect 12518 21534 12570 21586
rect 15934 21534 15986 21586
rect 16158 21534 16210 21586
rect 16494 21534 16546 21586
rect 16830 21534 16882 21586
rect 20078 21534 20130 21586
rect 20302 21534 20354 21586
rect 28814 21590 28866 21642
rect 34862 21646 34914 21698
rect 41246 21646 41298 21698
rect 23774 21534 23826 21586
rect 29038 21564 29090 21616
rect 34526 21534 34578 21586
rect 36766 21534 36818 21586
rect 37550 21534 37602 21586
rect 29206 21478 29258 21530
rect 39566 21534 39618 21586
rect 39902 21534 39954 21586
rect 40014 21534 40066 21586
rect 11342 21422 11394 21474
rect 19798 21422 19850 21474
rect 37942 21422 37994 21474
rect 39734 21478 39786 21530
rect 41078 21590 41130 21642
rect 40910 21534 40962 21586
rect 41358 21534 41410 21586
rect 42814 21534 42866 21586
rect 16606 21366 16658 21418
rect 9774 21310 9826 21362
rect 15654 21310 15706 21362
rect 23438 21310 23490 21362
rect 40294 21310 40346 21362
rect 41638 21310 41690 21362
rect 42646 21310 42698 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 29542 20974 29594 21026
rect 12014 20918 12066 20970
rect 5630 20862 5682 20914
rect 13918 20862 13970 20914
rect 21870 20862 21922 20914
rect 23774 20862 23826 20914
rect 41470 20862 41522 20914
rect 5742 20706 5794 20758
rect 5966 20750 6018 20802
rect 11566 20750 11618 20802
rect 11902 20750 11954 20802
rect 13470 20750 13522 20802
rect 24558 20750 24610 20802
rect 13750 20694 13802 20746
rect 29038 20750 29090 20802
rect 41638 20806 41690 20858
rect 29262 20750 29314 20802
rect 41246 20750 41298 20802
rect 40910 20694 40962 20746
rect 24950 20526 25002 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 4286 20134 4338 20186
rect 11006 20078 11058 20130
rect 4622 20022 4674 20074
rect 12630 20078 12682 20130
rect 27806 20078 27858 20130
rect 33126 20134 33178 20186
rect 35366 20078 35418 20130
rect 35982 20078 36034 20130
rect 3502 19966 3554 20018
rect 4286 19966 4338 20018
rect 4846 19966 4898 20018
rect 5574 19966 5626 20018
rect 6190 19966 6242 20018
rect 6302 19966 6354 20018
rect 11249 19966 11301 20018
rect 12126 19966 12178 20018
rect 25118 19966 25170 20018
rect 28702 19966 28754 20018
rect 35814 20022 35866 20074
rect 29094 19966 29146 20018
rect 32062 19966 32114 20018
rect 33294 19966 33346 20018
rect 35646 19966 35698 20018
rect 36094 19966 36146 20018
rect 25902 19854 25954 19906
rect 3166 19742 3218 19794
rect 5910 19742 5962 19794
rect 28366 19742 28418 19794
rect 32230 19742 32282 19794
rect 36374 19742 36426 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 5910 19406 5962 19458
rect 11006 19406 11058 19458
rect 25902 19406 25954 19458
rect 39566 19406 39618 19458
rect 2606 19294 2658 19346
rect 4510 19294 4562 19346
rect 18174 19294 18226 19346
rect 1822 19182 1874 19234
rect 5126 19182 5178 19234
rect 6190 19182 6242 19234
rect 6414 19182 6466 19234
rect 6694 19182 6746 19234
rect 6974 19182 7026 19234
rect 7198 19182 7250 19234
rect 9438 19182 9490 19234
rect 9774 19155 9826 19207
rect 10110 19182 10162 19234
rect 10670 19182 10722 19234
rect 17782 19182 17834 19234
rect 20078 19182 20130 19234
rect 20862 19182 20914 19234
rect 34974 19238 35026 19290
rect 35814 19238 35866 19290
rect 26238 19182 26290 19234
rect 39230 19182 39282 19234
rect 40742 19238 40794 19290
rect 41134 19182 41186 19234
rect 35254 19126 35306 19178
rect 41358 19154 41410 19206
rect 35646 19070 35698 19122
rect 9998 19014 10050 19066
rect 40910 19070 40962 19122
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 41190 18622 41242 18674
rect 10390 18510 10442 18562
rect 26574 18566 26626 18618
rect 15598 18510 15650 18562
rect 33406 18510 33458 18562
rect 9998 18398 10050 18450
rect 14702 18398 14754 18450
rect 14814 18398 14866 18450
rect 15206 18398 15258 18450
rect 15486 18398 15538 18450
rect 14086 18286 14138 18338
rect 15766 18342 15818 18394
rect 15934 18398 15986 18450
rect 16326 18398 16378 18450
rect 16606 18398 16658 18450
rect 16718 18398 16770 18450
rect 17838 18398 17890 18450
rect 19966 18398 20018 18450
rect 26910 18454 26962 18506
rect 20078 18398 20130 18450
rect 20358 18398 20410 18450
rect 20638 18398 20690 18450
rect 26462 18398 26514 18450
rect 27134 18398 27186 18450
rect 27806 18413 27858 18465
rect 28142 18398 28194 18450
rect 28758 18398 28810 18450
rect 28926 18398 28978 18450
rect 29150 18398 29202 18450
rect 31034 18454 31086 18506
rect 30158 18398 30210 18450
rect 31278 18398 31330 18450
rect 35310 18398 35362 18450
rect 36094 18398 36146 18450
rect 36486 18398 36538 18450
rect 38670 18398 38722 18450
rect 39006 18398 39058 18450
rect 39118 18398 39170 18450
rect 39454 18398 39506 18450
rect 41022 18398 41074 18450
rect 21590 18286 21642 18338
rect 26182 18286 26234 18338
rect 27694 18286 27746 18338
rect 29430 18286 29482 18338
rect 9662 18174 9714 18226
rect 14422 18174 14474 18226
rect 17502 18174 17554 18226
rect 20974 18174 21026 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 21366 17838 21418 17890
rect 37326 17838 37378 17890
rect 37998 17838 38050 17890
rect 38558 17838 38610 17890
rect 39118 17838 39170 17890
rect 39454 17838 39506 17890
rect 8766 17726 8818 17778
rect 10670 17726 10722 17778
rect 14198 17726 14250 17778
rect 15374 17726 15426 17778
rect 40742 17726 40794 17778
rect 41694 17726 41746 17778
rect 43598 17726 43650 17778
rect 7982 17614 8034 17666
rect 14702 17614 14754 17666
rect 15038 17614 15090 17666
rect 15710 17614 15762 17666
rect 17390 17614 17442 17666
rect 15430 17558 15482 17610
rect 21646 17614 21698 17666
rect 21870 17614 21922 17666
rect 22262 17614 22314 17666
rect 33406 17586 33458 17638
rect 35646 17614 35698 17666
rect 36990 17614 37042 17666
rect 37662 17614 37714 17666
rect 40910 17614 40962 17666
rect 11286 17390 11338 17442
rect 17726 17390 17778 17442
rect 27414 17390 27466 17442
rect 33126 17390 33178 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 21702 17054 21754 17106
rect 22206 17054 22258 17106
rect 33686 17054 33738 17106
rect 34190 17054 34242 17106
rect 37494 16942 37546 16994
rect 14478 16830 14530 16882
rect 14702 16830 14754 16882
rect 21030 16886 21082 16938
rect 20750 16830 20802 16882
rect 20862 16830 20914 16882
rect 21198 16830 21250 16882
rect 21870 16830 21922 16882
rect 28030 16830 28082 16882
rect 28366 16830 28418 16882
rect 28870 16830 28922 16882
rect 29150 16830 29202 16882
rect 29262 16830 29314 16882
rect 33854 16830 33906 16882
rect 39174 16886 39226 16938
rect 39006 16830 39058 16882
rect 39342 16830 39394 16882
rect 39454 16830 39506 16882
rect 14982 16606 15034 16658
rect 20470 16606 20522 16658
rect 39734 16606 39786 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 30158 16270 30210 16322
rect 24950 16158 25002 16210
rect 27862 16158 27914 16210
rect 14926 16046 14978 16098
rect 21478 16046 21530 16098
rect 23046 16046 23098 16098
rect 23214 16046 23266 16098
rect 28142 16046 28194 16098
rect 28254 16046 28306 16098
rect 29150 16018 29202 16070
rect 39566 16046 39618 16098
rect 28534 15934 28586 15986
rect 15262 15822 15314 15874
rect 23550 15822 23602 15874
rect 39230 15822 39282 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 17558 15486 17610 15538
rect 23886 15486 23938 15538
rect 32566 15486 32618 15538
rect 27806 15374 27858 15426
rect 30046 15374 30098 15426
rect 4510 15262 4562 15314
rect 7814 15262 7866 15314
rect 9438 15262 9490 15314
rect 10334 15289 10386 15341
rect 14030 15262 14082 15314
rect 14814 15262 14866 15314
rect 23550 15262 23602 15314
rect 24782 15262 24834 15314
rect 29878 15318 29930 15370
rect 38334 15374 38386 15426
rect 25118 15262 25170 15314
rect 28366 15262 28418 15314
rect 28590 15262 28642 15314
rect 29038 15262 29090 15314
rect 29710 15262 29762 15314
rect 30158 15262 30210 15314
rect 30438 15262 30490 15314
rect 30942 15262 30994 15314
rect 31166 15306 31218 15358
rect 31614 15262 31666 15314
rect 31950 15277 32002 15329
rect 34638 15306 34690 15358
rect 34974 15262 35026 15314
rect 37998 15262 38050 15314
rect 38166 15262 38218 15314
rect 38446 15262 38498 15314
rect 38726 15262 38778 15314
rect 39566 15262 39618 15314
rect 39678 15262 39730 15314
rect 39824 15299 39876 15351
rect 5294 15150 5346 15202
rect 7198 15150 7250 15202
rect 11006 15150 11058 15202
rect 12966 15150 13018 15202
rect 13862 15150 13914 15202
rect 16718 15150 16770 15202
rect 24446 15150 24498 15202
rect 25902 15150 25954 15202
rect 31278 15150 31330 15202
rect 32062 15150 32114 15202
rect 34246 15150 34298 15202
rect 34526 15150 34578 15202
rect 28366 15094 28418 15146
rect 40238 15038 40290 15090
rect 41022 15038 41074 15090
rect 41918 15038 41970 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 15374 14702 15426 14754
rect 40798 14702 40850 14754
rect 5854 14590 5906 14642
rect 17334 14590 17386 14642
rect 25622 14590 25674 14642
rect 27022 14590 27074 14642
rect 28198 14590 28250 14642
rect 29542 14590 29594 14642
rect 30046 14590 30098 14642
rect 31950 14590 32002 14642
rect 33126 14590 33178 14642
rect 40294 14590 40346 14642
rect 41918 14590 41970 14642
rect 43822 14590 43874 14642
rect 5966 14463 6018 14515
rect 6302 14478 6354 14530
rect 6750 14478 6802 14530
rect 7870 14478 7922 14530
rect 6993 14422 7045 14474
rect 12126 14434 12178 14486
rect 12462 14478 12514 14530
rect 14142 14478 14194 14530
rect 14702 14450 14754 14502
rect 25230 14478 25282 14530
rect 27134 14434 27186 14486
rect 27470 14478 27522 14530
rect 32734 14478 32786 14530
rect 33798 14478 33850 14530
rect 34078 14478 34130 14530
rect 34414 14451 34466 14503
rect 34750 14478 34802 14530
rect 38894 14478 38946 14530
rect 39006 14478 39058 14530
rect 39342 14478 39394 14530
rect 9942 14366 9994 14418
rect 39174 14422 39226 14474
rect 40462 14478 40514 14530
rect 41134 14478 41186 14530
rect 38614 14366 38666 14418
rect 12350 14310 12402 14362
rect 20358 14254 20410 14306
rect 34302 14310 34354 14362
rect 24894 14254 24946 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 7198 13918 7250 13970
rect 7870 13918 7922 13970
rect 15654 13918 15706 13970
rect 27134 13918 27186 13970
rect 28366 13918 28418 13970
rect 36934 13918 36986 13970
rect 14814 13862 14866 13914
rect 36318 13806 36370 13858
rect 10446 13694 10498 13746
rect 13134 13694 13186 13746
rect 13582 13694 13634 13746
rect 13694 13694 13746 13746
rect 13862 13694 13914 13746
rect 14702 13694 14754 13746
rect 15038 13738 15090 13790
rect 19742 13738 19794 13790
rect 20078 13694 20130 13746
rect 20302 13694 20354 13746
rect 20526 13694 20578 13746
rect 21086 13694 21138 13746
rect 21310 13694 21362 13746
rect 33630 13694 33682 13746
rect 11230 13582 11282 13634
rect 19630 13582 19682 13634
rect 34414 13582 34466 13634
rect 14254 13470 14306 13522
rect 20806 13470 20858 13522
rect 21590 13470 21642 13522
rect 27470 13470 27522 13522
rect 28142 13470 28194 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 8654 13078 8706 13130
rect 13526 13134 13578 13186
rect 34638 13134 34690 13186
rect 9438 13022 9490 13074
rect 11230 13022 11282 13074
rect 17558 13022 17610 13074
rect 18510 13022 18562 13074
rect 20414 13022 20466 13074
rect 38222 13022 38274 13074
rect 40574 13022 40626 13074
rect 7422 12910 7474 12962
rect 7030 12854 7082 12906
rect 7646 12882 7698 12934
rect 8206 12910 8258 12962
rect 8542 12910 8594 12962
rect 8990 12910 9042 12962
rect 9326 12895 9378 12947
rect 11342 12895 11394 12947
rect 11566 12910 11618 12962
rect 12238 12910 12290 12962
rect 12574 12883 12626 12935
rect 12910 12910 12962 12962
rect 13694 12910 13746 12962
rect 17726 12910 17778 12962
rect 21310 12910 21362 12962
rect 21982 12910 22034 12962
rect 21758 12854 21810 12906
rect 34302 12910 34354 12962
rect 38334 12866 38386 12918
rect 38670 12910 38722 12962
rect 39902 12910 39954 12962
rect 40014 12910 40066 12962
rect 40180 12910 40232 12962
rect 7198 12798 7250 12850
rect 12574 12742 12626 12794
rect 14086 12686 14138 12738
rect 21646 12742 21698 12794
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4958 12238 5010 12290
rect 20078 12238 20130 12290
rect 2270 12126 2322 12178
rect 5574 12126 5626 12178
rect 12574 12126 12626 12178
rect 12910 12153 12962 12205
rect 13246 12126 13298 12178
rect 13582 12126 13634 12178
rect 16886 12126 16938 12178
rect 17390 12126 17442 12178
rect 20638 12126 20690 12178
rect 20974 12126 21026 12178
rect 39156 12164 39208 12216
rect 39342 12126 39394 12178
rect 39454 12126 39506 12178
rect 41134 12126 41186 12178
rect 3054 12014 3106 12066
rect 12798 12014 12850 12066
rect 18174 12014 18226 12066
rect 20526 11958 20578 12010
rect 21478 12014 21530 12066
rect 38782 11902 38834 11954
rect 41470 11902 41522 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 3726 11566 3778 11618
rect 19742 11454 19794 11506
rect 40854 11454 40906 11506
rect 41806 11454 41858 11506
rect 43710 11454 43762 11506
rect 4062 11342 4114 11394
rect 6750 11342 6802 11394
rect 7198 11303 7250 11355
rect 7422 11342 7474 11394
rect 19854 11327 19906 11379
rect 20190 11342 20242 11394
rect 27918 11342 27970 11394
rect 38894 11342 38946 11394
rect 41022 11342 41074 11394
rect 6862 11174 6914 11226
rect 28254 11118 28306 11170
rect 38558 11118 38610 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 12966 10782 13018 10834
rect 24614 10726 24666 10778
rect 26518 10782 26570 10834
rect 36710 10782 36762 10834
rect 22486 10670 22538 10722
rect 39566 10670 39618 10722
rect 9998 10558 10050 10610
rect 12686 10558 12738 10610
rect 13134 10558 13186 10610
rect 21982 10558 22034 10610
rect 22206 10558 22258 10610
rect 24446 10558 24498 10610
rect 25756 10596 25808 10648
rect 25902 10558 25954 10610
rect 26014 10558 26066 10610
rect 27470 10558 27522 10610
rect 28254 10558 28306 10610
rect 30606 10558 30658 10610
rect 31482 10558 31534 10610
rect 32958 10558 33010 10610
rect 33182 10558 33234 10610
rect 36878 10558 36930 10610
rect 37662 10558 37714 10610
rect 10390 10446 10442 10498
rect 30158 10446 30210 10498
rect 9662 10334 9714 10386
rect 12350 10334 12402 10386
rect 25342 10334 25394 10386
rect 31726 10334 31778 10386
rect 33462 10334 33514 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 28086 9998 28138 10050
rect 32566 9998 32618 10050
rect 4958 9886 5010 9938
rect 5798 9886 5850 9938
rect 7870 9886 7922 9938
rect 11510 9886 11562 9938
rect 23774 9886 23826 9938
rect 27134 9886 27186 9938
rect 30550 9886 30602 9938
rect 37158 9886 37210 9938
rect 2270 9774 2322 9826
rect 3054 9774 3106 9826
rect 7086 9774 7138 9826
rect 7422 9774 7474 9826
rect 7982 9759 8034 9811
rect 8206 9774 8258 9826
rect 8990 9774 9042 9826
rect 9102 9774 9154 9826
rect 25678 9774 25730 9826
rect 26462 9774 26514 9826
rect 26686 9774 26738 9826
rect 27022 9759 27074 9811
rect 27582 9774 27634 9826
rect 27806 9774 27858 9826
rect 30942 9774 30994 9826
rect 31614 9774 31666 9826
rect 31390 9718 31442 9770
rect 32062 9774 32114 9826
rect 32286 9774 32338 9826
rect 35422 9774 35474 9826
rect 36206 9774 36258 9826
rect 8710 9662 8762 9714
rect 33518 9662 33570 9714
rect 31726 9606 31778 9658
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4174 9214 4226 9266
rect 27414 9214 27466 9266
rect 7310 9158 7362 9210
rect 10782 9102 10834 9154
rect 7646 9046 7698 9098
rect 25566 9158 25618 9210
rect 34078 9214 34130 9266
rect 13470 9102 13522 9154
rect 33126 9102 33178 9154
rect 4510 8990 4562 9042
rect 7198 8990 7250 9042
rect 7870 8990 7922 9042
rect 9774 9034 9826 9086
rect 10110 8990 10162 9042
rect 10446 8990 10498 9042
rect 10614 8990 10666 9042
rect 10894 8990 10946 9042
rect 11790 8990 11842 9042
rect 12350 9046 12402 9098
rect 13302 9046 13354 9098
rect 12126 8990 12178 9042
rect 12798 8990 12850 9042
rect 13134 8990 13186 9042
rect 13582 8990 13634 9042
rect 19742 8990 19794 9042
rect 19966 9034 20018 9086
rect 25398 9046 25450 9098
rect 25678 8990 25730 9042
rect 32174 8990 32226 9042
rect 32398 8990 32450 9042
rect 33406 8990 33458 9042
rect 33518 8990 33570 9042
rect 33742 8990 33794 9042
rect 9662 8878 9714 8930
rect 12574 8878 12626 8930
rect 20078 8878 20130 8930
rect 20806 8878 20858 8930
rect 26630 8878 26682 8930
rect 11174 8766 11226 8818
rect 32286 8822 32338 8874
rect 13862 8766 13914 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 7534 8430 7586 8482
rect 8206 8430 8258 8482
rect 16326 8318 16378 8370
rect 19182 8318 19234 8370
rect 21646 8318 21698 8370
rect 10670 8206 10722 8258
rect 11006 8191 11058 8243
rect 13470 8206 13522 8258
rect 14142 8206 14194 8258
rect 14758 8206 14810 8258
rect 16494 8206 16546 8258
rect 17278 8206 17330 8258
rect 19742 8206 19794 8258
rect 20078 8167 20130 8219
rect 20302 8206 20354 8258
rect 21310 8206 21362 8258
rect 21758 8167 21810 8219
rect 21982 8206 22034 8258
rect 22318 8206 22370 8258
rect 24222 8206 24274 8258
rect 24446 8206 24498 8258
rect 23942 8094 23994 8146
rect 10894 8038 10946 8090
rect 14254 8038 14306 8090
rect 19742 8038 19794 8090
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 18062 7646 18114 7698
rect 20582 7534 20634 7586
rect 22150 7534 22202 7586
rect 14142 7422 14194 7474
rect 14366 7422 14418 7474
rect 18398 7422 18450 7474
rect 20190 7422 20242 7474
rect 20302 7422 20354 7474
rect 21646 7422 21698 7474
rect 21870 7422 21922 7474
rect 14646 7198 14698 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 21870 6862 21922 6914
rect 22430 6862 22482 6914
rect 8374 6694 8426 6746
rect 7646 6600 7698 6652
rect 7982 6638 8034 6690
rect 12686 6638 12738 6690
rect 13022 6638 13074 6690
rect 14142 6638 14194 6690
rect 14646 6638 14698 6690
rect 30830 6638 30882 6690
rect 30942 6638 30994 6690
rect 31222 6638 31274 6690
rect 31502 6638 31554 6690
rect 31726 6638 31778 6690
rect 32006 6638 32058 6690
rect 8206 6526 8258 6578
rect 20358 6414 20410 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 27190 6078 27242 6130
rect 12126 6022 12178 6074
rect 30774 6078 30826 6130
rect 28478 6022 28530 6074
rect 31838 6022 31890 6074
rect 7758 5854 7810 5906
rect 7870 5854 7922 5906
rect 8150 5854 8202 5906
rect 8430 5854 8482 5906
rect 8654 5854 8706 5906
rect 9774 5854 9826 5906
rect 12014 5854 12066 5906
rect 12462 5893 12514 5945
rect 12686 5854 12738 5906
rect 14142 5854 14194 5906
rect 19742 5854 19794 5906
rect 19966 5854 20018 5906
rect 20470 5854 20522 5906
rect 20750 5854 20802 5906
rect 20862 5854 20914 5906
rect 21086 5854 21138 5906
rect 21310 5854 21362 5906
rect 22430 5854 22482 5906
rect 22542 5854 22594 5906
rect 22822 5854 22874 5906
rect 23550 5854 23602 5906
rect 23774 5854 23826 5906
rect 27582 5898 27634 5950
rect 27918 5854 27970 5906
rect 28254 5854 28306 5906
rect 28590 5881 28642 5933
rect 28926 5854 28978 5906
rect 29486 5854 29538 5906
rect 29598 5854 29650 5906
rect 31054 5854 31106 5906
rect 31502 5893 31554 5945
rect 31726 5854 31778 5906
rect 32958 5854 33010 5906
rect 9606 5686 9658 5738
rect 27470 5742 27522 5794
rect 29878 5742 29930 5794
rect 8934 5630 8986 5682
rect 13806 5630 13858 5682
rect 20078 5686 20130 5738
rect 21590 5630 21642 5682
rect 24054 5630 24106 5682
rect 33294 5630 33346 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 9214 5182 9266 5234
rect 9830 5182 9882 5234
rect 10894 5182 10946 5234
rect 12798 5182 12850 5234
rect 13638 5182 13690 5234
rect 14030 5182 14082 5234
rect 15934 5182 15986 5234
rect 17446 5182 17498 5234
rect 20302 5182 20354 5234
rect 23214 5182 23266 5234
rect 31614 5182 31666 5234
rect 34078 5182 34130 5234
rect 35254 5182 35306 5234
rect 6526 5070 6578 5122
rect 7310 5070 7362 5122
rect 10110 5070 10162 5122
rect 16718 5070 16770 5122
rect 17614 5070 17666 5122
rect 18398 5070 18450 5122
rect 25118 5070 25170 5122
rect 25902 5070 25954 5122
rect 26294 5070 26346 5122
rect 28478 5070 28530 5122
rect 31278 5070 31330 5122
rect 31558 5040 31610 5092
rect 32174 5070 32226 5122
rect 34862 5070 34914 5122
rect 28142 4846 28194 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 7534 4510 7586 4562
rect 16886 4510 16938 4562
rect 24222 4510 24274 4562
rect 29598 4398 29650 4450
rect 7870 4286 7922 4338
rect 20078 4330 20130 4382
rect 20414 4286 20466 4338
rect 23886 4286 23938 4338
rect 26910 4286 26962 4338
rect 27694 4286 27746 4338
rect 30214 4286 30266 4338
rect 19966 4174 20018 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 1792 45200 1904 46000
rect 5600 45200 5712 46000
rect 9408 45200 9520 46000
rect 13216 45200 13328 46000
rect 17024 45200 17136 46000
rect 20832 45200 20944 46000
rect 24640 45200 24752 46000
rect 28448 45200 28560 46000
rect 32256 45200 32368 46000
rect 36064 45200 36176 46000
rect 39872 45200 39984 46000
rect 43680 45200 43792 46000
rect 1820 43708 1876 45200
rect 1708 43652 1876 43708
rect 5628 43708 5684 45200
rect 9436 43708 9492 45200
rect 5628 43652 5796 43708
rect 9436 43652 9604 43708
rect 1708 23268 1764 43652
rect 5012 41972 5068 41982
rect 5740 41972 5796 43652
rect 5012 41970 5796 41972
rect 5012 41918 5014 41970
rect 5066 41918 5742 41970
rect 5794 41918 5796 41970
rect 5012 41916 5796 41918
rect 5012 41906 5068 41916
rect 5740 41906 5796 41916
rect 8820 41972 8876 41982
rect 9548 41972 9604 43652
rect 8820 41970 9604 41972
rect 8820 41918 8822 41970
rect 8874 41918 9550 41970
rect 9602 41918 9604 41970
rect 8820 41916 9604 41918
rect 8820 41906 8876 41916
rect 9548 41906 9604 41916
rect 13244 41860 13300 45200
rect 13244 41794 13300 41804
rect 13468 41997 13524 42009
rect 13468 41945 13470 41997
rect 13522 41945 13524 41997
rect 6076 41748 6132 41758
rect 6076 41746 6244 41748
rect 6076 41694 6078 41746
rect 6130 41694 6244 41746
rect 6076 41692 6244 41694
rect 6076 41682 6132 41692
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 2156 40404 2212 40414
rect 2156 40310 2212 40348
rect 5460 40404 5516 40414
rect 5460 40310 5516 40348
rect 5740 40404 5796 40414
rect 5740 40310 5796 40348
rect 2940 40290 2996 40302
rect 2940 40238 2942 40290
rect 2994 40238 2996 40290
rect 2828 38948 2884 38958
rect 2940 38948 2996 40238
rect 4844 40290 4900 40302
rect 4844 40238 4846 40290
rect 4898 40238 4900 40290
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 2828 38946 2996 38948
rect 2828 38894 2830 38946
rect 2882 38894 2996 38946
rect 2828 38892 2996 38894
rect 3052 39620 3108 39630
rect 2828 38882 2884 38892
rect 2660 38836 2716 38846
rect 2660 38742 2716 38780
rect 3052 38834 3108 39564
rect 4060 39620 4116 39630
rect 3052 38782 3054 38834
rect 3106 38782 3108 38834
rect 3052 38770 3108 38782
rect 3276 38862 3332 38874
rect 3276 38810 3278 38862
rect 3330 38810 3332 38862
rect 3276 38612 3332 38810
rect 3948 38872 4004 38884
rect 3948 38820 3950 38872
rect 4002 38820 4004 38872
rect 3948 38724 4004 38820
rect 3948 38658 4004 38668
rect 3276 38546 3332 38556
rect 3836 38612 3892 38622
rect 3836 37098 3892 38556
rect 3948 38276 4004 38286
rect 4060 38276 4116 39564
rect 4620 39620 4676 39630
rect 4620 39526 4676 39564
rect 4844 39620 4900 40238
rect 5068 40292 5124 40302
rect 5068 39730 5124 40236
rect 5068 39678 5070 39730
rect 5122 39678 5124 39730
rect 5068 39666 5124 39678
rect 4284 38948 4340 38958
rect 4284 38834 4340 38892
rect 4284 38782 4286 38834
rect 4338 38782 4340 38834
rect 4284 38770 4340 38782
rect 4508 38836 4564 38846
rect 4844 38836 4900 39564
rect 4508 38742 4564 38780
rect 4676 38780 4900 38836
rect 4956 39574 5012 39586
rect 4956 39522 4958 39574
rect 5010 39522 5012 39574
rect 4676 38778 4732 38780
rect 4676 38726 4678 38778
rect 4730 38726 4732 38778
rect 3948 38274 4116 38276
rect 3948 38222 3950 38274
rect 4002 38222 4116 38274
rect 3948 38220 4116 38222
rect 4172 38612 4228 38622
rect 3948 38210 4004 38220
rect 3948 37268 4004 37278
rect 3948 37174 4004 37212
rect 3836 37046 3838 37098
rect 3890 37046 3892 37098
rect 4060 37156 4116 37166
rect 4172 37156 4228 38556
rect 4676 38612 4732 38726
rect 4956 38722 5012 39522
rect 5292 38948 5348 38958
rect 4956 38670 4958 38722
rect 5010 38670 5012 38722
rect 4956 38658 5012 38670
rect 5068 38849 5124 38861
rect 5068 38797 5070 38849
rect 5122 38797 5124 38849
rect 5068 38724 5124 38797
rect 4676 38546 4732 38556
rect 5068 38500 5124 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4844 38444 5124 38500
rect 5292 38834 5348 38892
rect 5292 38782 5294 38834
rect 5346 38782 5348 38834
rect 4844 38276 4900 38444
rect 4508 38220 4900 38276
rect 4508 38050 4564 38220
rect 4342 37994 4398 38006
rect 4342 37942 4344 37994
rect 4396 37942 4398 37994
rect 4342 37828 4398 37942
rect 4342 37762 4398 37772
rect 4508 37998 4510 38050
rect 4562 37998 4564 38050
rect 4116 37100 4228 37156
rect 4060 37090 4116 37100
rect 3836 37034 3892 37046
rect 4508 37044 4564 37998
rect 4620 38050 4676 38062
rect 4620 37998 4622 38050
rect 4674 37998 4676 38050
rect 4620 37492 4676 37998
rect 5124 37828 5180 37838
rect 5124 37734 5180 37772
rect 5292 37492 5348 38782
rect 4620 37436 5348 37492
rect 4688 37304 4744 37316
rect 4688 37252 4690 37304
rect 4742 37252 4744 37304
rect 4688 37156 4744 37252
rect 4688 37090 4744 37100
rect 4844 37268 4900 37278
rect 4172 36988 4564 37044
rect 3276 34145 3332 34157
rect 3276 34093 3278 34145
rect 3330 34093 3332 34145
rect 3164 34020 3220 34030
rect 2604 34018 3220 34020
rect 2604 33966 3166 34018
rect 3218 33966 3220 34018
rect 2604 33964 3220 33966
rect 2604 33458 2660 33964
rect 3164 33954 3220 33964
rect 3276 33908 3332 34093
rect 3612 34132 3668 34142
rect 3612 34130 3780 34132
rect 3612 34078 3614 34130
rect 3666 34078 3780 34130
rect 3612 34076 3780 34078
rect 3612 34066 3668 34076
rect 3276 33842 3332 33852
rect 2604 33406 2606 33458
rect 2658 33406 2660 33458
rect 2604 33394 2660 33406
rect 1820 33346 1876 33358
rect 1820 33294 1822 33346
rect 1874 33294 1876 33346
rect 1820 28644 1876 33294
rect 3724 32452 3780 34076
rect 4172 33908 4228 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4732 34130 4788 34142
rect 4732 34078 4734 34130
rect 4786 34078 4788 34130
rect 4732 34020 4788 34078
rect 4172 33842 4228 33852
rect 4284 33964 4788 34020
rect 4284 32564 4340 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 32470 4340 32508
rect 4508 33234 4564 33246
rect 4508 33182 4510 33234
rect 4562 33182 4564 33234
rect 4508 32564 4564 33182
rect 4508 32498 4564 32508
rect 4620 32562 4676 32574
rect 4620 32510 4622 32562
rect 4674 32510 4676 32562
rect 4060 32452 4116 32462
rect 3724 32450 4116 32452
rect 3724 32398 4062 32450
rect 4114 32398 4116 32450
rect 3724 32396 4116 32398
rect 4060 32386 4116 32396
rect 4620 32452 4676 32510
rect 4844 32564 4900 37212
rect 4956 37044 5012 37436
rect 5124 37268 5180 37278
rect 5124 37174 5180 37212
rect 4956 36988 5124 37044
rect 4956 34132 5012 34142
rect 4956 34038 5012 34076
rect 5068 33796 5124 36988
rect 5852 34914 5908 34926
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5628 34132 5684 34142
rect 5236 34020 5292 34030
rect 5236 34018 5460 34020
rect 5236 33966 5238 34018
rect 5290 33966 5460 34018
rect 5236 33964 5460 33966
rect 5236 33954 5292 33964
rect 5068 33740 5236 33796
rect 5180 33684 5236 33740
rect 5180 33628 5348 33684
rect 5124 33460 5180 33470
rect 5180 33404 5236 33460
rect 5124 33366 5236 33404
rect 4956 32564 5012 32574
rect 4844 32562 5012 32564
rect 4844 32510 4958 32562
rect 5010 32510 5012 32562
rect 4844 32508 5012 32510
rect 4676 32396 4900 32452
rect 4620 32386 4676 32396
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 3724 29441 3780 29466
rect 3724 29428 3726 29441
rect 3778 29428 3780 29441
rect 3724 29362 3780 29372
rect 4060 29426 4116 29438
rect 4060 29374 4062 29426
rect 4114 29374 4116 29426
rect 2604 29316 2660 29326
rect 2604 28754 2660 29260
rect 3612 29316 3668 29326
rect 3612 29222 3668 29260
rect 2604 28702 2606 28754
rect 2658 28702 2660 28754
rect 2604 28690 2660 28702
rect 1820 28550 1876 28588
rect 4060 28532 4116 29374
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4508 28642 4564 28654
rect 4508 28590 4510 28642
rect 4562 28590 4564 28642
rect 4060 28476 4452 28532
rect 4060 27972 4116 27982
rect 4396 27972 4452 28476
rect 4508 28420 4564 28590
rect 4508 28354 4564 28364
rect 4844 28084 4900 32396
rect 4956 31220 5012 32508
rect 4956 31154 5012 31164
rect 5180 28654 5236 33366
rect 5292 32788 5348 33628
rect 5404 33460 5460 33964
rect 5404 33394 5460 33404
rect 5516 33796 5572 33806
rect 5292 32722 5348 32732
rect 5404 33236 5460 33246
rect 5404 32562 5460 33180
rect 5404 32510 5406 32562
rect 5458 32510 5460 32562
rect 5404 32498 5460 32510
rect 5124 28644 5236 28654
rect 5180 28588 5236 28644
rect 5124 28550 5236 28588
rect 4620 27972 4676 27982
rect 4396 27970 4676 27972
rect 4396 27918 4622 27970
rect 4674 27918 4676 27970
rect 4396 27916 4676 27918
rect 4060 27858 4116 27916
rect 4620 27906 4676 27916
rect 4060 27806 4062 27858
rect 4114 27806 4116 27858
rect 4060 27794 4116 27806
rect 4284 27858 4340 27870
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 1932 24722 1988 24734
rect 1932 24670 1934 24722
rect 1986 24670 1988 24722
rect 1932 24612 1988 24670
rect 1932 24546 1988 24556
rect 2716 24612 2772 24622
rect 2716 24610 2996 24612
rect 2716 24558 2718 24610
rect 2770 24558 2996 24610
rect 2716 24556 2996 24558
rect 2716 24546 2772 24556
rect 2940 24276 2996 24556
rect 2940 24220 3220 24276
rect 3164 24162 3220 24220
rect 3164 24110 3166 24162
rect 3218 24110 3220 24162
rect 3164 24098 3220 24110
rect 4172 24052 4228 24062
rect 3500 23938 3556 23950
rect 3500 23886 3502 23938
rect 3554 23886 3556 23938
rect 3500 23604 3556 23886
rect 3500 23548 3892 23604
rect 3836 23322 3892 23548
rect 3836 23270 3838 23322
rect 3890 23270 3892 23322
rect 3836 23258 3892 23270
rect 1708 23202 1764 23212
rect 3948 23154 4004 23166
rect 3948 23102 3950 23154
rect 4002 23102 4004 23154
rect 3948 22484 4004 23102
rect 3948 22418 4004 22428
rect 4172 20916 4228 23996
rect 4284 23210 4340 27806
rect 4844 27858 4900 28028
rect 4844 27806 4846 27858
rect 4898 27806 4900 27858
rect 4844 27794 4900 27806
rect 5068 28420 5124 28430
rect 5068 27858 5124 28364
rect 5068 27806 5070 27858
rect 5122 27806 5124 27858
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4620 24724 4676 24734
rect 4620 24630 4676 24668
rect 5068 24388 5124 27806
rect 5180 24622 5236 28550
rect 5516 30884 5572 33740
rect 5628 33346 5684 34076
rect 5852 33684 5908 34862
rect 6076 34858 6132 34870
rect 6076 34806 6078 34858
rect 6130 34806 6132 34858
rect 5964 34145 6020 34157
rect 5964 34093 5966 34145
rect 6018 34093 6020 34145
rect 5964 33796 6020 34093
rect 6076 34018 6132 34806
rect 6076 33966 6078 34018
rect 6130 33966 6132 34018
rect 6076 33954 6132 33966
rect 6188 34020 6244 41692
rect 9884 41746 9940 41758
rect 9884 41694 9886 41746
rect 9938 41694 9940 41746
rect 9324 40964 9380 40974
rect 8876 40962 9380 40964
rect 8876 40910 9326 40962
rect 9378 40910 9380 40962
rect 8876 40908 9380 40910
rect 6636 40404 6692 40414
rect 6524 40292 6580 40302
rect 6524 40198 6580 40236
rect 6412 37828 6468 37838
rect 6300 35698 6356 35710
rect 6300 35646 6302 35698
rect 6354 35646 6356 35698
rect 6300 34746 6356 35646
rect 6300 34694 6302 34746
rect 6354 34694 6356 34746
rect 6300 34682 6356 34694
rect 6412 34916 6468 37772
rect 6188 33954 6244 33964
rect 6412 33796 6468 34860
rect 5964 33740 6356 33796
rect 5852 33628 6076 33684
rect 5628 33294 5630 33346
rect 5682 33294 5684 33346
rect 5628 33124 5684 33294
rect 5628 33058 5684 33068
rect 5740 33346 5796 33358
rect 5740 33294 5742 33346
rect 5794 33294 5796 33346
rect 5740 33012 5796 33294
rect 5852 33348 5908 33628
rect 6020 33570 6076 33628
rect 6020 33518 6022 33570
rect 6074 33518 6076 33570
rect 6020 33506 6076 33518
rect 5852 33282 5908 33292
rect 6300 33346 6356 33740
rect 6412 33730 6468 33740
rect 6524 36484 6580 36494
rect 6636 36484 6692 40348
rect 8428 40402 8484 40414
rect 8428 40350 8430 40402
rect 8482 40350 8484 40402
rect 7756 38948 7812 38958
rect 7756 38854 7812 38892
rect 8092 38836 8148 38846
rect 8092 38742 8148 38780
rect 8428 38836 8484 40350
rect 8764 39508 8820 39518
rect 8764 39414 8820 39452
rect 8428 38770 8484 38780
rect 6524 36482 6692 36484
rect 6524 36430 6526 36482
rect 6578 36430 6692 36482
rect 6524 36428 6692 36430
rect 6860 37156 6916 37166
rect 6524 33572 6580 36428
rect 6636 35924 6692 35934
rect 6636 35830 6692 35868
rect 6860 34692 6916 37100
rect 7308 36482 7364 36494
rect 7308 36430 7310 36482
rect 7362 36430 7364 36482
rect 7308 35924 7364 36430
rect 7308 35858 7364 35868
rect 7028 34916 7084 34926
rect 7028 34822 7084 34860
rect 6860 34636 7028 34692
rect 6524 33506 6580 33516
rect 6804 33908 6860 33918
rect 6804 33570 6860 33852
rect 6804 33518 6806 33570
rect 6858 33518 6860 33570
rect 6804 33506 6860 33518
rect 6300 33294 6302 33346
rect 6354 33294 6356 33346
rect 6300 33012 6356 33294
rect 6412 33460 6468 33470
rect 6412 33348 6468 33404
rect 6524 33348 6580 33358
rect 6972 33348 7028 34636
rect 6412 33346 6580 33348
rect 6412 33294 6526 33346
rect 6578 33294 6580 33346
rect 6412 33292 6580 33294
rect 6524 33282 6580 33292
rect 6748 33292 7028 33348
rect 8764 33348 8820 33358
rect 5740 32956 6356 33012
rect 6524 33124 6580 33134
rect 5180 24612 5292 24622
rect 5180 24556 5236 24612
rect 5236 24518 5292 24556
rect 4476 24332 4740 24342
rect 5068 24332 5236 24388
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23158 4286 23210
rect 4338 23158 4340 23210
rect 4284 22708 4340 23158
rect 4620 24052 4676 24062
rect 4620 23154 4676 23996
rect 4900 24052 4956 24062
rect 4900 23958 4956 23996
rect 4620 23102 4622 23154
rect 4674 23102 4676 23154
rect 4620 23090 4676 23102
rect 5068 23604 5124 23614
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22642 4340 22652
rect 4620 22484 4676 22494
rect 4620 22390 4676 22428
rect 5068 22484 5124 23548
rect 5180 23156 5236 24332
rect 5516 24052 5572 30828
rect 5628 31220 5684 31230
rect 5628 27982 5684 31164
rect 5740 29428 5796 32956
rect 5852 32788 5908 32798
rect 5852 32562 5908 32732
rect 5852 32510 5854 32562
rect 5906 32510 5908 32562
rect 5852 32498 5908 32510
rect 6300 32601 6356 32613
rect 6300 32564 6302 32601
rect 6354 32564 6356 32601
rect 6300 32498 6356 32508
rect 6524 32562 6580 33068
rect 6524 32510 6526 32562
rect 6578 32510 6580 32562
rect 6524 32498 6580 32510
rect 6188 32450 6244 32462
rect 6188 32398 6190 32450
rect 6242 32398 6244 32450
rect 5908 31554 5964 31566
rect 5908 31502 5910 31554
rect 5962 31502 5964 31554
rect 5908 31218 5964 31502
rect 5908 31166 5910 31218
rect 5962 31166 5964 31218
rect 5908 31154 5964 31166
rect 6188 29540 6244 32398
rect 6636 31666 6692 31678
rect 6636 31614 6638 31666
rect 6690 31614 6692 31666
rect 6188 29484 6412 29540
rect 6356 29482 6412 29484
rect 5852 29428 5908 29438
rect 6076 29428 6132 29438
rect 5740 29372 5852 29428
rect 5628 27972 5740 27982
rect 5628 27916 5684 27972
rect 5684 27878 5740 27916
rect 5516 23986 5572 23996
rect 5740 24948 5796 24958
rect 5740 23604 5796 24892
rect 5852 24610 5908 29372
rect 5852 24558 5854 24610
rect 5906 24558 5908 24610
rect 5852 24546 5908 24558
rect 5964 29426 6132 29428
rect 5964 29374 6078 29426
rect 6130 29374 6132 29426
rect 6356 29430 6358 29482
rect 6410 29430 6412 29482
rect 6356 29418 6412 29430
rect 6524 29428 6580 29438
rect 5964 29372 6132 29374
rect 5964 24766 6020 29372
rect 6076 29362 6132 29372
rect 6524 29314 6580 29372
rect 6524 29262 6526 29314
rect 6578 29262 6580 29314
rect 6524 29250 6580 29262
rect 6636 28868 6692 31614
rect 6748 29426 6804 33292
rect 8428 33124 8484 33134
rect 8428 33030 8484 33068
rect 6860 32564 6916 32574
rect 6860 31948 6916 32508
rect 7252 32452 7308 32462
rect 7252 32358 7308 32396
rect 6860 31892 6935 31948
rect 6879 31778 6935 31892
rect 6879 31726 6881 31778
rect 6933 31726 6935 31778
rect 6879 31714 6935 31726
rect 7756 31778 7812 31790
rect 7756 31726 7758 31778
rect 7810 31726 7812 31778
rect 7756 30996 7812 31726
rect 7756 30930 7812 30940
rect 8764 30996 8820 33292
rect 8876 31948 8932 40908
rect 9324 40898 9380 40908
rect 9884 40962 9940 41694
rect 9884 40910 9886 40962
rect 9938 40910 9940 40962
rect 9884 40898 9940 40910
rect 11788 40628 11844 40638
rect 11788 40514 11844 40572
rect 13468 40628 13524 41945
rect 14476 41860 14532 41870
rect 14476 41766 14532 41804
rect 17052 41860 17108 45200
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 17052 41794 17108 41804
rect 17276 41997 17332 42009
rect 17276 41945 17278 41997
rect 17330 41945 17332 41997
rect 13468 40562 13524 40572
rect 11788 40462 11790 40514
rect 11842 40462 11844 40514
rect 11788 40450 11844 40462
rect 15820 40516 15876 40526
rect 9044 40404 9100 40414
rect 9044 39844 9100 40348
rect 13468 40404 13524 40414
rect 13468 40068 13524 40348
rect 14476 40404 14532 40414
rect 14476 40310 14532 40348
rect 13692 40292 13748 40302
rect 13692 40290 13972 40292
rect 13692 40238 13694 40290
rect 13746 40238 13972 40290
rect 13692 40236 13972 40238
rect 13692 40226 13748 40236
rect 13356 40012 13524 40068
rect 9044 39788 9268 39844
rect 9007 39620 9063 39630
rect 9007 39526 9063 39564
rect 9212 37492 9268 39788
rect 9884 39618 9940 39630
rect 9884 39566 9886 39618
rect 9938 39566 9940 39618
rect 9884 39508 9940 39566
rect 12236 39618 12292 39630
rect 12236 39566 12238 39618
rect 12290 39566 12292 39618
rect 10332 39508 10388 39518
rect 9884 39506 10388 39508
rect 9884 39454 10334 39506
rect 10386 39454 10388 39506
rect 9884 39452 10388 39454
rect 9884 38836 9940 38846
rect 9716 37492 9772 37502
rect 9212 37490 9772 37492
rect 9212 37438 9718 37490
rect 9770 37438 9772 37490
rect 9212 37436 9772 37438
rect 9716 37426 9772 37436
rect 9212 36370 9268 36382
rect 9212 36318 9214 36370
rect 9266 36318 9268 36370
rect 9212 33348 9268 36318
rect 9884 36260 9940 38780
rect 10332 38836 10388 39452
rect 10332 38770 10388 38780
rect 10892 39508 10948 39518
rect 10108 36372 10164 36382
rect 10108 36278 10164 36316
rect 10780 36372 10836 36382
rect 9884 36204 9959 36260
rect 9903 35754 9959 36204
rect 9903 35702 9905 35754
rect 9957 35702 9959 35754
rect 9903 35690 9959 35702
rect 10780 35700 10836 36316
rect 10892 35700 10948 39452
rect 12236 39060 12292 39566
rect 12236 38994 12292 39004
rect 13020 39620 13076 39630
rect 13356 39620 13412 40012
rect 13916 39842 13972 40236
rect 13916 39790 13918 39842
rect 13970 39790 13972 39842
rect 13916 39778 13972 39790
rect 15820 39730 15876 40460
rect 17276 40516 17332 41945
rect 18284 41860 18340 41870
rect 18284 41766 18340 41804
rect 20860 41860 20916 45200
rect 20860 41794 20916 41804
rect 21084 41997 21140 42009
rect 21084 41945 21086 41997
rect 21138 41945 21140 41997
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 17276 40450 17332 40460
rect 21084 40514 21140 41945
rect 22092 41860 22148 41870
rect 22092 41766 22148 41804
rect 24668 41860 24724 45200
rect 24668 41794 24724 41804
rect 24892 41997 24948 42009
rect 24892 41945 24894 41997
rect 24946 41945 24948 41997
rect 24892 41188 24948 41945
rect 25900 41860 25956 41870
rect 25900 41766 25956 41804
rect 28476 41860 28532 45200
rect 28476 41794 28532 41804
rect 28700 41997 28756 42009
rect 28700 41945 28702 41997
rect 28754 41945 28756 41997
rect 21084 40462 21086 40514
rect 21138 40462 21140 40514
rect 21084 40450 21140 40462
rect 24556 41132 24948 41188
rect 24556 40514 24612 41132
rect 24556 40462 24558 40514
rect 24610 40462 24612 40514
rect 24556 40450 24612 40462
rect 28700 40514 28756 41945
rect 29708 41860 29764 41870
rect 29708 41766 29764 41804
rect 32284 41860 32340 45200
rect 32284 41794 32340 41804
rect 32508 41997 32564 42009
rect 32508 41945 32510 41997
rect 32562 41945 32564 41997
rect 28700 40462 28702 40514
rect 28754 40462 28756 40514
rect 28700 40450 28756 40462
rect 32396 40516 32452 40526
rect 32508 40516 32564 41945
rect 33516 41860 33572 41870
rect 33516 41766 33572 41804
rect 36092 41860 36148 45200
rect 36092 41794 36148 41804
rect 36316 41997 36372 42009
rect 36316 41945 36318 41997
rect 36370 41945 36372 41997
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 36316 41188 36372 41945
rect 37324 41860 37380 41870
rect 37324 41766 37380 41804
rect 39900 41860 39956 45200
rect 39900 41794 39956 41804
rect 40124 41997 40180 42009
rect 40124 41945 40126 41997
rect 40178 41945 40180 41997
rect 35980 41132 36372 41188
rect 32396 40514 32564 40516
rect 32396 40462 32398 40514
rect 32450 40462 32564 40514
rect 32396 40460 32564 40462
rect 32788 40962 32844 40974
rect 32788 40910 32790 40962
rect 32842 40910 32844 40962
rect 32396 40450 32452 40460
rect 18396 40404 18452 40414
rect 21868 40404 21924 40414
rect 18452 40348 18564 40404
rect 18396 40310 18452 40348
rect 15820 39678 15822 39730
rect 15874 39678 15876 39730
rect 15820 39666 15876 39678
rect 17724 39732 17780 39742
rect 17724 39638 17780 39676
rect 13020 39618 13412 39620
rect 13020 39566 13022 39618
rect 13074 39566 13412 39618
rect 13020 39564 13412 39566
rect 14252 39620 14308 39630
rect 12012 36484 12068 36494
rect 12796 36484 12852 36494
rect 13020 36484 13076 39564
rect 14252 39526 14308 39564
rect 18508 39618 18564 40348
rect 21756 40348 21868 40404
rect 19180 40290 19236 40302
rect 19180 40238 19182 40290
rect 19234 40238 19236 40290
rect 19180 39844 19236 40238
rect 19180 39778 19236 39788
rect 20188 39844 20244 39854
rect 20188 39750 20244 39788
rect 18508 39566 18510 39618
rect 18562 39566 18564 39618
rect 18508 39554 18564 39566
rect 20524 39618 20580 39630
rect 20524 39566 20526 39618
rect 20578 39566 20580 39618
rect 20524 39508 20580 39566
rect 20524 39442 20580 39452
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 16044 39060 16100 39070
rect 16044 38966 16100 39004
rect 13468 38836 13524 38846
rect 13468 38742 13524 38780
rect 16380 38834 16436 38846
rect 16380 38782 16382 38834
rect 16434 38782 16436 38834
rect 13804 38612 13860 38622
rect 11788 36482 12068 36484
rect 11788 36430 12014 36482
rect 12066 36430 12068 36482
rect 11788 36428 12068 36430
rect 11676 35924 11732 35934
rect 11788 35924 11844 36428
rect 12012 36418 12068 36428
rect 12572 36482 13076 36484
rect 12572 36430 12798 36482
rect 12850 36430 13076 36482
rect 12572 36428 13076 36430
rect 13468 38610 13860 38612
rect 13468 38558 13806 38610
rect 13858 38558 13860 38610
rect 13468 38556 13860 38558
rect 11676 35922 11844 35924
rect 11676 35870 11678 35922
rect 11730 35870 11844 35922
rect 11676 35868 11844 35870
rect 11676 35858 11732 35868
rect 10892 35644 11060 35700
rect 10780 35634 10836 35644
rect 9212 33282 9268 33292
rect 9660 35474 9716 35486
rect 9660 35422 9662 35474
rect 9714 35422 9716 35474
rect 9660 31948 9716 35422
rect 11004 35252 11060 35644
rect 10668 35196 11060 35252
rect 12012 35698 12068 35710
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 8876 31892 9044 31948
rect 9660 31892 9828 31948
rect 8764 30930 8820 30940
rect 8148 30212 8204 30222
rect 8316 30212 8372 30222
rect 7980 30210 8316 30212
rect 7980 30158 8150 30210
rect 8202 30158 8316 30210
rect 7980 30156 8316 30158
rect 6748 29374 6750 29426
rect 6802 29374 6804 29426
rect 6748 29362 6804 29374
rect 6972 29428 7028 29438
rect 6972 29334 7028 29372
rect 7252 29204 7308 29214
rect 7252 29202 7700 29204
rect 7252 29150 7254 29202
rect 7306 29150 7700 29202
rect 7252 29148 7700 29150
rect 7252 29138 7308 29148
rect 6636 28802 6692 28812
rect 6300 28756 6356 28766
rect 6132 28084 6188 28094
rect 6132 27990 6188 28028
rect 6300 27298 6356 28700
rect 6300 27246 6302 27298
rect 6354 27246 6356 27298
rect 6300 27234 6356 27246
rect 7420 27076 7476 27086
rect 6543 27018 6599 27030
rect 6543 26966 6545 27018
rect 6597 26966 6599 27018
rect 7420 26982 7476 27020
rect 6543 26404 6599 26966
rect 5964 24714 5966 24766
rect 6018 24714 6020 24766
rect 5740 23210 5796 23548
rect 5964 23380 6020 24714
rect 5404 23156 5460 23166
rect 5180 23154 5460 23156
rect 5180 23102 5406 23154
rect 5458 23102 5460 23154
rect 5740 23158 5742 23210
rect 5794 23158 5796 23210
rect 5740 23146 5796 23158
rect 5852 23324 6020 23380
rect 6076 26348 6599 26404
rect 5180 23100 5460 23102
rect 4844 22372 4900 22382
rect 4788 22316 4844 22326
rect 4788 22314 4900 22316
rect 4788 22262 4790 22314
rect 4842 22262 4900 22314
rect 5068 22370 5124 22428
rect 5068 22318 5070 22370
rect 5122 22318 5124 22370
rect 5068 22306 5124 22318
rect 4788 22204 4900 22262
rect 4844 21924 4900 22204
rect 4844 21868 5124 21924
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4620 20916 4676 20926
rect 4172 20860 4452 20916
rect 4284 20188 4340 20198
rect 3500 20186 4340 20188
rect 3500 20134 4286 20186
rect 4338 20134 4340 20186
rect 3500 20132 4340 20134
rect 3500 20018 3556 20132
rect 4284 20122 4340 20132
rect 3500 19966 3502 20018
rect 3554 19966 3556 20018
rect 3500 19954 3556 19966
rect 4284 20020 4340 20030
rect 4396 20020 4452 20860
rect 4340 19964 4452 20020
rect 4620 20074 4676 20860
rect 5068 20188 5124 21868
rect 5404 21812 5460 23100
rect 5628 23044 5684 23054
rect 5852 23044 5908 23324
rect 5628 23042 5908 23044
rect 5628 22990 5630 23042
rect 5682 22990 5908 23042
rect 5628 22988 5908 22990
rect 5964 23156 6020 23166
rect 6076 23156 6132 26348
rect 6748 24948 6804 24958
rect 6748 24854 6804 24892
rect 6300 24724 6356 24734
rect 7084 24724 7140 24734
rect 6300 24722 6468 24724
rect 6300 24670 6302 24722
rect 6354 24670 6468 24722
rect 6300 24668 6468 24670
rect 6300 24658 6356 24668
rect 6300 23156 6356 23166
rect 5964 23154 6132 23156
rect 5964 23102 5966 23154
rect 6018 23102 6132 23154
rect 5964 23100 6132 23102
rect 6188 23154 6356 23156
rect 6188 23102 6302 23154
rect 6354 23102 6356 23154
rect 6188 23100 6356 23102
rect 5628 22978 5684 22988
rect 5684 22596 5740 22606
rect 5964 22596 6020 23100
rect 5684 22502 5740 22540
rect 5852 22540 6020 22596
rect 5404 21746 5460 21756
rect 5628 20916 5684 20926
rect 5628 20822 5684 20860
rect 5852 20804 5908 22540
rect 6076 22484 6132 22494
rect 5964 22372 6020 22382
rect 5964 22278 6020 22316
rect 6076 22370 6132 22428
rect 6076 22318 6078 22370
rect 6130 22318 6132 22370
rect 6076 22306 6132 22318
rect 5964 20804 6020 20814
rect 5852 20802 6132 20804
rect 4620 20022 4622 20074
rect 4674 20022 4676 20074
rect 4620 20010 4676 20022
rect 4844 20132 5124 20188
rect 5740 20758 5796 20770
rect 5740 20706 5742 20758
rect 5794 20706 5796 20758
rect 5852 20750 5966 20802
rect 6018 20750 6132 20802
rect 5852 20748 6132 20750
rect 5964 20738 6020 20748
rect 4844 20018 4900 20132
rect 4844 19966 4846 20018
rect 4898 19966 4900 20018
rect 4284 19926 4340 19964
rect 3164 19796 3220 19806
rect 2604 19794 3220 19796
rect 2604 19742 3166 19794
rect 3218 19742 3220 19794
rect 2604 19740 3220 19742
rect 2604 19346 2660 19740
rect 3164 19730 3220 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4844 19460 4900 19966
rect 5572 20020 5628 20030
rect 5572 19926 5628 19964
rect 4844 19394 4900 19404
rect 2604 19294 2606 19346
rect 2658 19294 2660 19346
rect 2604 19282 2660 19294
rect 4508 19348 4564 19358
rect 4508 19254 4564 19292
rect 1820 19236 1876 19246
rect 5124 19236 5180 19246
rect 1820 19142 1876 19180
rect 5068 19180 5124 19236
rect 5068 19142 5180 19180
rect 5740 19236 5796 20706
rect 6076 20132 6132 20748
rect 6076 20066 6132 20076
rect 6188 20020 6244 23100
rect 6300 23090 6356 23100
rect 6412 22260 6468 24668
rect 7084 24630 7140 24668
rect 6412 22194 6468 22204
rect 6188 19926 6244 19964
rect 6300 20132 6356 20142
rect 6300 20018 6356 20076
rect 6300 19966 6302 20018
rect 6354 19966 6356 20018
rect 5908 19796 5964 19806
rect 5908 19794 6244 19796
rect 5908 19742 5910 19794
rect 5962 19742 6244 19794
rect 5908 19740 6244 19742
rect 5908 19730 5964 19740
rect 5908 19460 5964 19470
rect 5908 19366 5964 19404
rect 5740 19170 5796 19180
rect 6188 19234 6244 19740
rect 6300 19348 6356 19966
rect 6300 19282 6356 19292
rect 7196 20020 7252 20030
rect 7196 19460 7252 19964
rect 6188 19182 6190 19234
rect 6242 19182 6244 19234
rect 6188 19170 6244 19182
rect 6412 19234 6468 19246
rect 6412 19182 6414 19234
rect 6466 19182 6468 19234
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4508 15316 4564 15326
rect 4508 15222 4564 15260
rect 5068 15316 5124 19142
rect 6412 19012 6468 19182
rect 6692 19236 6748 19246
rect 6692 19142 6748 19180
rect 6972 19234 7028 19246
rect 6972 19182 6974 19234
rect 7026 19182 7028 19234
rect 6412 18946 6468 18956
rect 6972 19012 7028 19182
rect 7196 19234 7252 19404
rect 7196 19182 7198 19234
rect 7250 19182 7252 19234
rect 7196 19170 7252 19182
rect 6972 18946 7028 18956
rect 7644 18340 7700 29148
rect 7756 28756 7812 28766
rect 7756 28642 7812 28700
rect 7756 28590 7758 28642
rect 7810 28590 7812 28642
rect 7756 28578 7812 28590
rect 7980 28644 8036 30156
rect 8148 30146 8204 30156
rect 8316 30118 8372 30156
rect 7980 28578 8036 28588
rect 8092 28868 8148 28878
rect 8092 28642 8148 28812
rect 8092 28590 8094 28642
rect 8146 28590 8148 28642
rect 8092 28578 8148 28590
rect 8204 28810 8260 28822
rect 8204 28758 8206 28810
rect 8258 28758 8260 28810
rect 8204 28308 8260 28758
rect 8204 28242 8260 28252
rect 7980 24612 8036 24622
rect 7980 22372 8036 24556
rect 8988 24052 9044 31892
rect 9436 30212 9492 30222
rect 9436 30118 9492 30156
rect 9772 28644 9828 31892
rect 9884 31668 9940 31678
rect 9884 31666 10052 31668
rect 9884 31614 9886 31666
rect 9938 31614 10052 31666
rect 9884 31612 10052 31614
rect 9884 31602 9940 31612
rect 9996 31044 10052 31612
rect 10668 31220 10724 35196
rect 12012 34244 12068 35646
rect 12012 34178 12068 34188
rect 11788 31780 11844 31790
rect 12572 31780 12628 36428
rect 12796 36418 12852 36428
rect 13356 35700 13412 35710
rect 13468 35700 13524 38556
rect 13804 38546 13860 38556
rect 16380 37156 16436 38782
rect 17500 37826 17556 37838
rect 17500 37774 17502 37826
rect 17554 37774 17556 37826
rect 16380 37090 16436 37100
rect 17388 37266 17444 37278
rect 17388 37214 17390 37266
rect 17442 37214 17444 37266
rect 13356 35698 13524 35700
rect 13356 35646 13358 35698
rect 13410 35646 13524 35698
rect 13356 35644 13524 35646
rect 13356 35634 13412 35644
rect 13468 35588 13524 35644
rect 13916 35700 13972 35710
rect 13916 35606 13972 35644
rect 14364 35700 14420 35710
rect 14364 35606 14420 35644
rect 16380 35700 16436 35710
rect 16044 35588 16100 35598
rect 13468 35522 13524 35532
rect 14140 35530 14196 35542
rect 14140 35478 14142 35530
rect 14194 35478 14196 35530
rect 14140 35140 14196 35478
rect 14700 35474 14756 35486
rect 14700 35422 14702 35474
rect 14754 35422 14756 35474
rect 14700 35364 14756 35422
rect 14700 35298 14756 35308
rect 14140 35084 14644 35140
rect 14383 34858 14439 34870
rect 14140 34804 14196 34814
rect 14383 34806 14385 34858
rect 14437 34806 14439 34858
rect 14140 34802 14308 34804
rect 14140 34750 14142 34802
rect 14194 34750 14308 34802
rect 14140 34748 14308 34750
rect 14140 34738 14196 34748
rect 13860 34244 13916 34254
rect 14252 34244 14308 34748
rect 14383 34468 14439 34806
rect 14383 34402 14439 34412
rect 14588 34356 14644 35084
rect 15260 34916 15316 34926
rect 15260 34822 15316 34860
rect 14476 34300 14644 34356
rect 14700 34580 14756 34590
rect 14252 34188 14364 34244
rect 13860 34150 13916 34188
rect 14308 34186 14364 34188
rect 14140 34158 14196 34170
rect 11788 31778 12180 31780
rect 11788 31726 11790 31778
rect 11842 31726 12180 31778
rect 11788 31724 12180 31726
rect 11788 31714 11844 31724
rect 11676 31220 11732 31230
rect 10668 31164 11396 31220
rect 9992 31032 10052 31044
rect 9992 30980 9994 31032
rect 10046 30980 10052 31032
rect 9992 30940 10052 30980
rect 10108 30996 10164 31006
rect 9992 30772 10048 30940
rect 9992 30706 10048 30716
rect 10108 29988 10164 30940
rect 10668 30996 10724 31006
rect 10668 30902 10724 30940
rect 10104 29932 10164 29988
rect 10780 30826 10836 30838
rect 10780 30774 10782 30826
rect 10834 30774 10836 30826
rect 10104 29464 10160 29932
rect 10780 29764 10836 30774
rect 10780 29708 11172 29764
rect 10104 29412 10106 29464
rect 10158 29412 10160 29464
rect 10104 29400 10160 29412
rect 10780 29428 10836 29438
rect 10780 29334 10836 29372
rect 10556 29258 10612 29270
rect 10556 29206 10558 29258
rect 10610 29206 10612 29258
rect 10556 28812 10612 29206
rect 10220 28756 10276 28766
rect 9996 28754 10276 28756
rect 9996 28702 10222 28754
rect 10274 28702 10276 28754
rect 9996 28700 10276 28702
rect 9884 28644 9940 28654
rect 9772 28642 9940 28644
rect 9772 28590 9886 28642
rect 9938 28590 9940 28642
rect 9772 28588 9940 28590
rect 9884 28578 9940 28588
rect 9324 28084 9380 28094
rect 9324 25674 9380 28028
rect 9996 27858 10052 28700
rect 10220 28690 10276 28700
rect 10332 28756 10612 28812
rect 10332 28598 10388 28756
rect 11004 28754 11060 28766
rect 11004 28702 11006 28754
rect 11058 28702 11060 28754
rect 10276 28586 10388 28598
rect 10276 28534 10278 28586
rect 10330 28534 10388 28586
rect 10276 28476 10388 28534
rect 10444 28642 10500 28654
rect 10444 28590 10446 28642
rect 10498 28590 10500 28642
rect 10332 28308 10388 28318
rect 9996 27806 9998 27858
rect 10050 27806 10052 27858
rect 9996 27794 10052 27806
rect 10108 28026 10164 28038
rect 10108 27974 10110 28026
rect 10162 27974 10164 28026
rect 9544 26328 9600 26340
rect 9544 26276 9546 26328
rect 9598 26276 9600 26328
rect 9544 25844 9600 26276
rect 9996 26292 10052 26302
rect 9544 25788 9604 25844
rect 9324 25622 9326 25674
rect 9378 25622 9380 25674
rect 9324 25610 9380 25622
rect 9324 25506 9380 25518
rect 9324 25454 9326 25506
rect 9378 25454 9380 25506
rect 9324 24948 9380 25454
rect 9324 24882 9380 24892
rect 9548 24724 9604 25788
rect 9996 25518 10052 26236
rect 10108 25620 10164 27974
rect 10332 27914 10388 28252
rect 10332 27862 10334 27914
rect 10386 27862 10388 27914
rect 10332 27850 10388 27862
rect 10444 27412 10500 28590
rect 10892 28642 10948 28654
rect 10892 28590 10894 28642
rect 10946 28590 10948 28642
rect 10892 28084 10948 28590
rect 10892 28018 10948 28028
rect 10668 27860 10724 27870
rect 11004 27860 11060 28702
rect 11116 28644 11172 29708
rect 11340 28644 11396 31164
rect 11676 30996 11732 31164
rect 11676 30902 11732 30940
rect 12124 30434 12180 31724
rect 14140 34106 14142 34158
rect 14194 34106 14196 34158
rect 14308 34134 14310 34186
rect 14362 34134 14364 34186
rect 14308 34122 14364 34134
rect 12572 31686 12628 31724
rect 13804 31750 13860 31762
rect 13804 31698 13806 31750
rect 13858 31698 13860 31750
rect 13804 31668 13860 31698
rect 12124 30382 12126 30434
rect 12178 30382 12180 30434
rect 12124 30370 12180 30382
rect 12236 30994 12292 31006
rect 12236 30942 12238 30994
rect 12290 30942 12292 30994
rect 12236 30772 12292 30942
rect 11676 30212 11732 30222
rect 11676 30130 11678 30156
rect 11730 30130 11732 30156
rect 11676 30118 11732 30130
rect 11564 29428 11620 29438
rect 11564 29334 11620 29372
rect 11900 29428 11956 29438
rect 12236 29428 12292 30716
rect 12460 30826 12516 30838
rect 12460 30774 12462 30826
rect 12514 30774 12516 30826
rect 12460 30436 12516 30774
rect 12460 30380 12628 30436
rect 12460 30210 12516 30222
rect 12460 30158 12462 30210
rect 12514 30158 12516 30210
rect 12460 30100 12516 30158
rect 12460 30034 12516 30044
rect 11900 29426 12292 29428
rect 11900 29374 11902 29426
rect 11954 29374 12292 29426
rect 11900 29372 12292 29374
rect 11900 29362 11956 29372
rect 11564 28644 11620 28654
rect 11116 28588 11228 28644
rect 11340 28642 11620 28644
rect 11340 28590 11566 28642
rect 11618 28590 11620 28642
rect 11340 28588 11620 28590
rect 11172 28586 11228 28588
rect 11172 28534 11174 28586
rect 11226 28534 11228 28586
rect 11564 28578 11620 28588
rect 12572 28644 12628 30380
rect 12852 30212 12908 30222
rect 12852 30118 12908 30156
rect 13804 30212 13860 31612
rect 13804 30146 13860 30156
rect 14140 29876 14196 34106
rect 14476 31948 14532 34300
rect 14700 34186 14756 34524
rect 14588 34158 14644 34170
rect 14588 34106 14590 34158
rect 14642 34106 14644 34158
rect 14700 34134 14702 34186
rect 14754 34134 14756 34186
rect 14700 34122 14756 34134
rect 16044 34130 16100 35532
rect 16268 34916 16324 34926
rect 16268 34692 16324 34860
rect 14588 34020 14644 34106
rect 16044 34078 16046 34130
rect 16098 34078 16100 34130
rect 16212 34636 16324 34692
rect 16212 34186 16268 34636
rect 16212 34134 16214 34186
rect 16266 34134 16268 34186
rect 16212 34122 16268 34134
rect 16380 34130 16436 35644
rect 16604 35588 16660 35598
rect 16604 34914 16660 35532
rect 17388 35588 17444 37214
rect 17500 37266 17556 37774
rect 18396 37826 18452 37838
rect 18396 37774 18398 37826
rect 18450 37774 18452 37826
rect 17500 37214 17502 37266
rect 17554 37214 17556 37266
rect 17500 37202 17556 37214
rect 17646 37303 17702 37315
rect 17646 37251 17648 37303
rect 17700 37251 17702 37303
rect 17646 36820 17702 37251
rect 18060 37156 18116 37166
rect 18060 37062 18116 37100
rect 17388 35522 17444 35532
rect 17500 36764 17702 36820
rect 16940 35028 16996 35038
rect 16940 35026 17108 35028
rect 16940 34974 16942 35026
rect 16994 34974 17108 35026
rect 16940 34972 17108 34974
rect 16940 34962 16996 34972
rect 16604 34862 16606 34914
rect 16658 34862 16660 34914
rect 16604 34850 16660 34862
rect 16940 34858 16996 34870
rect 16940 34806 16942 34858
rect 16994 34806 16996 34858
rect 16940 34804 16996 34806
rect 16940 34738 16996 34748
rect 16044 34066 16100 34078
rect 16380 34078 16382 34130
rect 16434 34078 16436 34130
rect 15204 34020 15260 34030
rect 14588 34018 15260 34020
rect 14588 33966 15206 34018
rect 15258 33966 15260 34018
rect 14588 33964 15260 33966
rect 12572 28578 12628 28588
rect 13468 28980 13524 28990
rect 11172 28522 11228 28534
rect 10668 27858 11060 27860
rect 10668 27806 10670 27858
rect 10722 27806 11060 27858
rect 10668 27804 11060 27806
rect 10668 27794 10724 27804
rect 10332 27356 10500 27412
rect 10220 26290 10276 26302
rect 10220 26238 10222 26290
rect 10274 26238 10276 26290
rect 10220 25844 10276 26238
rect 10332 26122 10388 27356
rect 10332 26070 10334 26122
rect 10386 26070 10388 26122
rect 10332 26058 10388 26070
rect 10220 25788 10724 25844
rect 10668 25732 10724 25788
rect 10668 25638 10724 25676
rect 10108 25564 10276 25620
rect 9996 25508 10056 25518
rect 9996 25452 10000 25508
rect 10000 25416 10002 25452
rect 10054 25416 10056 25452
rect 10000 25404 10056 25416
rect 9548 24658 9604 24668
rect 8988 23986 9044 23996
rect 10108 23940 10164 23950
rect 10108 23846 10164 23884
rect 9772 23716 9828 23726
rect 8764 23714 9828 23716
rect 8764 23662 9774 23714
rect 9826 23662 9828 23714
rect 8764 23660 9828 23662
rect 8764 22482 8820 23660
rect 9772 23650 9828 23660
rect 10220 22596 10276 25564
rect 10332 25508 10388 25518
rect 10332 25414 10388 25452
rect 11900 25172 11956 25182
rect 11900 24162 11956 25116
rect 13468 24836 13524 28924
rect 14140 28980 14196 29820
rect 14140 28914 14196 28924
rect 14364 31892 14532 31948
rect 15036 32452 15092 33964
rect 15204 33954 15260 33964
rect 16380 33908 16436 34078
rect 13692 28644 13748 28654
rect 13692 27858 13748 28588
rect 13692 27806 13694 27858
rect 13746 27806 13748 27858
rect 13692 27794 13748 27806
rect 14028 27885 14084 27897
rect 14028 27833 14030 27885
rect 14082 27833 14084 27885
rect 13916 27748 13972 27758
rect 13916 27654 13972 27692
rect 13916 26305 13972 26330
rect 13580 26290 13636 26302
rect 13580 26238 13582 26290
rect 13634 26238 13636 26290
rect 13580 25508 13636 26238
rect 13916 26292 13918 26305
rect 13970 26292 13972 26305
rect 13916 26226 13972 26236
rect 14028 26178 14084 27833
rect 14364 27858 14420 31892
rect 14812 31780 14868 31790
rect 14812 31556 14868 31724
rect 14812 31554 14980 31556
rect 14812 31502 14814 31554
rect 14866 31502 14980 31554
rect 14812 31500 14980 31502
rect 14812 31490 14868 31500
rect 14924 31021 14980 31500
rect 14924 30969 14926 31021
rect 14978 30969 14980 31021
rect 14924 30957 14980 30969
rect 14924 30210 14980 30222
rect 14924 30158 14926 30210
rect 14978 30158 14980 30210
rect 14924 29316 14980 30158
rect 14364 27806 14366 27858
rect 14418 27806 14420 27858
rect 14364 27794 14420 27806
rect 14700 27858 14756 27870
rect 14700 27806 14702 27858
rect 14754 27806 14756 27858
rect 14700 27188 14756 27806
rect 14812 27188 14868 27198
rect 14700 27186 14868 27188
rect 14700 27134 14814 27186
rect 14866 27134 14868 27186
rect 14700 27132 14868 27134
rect 14812 27122 14868 27132
rect 14364 27076 14420 27086
rect 14364 26982 14420 27020
rect 14700 27030 14756 27042
rect 14700 26978 14702 27030
rect 14754 26978 14756 27030
rect 14700 26964 14756 26978
rect 14700 26898 14756 26908
rect 14588 26292 14644 26302
rect 14028 26126 14030 26178
rect 14082 26126 14084 26178
rect 14028 26114 14084 26126
rect 14476 26290 14644 26292
rect 14476 26238 14590 26290
rect 14642 26238 14644 26290
rect 14476 26236 14644 26238
rect 13804 25508 13860 25518
rect 13580 25506 13860 25508
rect 13580 25454 13806 25506
rect 13858 25454 13860 25506
rect 13580 25452 13860 25454
rect 13804 25172 13860 25452
rect 14476 25284 14532 26236
rect 14588 26226 14644 26236
rect 14924 25844 14980 29260
rect 14924 25778 14980 25788
rect 14680 25508 14736 25518
rect 14680 25414 14736 25452
rect 14476 25218 14532 25228
rect 14924 25394 14980 25406
rect 14924 25342 14926 25394
rect 14978 25342 14980 25394
rect 14924 25172 14980 25342
rect 13804 25106 13860 25116
rect 14588 25116 14980 25172
rect 14588 25060 14644 25116
rect 14252 25004 14644 25060
rect 13468 24780 14028 24836
rect 13972 24778 14028 24780
rect 13972 24726 13974 24778
rect 14026 24726 14028 24778
rect 13972 24714 14028 24726
rect 14252 24778 14308 25004
rect 15036 24958 15092 32396
rect 16044 33852 16436 33908
rect 16492 34130 16548 34142
rect 16492 34078 16494 34130
rect 16546 34078 16548 34130
rect 15484 31780 15540 31790
rect 15372 30154 15428 30166
rect 15148 30100 15204 30110
rect 15148 30042 15204 30044
rect 15148 29990 15150 30042
rect 15202 29990 15204 30042
rect 15372 30102 15374 30154
rect 15426 30102 15428 30154
rect 15372 30100 15428 30102
rect 15372 30034 15428 30044
rect 15148 29978 15204 29990
rect 15484 29467 15540 31724
rect 16044 30996 16100 33852
rect 16212 32450 16268 32462
rect 16212 32398 16214 32450
rect 16266 32398 16268 32450
rect 16212 31948 16268 32398
rect 16492 31948 16548 34078
rect 16772 34132 16828 34142
rect 16772 34038 16828 34076
rect 17052 34020 17108 34972
rect 17276 34916 17332 34926
rect 17276 34822 17332 34860
rect 17500 34254 17556 36764
rect 18396 36270 18452 37774
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 21756 37502 21812 40348
rect 21868 40310 21924 40348
rect 25396 40404 25452 40414
rect 25396 40310 25452 40348
rect 26012 40404 26068 40414
rect 26012 40310 26068 40348
rect 28588 40404 28644 40414
rect 22652 40290 22708 40302
rect 26796 40292 26852 40302
rect 22652 40238 22654 40290
rect 22706 40238 22708 40290
rect 22652 39844 22708 40238
rect 26684 40290 26852 40292
rect 26684 40238 26798 40290
rect 26850 40238 26852 40290
rect 26684 40236 26852 40238
rect 24444 39844 24500 39854
rect 22652 39778 22708 39788
rect 23660 39786 23716 39798
rect 23660 39734 23662 39786
rect 23714 39734 23716 39786
rect 24444 39750 24500 39788
rect 23660 39732 23716 39734
rect 23660 39666 23716 39676
rect 23436 39620 23492 39630
rect 23436 38274 23492 39564
rect 23548 39618 23604 39630
rect 23548 39566 23550 39618
rect 23602 39566 23604 39618
rect 23548 38836 23604 39566
rect 23772 39618 23828 39630
rect 24108 39620 24164 39630
rect 23772 39566 23774 39618
rect 23826 39566 23828 39618
rect 23772 38948 23828 39566
rect 23548 38770 23604 38780
rect 23660 38892 23828 38948
rect 23884 39618 24164 39620
rect 23884 39566 24110 39618
rect 24162 39566 24164 39618
rect 23884 39564 24164 39566
rect 23436 38222 23438 38274
rect 23490 38222 23492 38274
rect 23436 38210 23492 38222
rect 23660 37940 23716 38892
rect 23772 38724 23828 38734
rect 23884 38724 23940 39564
rect 24108 39554 24164 39564
rect 23772 38722 23940 38724
rect 23772 38670 23774 38722
rect 23826 38670 23940 38722
rect 23772 38668 23940 38670
rect 24166 38834 24222 38846
rect 24166 38782 24168 38834
rect 24220 38782 24222 38834
rect 23772 38658 23828 38668
rect 24166 38276 24222 38782
rect 24332 38836 24388 38846
rect 24332 38742 24388 38780
rect 24444 38834 24500 38846
rect 24444 38782 24446 38834
rect 24498 38782 24500 38834
rect 23884 38220 24222 38276
rect 24444 38276 24500 38782
rect 23884 38062 23940 38220
rect 24444 38210 24500 38220
rect 23660 37874 23716 37884
rect 23830 38050 23940 38062
rect 23830 37998 23832 38050
rect 23884 37998 23940 38050
rect 23830 37996 23940 37998
rect 23996 38050 24052 38062
rect 23996 37998 23998 38050
rect 24050 37998 24052 38050
rect 23830 37828 23886 37996
rect 23996 37940 24052 37998
rect 24108 38052 24164 38062
rect 24108 38050 24612 38052
rect 24108 37998 24110 38050
rect 24162 37998 24612 38050
rect 24108 37996 24612 37998
rect 24108 37986 24164 37996
rect 23996 37874 24052 37884
rect 23830 37762 23886 37772
rect 21700 37492 21812 37502
rect 21308 37490 21812 37492
rect 21308 37438 21702 37490
rect 21754 37438 21812 37490
rect 21308 37436 21812 37438
rect 21308 37266 21364 37436
rect 21700 37426 21756 37436
rect 21308 37214 21310 37266
rect 21362 37214 21364 37266
rect 21308 37202 21364 37214
rect 18620 37154 18676 37166
rect 18620 37102 18622 37154
rect 18674 37102 18676 37154
rect 18396 36258 18508 36270
rect 18396 36206 18454 36258
rect 18506 36206 18508 36258
rect 18396 36204 18508 36206
rect 18452 35924 18508 36204
rect 18284 35868 18508 35924
rect 17612 34914 17668 34926
rect 17612 34862 17614 34914
rect 17666 34862 17668 34914
rect 17612 34468 17668 34862
rect 17612 34402 17668 34412
rect 18004 34692 18060 34702
rect 17444 34242 17556 34254
rect 17444 34190 17446 34242
rect 17498 34190 17556 34242
rect 17444 34188 17556 34190
rect 17444 34178 17500 34188
rect 17724 34132 17780 34142
rect 17612 34130 17780 34132
rect 17612 34078 17726 34130
rect 17778 34078 17780 34130
rect 17612 34076 17780 34078
rect 17612 34020 17668 34076
rect 17724 34066 17780 34076
rect 17836 34132 17892 34142
rect 17836 34038 17892 34076
rect 18004 34074 18060 34636
rect 18284 34356 18340 35868
rect 18396 35700 18452 35710
rect 18620 35700 18676 37102
rect 20524 37154 20580 37166
rect 20524 37102 20526 37154
rect 20578 37102 20580 37154
rect 20524 37044 20580 37102
rect 20524 36978 20580 36988
rect 19516 36932 19572 36942
rect 19516 36706 19572 36876
rect 19516 36654 19518 36706
rect 19570 36654 19572 36706
rect 19516 36642 19572 36654
rect 18452 35644 18676 35700
rect 19180 36482 19236 36494
rect 19180 36430 19182 36482
rect 19234 36430 19236 36482
rect 18396 35606 18452 35644
rect 18732 35476 18788 35486
rect 18508 35474 18788 35476
rect 18508 35422 18734 35474
rect 18786 35422 18788 35474
rect 18508 35420 18788 35422
rect 18508 35140 18564 35420
rect 18732 35410 18788 35420
rect 18284 34290 18340 34300
rect 18396 35084 18564 35140
rect 19180 35150 19236 36430
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19180 35138 19292 35150
rect 19180 35086 19238 35138
rect 19290 35086 19292 35138
rect 19180 35084 19292 35086
rect 18396 34916 18452 35084
rect 19236 35074 19292 35084
rect 17052 33964 17668 34020
rect 18004 34022 18006 34074
rect 18058 34022 18060 34074
rect 18172 34132 18228 34142
rect 18396 34132 18452 34860
rect 18172 34130 18340 34132
rect 18172 34078 18174 34130
rect 18226 34078 18340 34130
rect 18172 34076 18340 34078
rect 18172 34066 18228 34076
rect 18004 33684 18060 34022
rect 17948 33628 18060 33684
rect 18172 33796 18228 33806
rect 16212 31892 16324 31948
rect 16492 31902 16660 31948
rect 16492 31892 16716 31902
rect 16156 31778 16212 31790
rect 16156 31726 16158 31778
rect 16210 31726 16212 31778
rect 16156 31556 16212 31726
rect 16156 31490 16212 31500
rect 16268 31668 16324 31892
rect 16604 31890 16716 31892
rect 16604 31838 16662 31890
rect 16714 31838 16716 31890
rect 16604 31836 16716 31838
rect 16380 31780 16436 31790
rect 16380 31686 16436 31724
rect 16660 31780 16716 31836
rect 16660 31714 16716 31724
rect 17164 31780 17220 31790
rect 17164 31686 17220 31724
rect 16268 31220 16324 31612
rect 16716 31556 16772 31566
rect 16268 31164 16436 31220
rect 16044 30930 16100 30940
rect 16268 30996 16324 31006
rect 16268 30902 16324 30940
rect 16156 30884 16212 30894
rect 16156 30826 16212 30828
rect 16156 30774 16158 30826
rect 16210 30774 16212 30826
rect 16156 30762 16212 30774
rect 16380 30324 16436 31164
rect 16604 30994 16660 31006
rect 16604 30942 16606 30994
rect 16658 30942 16660 30994
rect 16604 30772 16660 30942
rect 16604 30706 16660 30716
rect 16380 30258 16436 30268
rect 15596 30212 15652 30222
rect 15596 30210 15764 30212
rect 15596 30158 15598 30210
rect 15650 30158 15764 30210
rect 16716 30210 16772 31500
rect 17500 31556 17556 31566
rect 17500 31462 17556 31500
rect 17948 31220 18004 33628
rect 18060 33460 18116 33470
rect 18060 31556 18116 33404
rect 18172 33346 18228 33740
rect 18284 33572 18340 34076
rect 18396 33796 18452 34076
rect 18396 33730 18452 33740
rect 18508 34914 18564 34926
rect 18508 34862 18510 34914
rect 18562 34862 18564 34914
rect 18956 34914 19012 34926
rect 18508 33572 18564 34862
rect 18676 34858 18732 34870
rect 18676 34806 18678 34858
rect 18730 34806 18732 34858
rect 18956 34862 18958 34914
rect 19010 34862 19012 34914
rect 18676 34692 18732 34806
rect 18676 34626 18732 34636
rect 18844 34802 18900 34814
rect 18844 34750 18846 34802
rect 18898 34750 18900 34802
rect 18620 34468 18676 34478
rect 18620 34130 18676 34412
rect 18844 34254 18900 34750
rect 18956 34580 19012 34862
rect 23660 34916 23716 34926
rect 18956 34514 19012 34524
rect 19292 34580 19348 34590
rect 18844 34242 18956 34254
rect 18844 34190 18902 34242
rect 18954 34190 18956 34242
rect 18844 34188 18956 34190
rect 18900 34178 18956 34188
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18620 33796 18676 34078
rect 19292 33962 19348 34524
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 23660 34354 23716 34860
rect 23660 34302 23662 34354
rect 23714 34302 23716 34354
rect 19292 33910 19294 33962
rect 19346 33910 19348 33962
rect 19292 33898 19348 33910
rect 19404 34130 19460 34142
rect 19404 34078 19406 34130
rect 19458 34078 19460 34130
rect 18620 33730 18676 33740
rect 19404 33796 19460 34078
rect 19628 34132 19684 34142
rect 19628 34038 19684 34076
rect 21980 34130 22036 34142
rect 21980 34078 21982 34130
rect 22034 34078 22036 34130
rect 19404 33730 19460 33740
rect 20244 34018 20300 34030
rect 20244 33966 20246 34018
rect 20298 33966 20300 34018
rect 18844 33572 18900 33582
rect 18284 33516 18452 33572
rect 18508 33570 18900 33572
rect 18508 33518 18846 33570
rect 18898 33518 18900 33570
rect 18508 33516 18900 33518
rect 18396 33358 18452 33516
rect 18844 33506 18900 33516
rect 20244 33460 20300 33966
rect 21252 34020 21308 34030
rect 21252 33926 21308 33964
rect 21980 34020 22036 34078
rect 21980 33954 22036 33964
rect 22316 34130 22372 34142
rect 22316 34078 22318 34130
rect 22370 34078 22372 34130
rect 22316 34020 22372 34078
rect 23324 34130 23380 34142
rect 23324 34078 23326 34130
rect 23378 34078 23380 34130
rect 22316 33954 22372 33964
rect 23044 34020 23100 34030
rect 23044 33926 23100 33964
rect 21644 33908 21700 33918
rect 20244 33394 20300 33404
rect 21532 33906 21700 33908
rect 21532 33854 21646 33906
rect 21698 33854 21700 33906
rect 21532 33852 21700 33854
rect 18172 33294 18174 33346
rect 18226 33294 18228 33346
rect 18172 33282 18228 33294
rect 18284 33346 18340 33358
rect 18284 33294 18286 33346
rect 18338 33294 18340 33346
rect 18060 31490 18116 31500
rect 17948 31164 18228 31220
rect 17948 30996 18004 31006
rect 17556 30882 17612 30894
rect 17556 30830 17558 30882
rect 17610 30830 17612 30882
rect 15596 30156 15764 30158
rect 15596 30146 15652 30156
rect 15484 29455 15596 29467
rect 15260 29428 15316 29438
rect 15260 29334 15316 29372
rect 15484 29403 15542 29455
rect 15594 29403 15596 29455
rect 15484 29372 15596 29403
rect 15316 26974 15372 26984
rect 15260 26964 15372 26974
rect 15316 26962 15372 26964
rect 15316 26910 15318 26962
rect 15370 26910 15372 26962
rect 15316 26908 15372 26910
rect 15260 26898 15372 26908
rect 15148 26290 15204 26302
rect 15148 26238 15150 26290
rect 15202 26238 15204 26290
rect 15148 25508 15204 26238
rect 15148 25442 15204 25452
rect 15036 24946 15148 24958
rect 15036 24894 15094 24946
rect 15146 24894 15148 24946
rect 15036 24882 15148 24894
rect 14252 24726 14254 24778
rect 14306 24726 14308 24778
rect 14588 24836 14644 24846
rect 14588 24778 14644 24780
rect 14252 24714 14308 24726
rect 14476 24750 14532 24762
rect 14476 24724 14478 24750
rect 14530 24724 14532 24750
rect 14588 24726 14590 24778
rect 14642 24726 14644 24778
rect 14588 24714 14644 24726
rect 14700 24724 14756 24734
rect 14476 24658 14532 24668
rect 14588 24612 14644 24622
rect 11900 24110 11902 24162
rect 11954 24110 11956 24162
rect 11900 24098 11956 24110
rect 13748 24498 13804 24510
rect 13748 24446 13750 24498
rect 13802 24446 13804 24498
rect 11564 23940 11620 23950
rect 10220 22530 10276 22540
rect 10668 23938 11620 23940
rect 10668 23886 11566 23938
rect 11618 23886 11620 23938
rect 10668 23884 11620 23886
rect 8764 22430 8766 22482
rect 8818 22430 8820 22482
rect 8764 22418 8820 22430
rect 10668 22484 10724 23884
rect 11564 23874 11620 23884
rect 13748 23940 13804 24446
rect 13748 23874 13804 23884
rect 13580 22596 13636 22606
rect 12012 22484 12068 22494
rect 10668 22482 10948 22484
rect 10668 22430 10670 22482
rect 10722 22430 10948 22482
rect 10668 22428 10948 22430
rect 10668 22418 10724 22428
rect 7980 22278 8036 22316
rect 10015 21812 10071 21822
rect 10015 21642 10071 21756
rect 10015 21590 10017 21642
rect 10069 21590 10071 21642
rect 10015 21578 10071 21590
rect 10892 21586 10948 22428
rect 11284 22372 11340 22382
rect 11284 22278 11340 22316
rect 12012 21642 12068 22428
rect 13580 22370 13636 22540
rect 13692 22538 13748 22550
rect 13692 22486 13694 22538
rect 13746 22486 13748 22538
rect 13692 22484 13748 22486
rect 13692 22418 13748 22428
rect 13580 22318 13582 22370
rect 13634 22318 13636 22370
rect 13580 22306 13636 22318
rect 13916 22370 13972 22382
rect 13916 22318 13918 22370
rect 13970 22318 13972 22370
rect 10892 21534 10894 21586
rect 10946 21534 10948 21586
rect 11900 21624 11956 21636
rect 11900 21588 11902 21624
rect 11954 21588 11956 21624
rect 12012 21590 12014 21642
rect 12066 21590 12068 21642
rect 13916 22036 13972 22318
rect 12012 21578 12068 21590
rect 12516 21588 12572 21598
rect 10892 21522 10948 21534
rect 11172 21530 11228 21542
rect 11172 21478 11174 21530
rect 11226 21478 11228 21530
rect 11900 21522 11956 21532
rect 12516 21494 12572 21532
rect 9772 21362 9828 21374
rect 9772 21310 9774 21362
rect 9826 21310 9828 21362
rect 9772 20804 9828 21310
rect 11172 20916 11228 21478
rect 9772 20738 9828 20748
rect 11116 20860 11228 20916
rect 11340 21474 11396 21486
rect 11340 21422 11342 21474
rect 11394 21422 11396 21474
rect 9772 20580 9828 20590
rect 9436 19236 9492 19246
rect 9436 19142 9492 19180
rect 9772 19207 9828 20524
rect 11004 20468 11060 20478
rect 11004 20130 11060 20412
rect 11004 20078 11006 20130
rect 11058 20078 11060 20130
rect 11004 20066 11060 20078
rect 11004 19460 11060 19470
rect 11116 19460 11172 20860
rect 11340 20580 11396 21422
rect 12012 20970 12068 20982
rect 12012 20918 12014 20970
rect 12066 20918 12068 20970
rect 11564 20804 11620 20814
rect 11564 20710 11620 20748
rect 11900 20802 11956 20814
rect 11900 20750 11902 20802
rect 11954 20750 11956 20802
rect 11340 20514 11396 20524
rect 11900 20468 11956 20750
rect 12012 20804 12068 20918
rect 13916 20914 13972 21980
rect 13916 20862 13918 20914
rect 13970 20862 13972 20914
rect 13916 20850 13972 20862
rect 12012 20738 12068 20748
rect 13468 20804 13524 20814
rect 13468 20710 13524 20748
rect 13748 20746 13804 20758
rect 13748 20694 13750 20746
rect 13802 20694 13804 20746
rect 13748 20692 13804 20694
rect 11900 20402 11956 20412
rect 13580 20636 13804 20692
rect 13580 20188 13636 20636
rect 12124 20132 12180 20142
rect 11247 20020 11303 20030
rect 11060 19404 11172 19460
rect 11228 20018 11303 20020
rect 11228 19966 11249 20018
rect 11301 19966 11303 20018
rect 11228 19954 11303 19966
rect 12124 20018 12180 20076
rect 12628 20132 12684 20142
rect 12628 20038 12684 20076
rect 13468 20132 13636 20188
rect 12124 19966 12126 20018
rect 12178 19966 12180 20018
rect 12124 19954 12180 19966
rect 11004 19366 11060 19404
rect 9772 19155 9774 19207
rect 9826 19155 9828 19207
rect 9772 19143 9828 19155
rect 10108 19234 10164 19246
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 9996 19066 10052 19078
rect 9996 19014 9998 19066
rect 10050 19014 10052 19066
rect 9996 18450 10052 19014
rect 10108 18564 10164 19182
rect 10668 19236 10724 19246
rect 11228 19236 11284 19954
rect 10668 19234 11284 19236
rect 10668 19182 10670 19234
rect 10722 19182 11284 19234
rect 10668 19180 11284 19182
rect 10108 18498 10164 18508
rect 10388 18564 10444 18574
rect 10388 18470 10444 18508
rect 9996 18398 9998 18450
rect 10050 18398 10052 18450
rect 9996 18386 10052 18398
rect 7644 18274 7700 18284
rect 9660 18228 9716 18238
rect 8764 18226 9716 18228
rect 8764 18174 9662 18226
rect 9714 18174 9716 18226
rect 8764 18172 9716 18174
rect 8764 17778 8820 18172
rect 9660 18162 9716 18172
rect 8764 17726 8766 17778
rect 8818 17726 8820 17778
rect 8764 17714 8820 17726
rect 10668 17778 10724 19180
rect 10668 17726 10670 17778
rect 10722 17726 10724 17778
rect 10668 17714 10724 17726
rect 7980 17666 8036 17678
rect 7980 17614 7982 17666
rect 8034 17614 8036 17666
rect 5068 15250 5124 15260
rect 5516 15316 5572 15326
rect 5292 15202 5348 15214
rect 5292 15150 5294 15202
rect 5346 15150 5348 15202
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5292 14644 5348 15150
rect 5292 14578 5348 14588
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4956 12740 5012 12750
rect 4956 12290 5012 12684
rect 4956 12238 4958 12290
rect 5010 12238 5012 12290
rect 4956 12226 5012 12238
rect 5516 12200 5572 15260
rect 7812 15316 7868 15326
rect 7980 15316 8036 17614
rect 11284 17444 11340 17454
rect 11004 17442 11340 17444
rect 11004 17390 11286 17442
rect 11338 17390 11340 17442
rect 11004 17388 11340 17390
rect 10332 15341 10388 15353
rect 7868 15260 8036 15316
rect 9436 15316 9492 15326
rect 7812 15222 7868 15260
rect 9436 15222 9492 15260
rect 10332 15289 10334 15341
rect 10386 15289 10388 15341
rect 7196 15202 7252 15214
rect 7196 15150 7198 15202
rect 7250 15150 7252 15202
rect 5852 14644 5908 14654
rect 5852 14550 5908 14588
rect 5964 14532 6020 14542
rect 5964 14463 5966 14476
rect 6018 14463 6020 14476
rect 6300 14532 6356 14542
rect 6748 14532 6804 14542
rect 6300 14530 6692 14532
rect 6300 14478 6302 14530
rect 6354 14478 6692 14530
rect 6300 14476 6692 14478
rect 6300 14466 6356 14476
rect 5964 14438 6020 14463
rect 2268 12180 2324 12190
rect 2268 9826 2324 12124
rect 5516 12180 5628 12200
rect 5572 12178 5628 12180
rect 5572 12126 5574 12178
rect 5626 12126 5628 12178
rect 5572 12124 5628 12126
rect 5516 12114 5628 12124
rect 3052 12066 3108 12078
rect 3052 12014 3054 12066
rect 3106 12014 3108 12066
rect 3052 11620 3108 12014
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 3052 11554 3108 11564
rect 3724 11620 3780 11630
rect 3724 11526 3780 11564
rect 4060 11396 4116 11406
rect 4060 11302 4116 11340
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4956 9940 5012 9950
rect 5516 9940 5572 12114
rect 6636 11396 6692 14476
rect 6748 14438 6804 14476
rect 6991 14474 7047 14486
rect 6991 14422 6993 14474
rect 7045 14422 7047 14474
rect 6991 13860 7047 14422
rect 7196 13970 7252 15150
rect 10332 15204 10388 15289
rect 10332 15138 10388 15148
rect 10444 15316 10500 15326
rect 7196 13918 7198 13970
rect 7250 13918 7252 13970
rect 7196 13906 7252 13918
rect 7868 14530 7924 14542
rect 7868 14478 7870 14530
rect 7922 14478 7924 14530
rect 7868 13970 7924 14478
rect 9940 14420 9996 14430
rect 10444 14420 10500 15260
rect 11004 15316 11060 17388
rect 11284 17378 11340 17388
rect 11004 15202 11060 15260
rect 11004 15150 11006 15202
rect 11058 15150 11060 15202
rect 11004 15138 11060 15150
rect 12964 15204 13020 15214
rect 12964 15110 13020 15148
rect 12460 14532 12516 14542
rect 9940 14418 10500 14420
rect 9940 14366 9942 14418
rect 9994 14366 10500 14418
rect 9940 14364 10500 14366
rect 9940 14354 9996 14364
rect 7868 13918 7870 13970
rect 7922 13918 7924 13970
rect 6972 13804 7047 13860
rect 6972 13188 7028 13804
rect 6972 13122 7028 13132
rect 7644 13188 7700 13198
rect 7420 12964 7476 12974
rect 7028 12906 7084 12918
rect 7028 12854 7030 12906
rect 7082 12854 7084 12906
rect 7420 12870 7476 12908
rect 7644 12934 7700 13132
rect 7644 12882 7646 12934
rect 7698 12882 7700 12934
rect 7868 12964 7924 13918
rect 10444 13746 10500 14364
rect 12124 14486 12180 14498
rect 12124 14434 12126 14486
rect 12178 14434 12180 14486
rect 12460 14438 12516 14476
rect 12908 14532 12964 14542
rect 12124 13972 12180 14434
rect 12124 13906 12180 13916
rect 12348 14362 12404 14374
rect 12348 14310 12350 14362
rect 12402 14310 12404 14362
rect 10444 13694 10446 13746
rect 10498 13694 10500 13746
rect 10444 13682 10500 13694
rect 11228 13634 11284 13646
rect 11228 13582 11230 13634
rect 11282 13582 11284 13634
rect 8652 13130 8708 13142
rect 8652 13078 8654 13130
rect 8706 13078 8708 13130
rect 8652 13076 8708 13078
rect 8652 13010 8708 13020
rect 9436 13074 9492 13086
rect 9436 13022 9438 13074
rect 9490 13022 9492 13074
rect 7868 12898 7924 12908
rect 8204 12962 8260 12974
rect 8204 12910 8206 12962
rect 8258 12910 8260 12962
rect 7028 12740 7084 12854
rect 7028 12674 7084 12684
rect 7196 12850 7252 12862
rect 7196 12798 7198 12850
rect 7250 12798 7252 12850
rect 6748 11396 6804 11406
rect 6636 11394 6804 11396
rect 6636 11342 6750 11394
rect 6802 11342 6804 11394
rect 6636 11340 6804 11342
rect 6748 10388 6804 11340
rect 6860 11396 6916 11406
rect 6860 11226 6916 11340
rect 7196 11355 7252 12798
rect 7644 12740 7700 12882
rect 8204 12852 8260 12910
rect 8540 12964 8596 12974
rect 8540 12870 8596 12908
rect 8988 12962 9044 12974
rect 8988 12910 8990 12962
rect 9042 12910 9044 12962
rect 8204 12786 8260 12796
rect 8988 12852 9044 12910
rect 9324 12964 9380 12974
rect 9324 12895 9326 12908
rect 9378 12895 9380 12908
rect 9324 12870 9380 12895
rect 8988 12786 9044 12796
rect 7644 12674 7700 12684
rect 9436 12180 9492 13022
rect 11228 13074 11284 13582
rect 11228 13022 11230 13074
rect 11282 13022 11284 13074
rect 11228 13010 11284 13022
rect 11340 13524 11396 13534
rect 11340 12947 11396 13468
rect 12236 13076 12292 13086
rect 11340 12895 11342 12947
rect 11394 12895 11396 12947
rect 11340 12883 11396 12895
rect 11564 12962 11620 12974
rect 11564 12910 11566 12962
rect 11618 12910 11620 12962
rect 11564 12740 11620 12910
rect 12236 12962 12292 13020
rect 12236 12910 12238 12962
rect 12290 12910 12292 12962
rect 12236 12898 12292 12910
rect 11564 12674 11620 12684
rect 12348 12740 12404 14310
rect 12572 13860 12628 13870
rect 12572 12935 12628 13804
rect 12572 12883 12574 12935
rect 12626 12883 12628 12935
rect 12572 12871 12628 12883
rect 12796 13412 12852 13422
rect 12348 12674 12404 12684
rect 12572 12794 12628 12806
rect 12572 12742 12574 12794
rect 12626 12742 12628 12794
rect 12572 12404 12628 12742
rect 9436 12114 9492 12124
rect 12460 12348 12628 12404
rect 12236 11508 12292 11518
rect 7196 11303 7198 11355
rect 7250 11303 7252 11355
rect 7196 11291 7252 11303
rect 7420 11394 7476 11406
rect 7420 11342 7422 11394
rect 7474 11342 7476 11394
rect 6860 11174 6862 11226
rect 6914 11174 6916 11226
rect 6860 11162 6916 11174
rect 5796 9940 5852 9950
rect 5516 9938 5908 9940
rect 5516 9886 5798 9938
rect 5850 9886 5908 9938
rect 5516 9884 5908 9886
rect 4956 9846 5012 9884
rect 5796 9874 5908 9884
rect 2268 9774 2270 9826
rect 2322 9774 2324 9826
rect 2268 9762 2324 9774
rect 3052 9826 3108 9838
rect 3052 9774 3054 9826
rect 3106 9774 3108 9826
rect 3052 9268 3108 9774
rect 3052 9202 3108 9212
rect 4172 9268 4228 9278
rect 4172 9174 4228 9212
rect 4508 9044 4564 9054
rect 4508 8950 4564 8988
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 5852 5124 5908 9874
rect 6748 9044 6804 10332
rect 7420 10052 7476 11342
rect 9996 10610 10052 10622
rect 9996 10558 9998 10610
rect 10050 10558 10052 10610
rect 9996 10500 10052 10558
rect 10388 10500 10444 10510
rect 9996 10498 10500 10500
rect 9996 10446 10390 10498
rect 10442 10446 10500 10498
rect 9996 10444 10500 10446
rect 10388 10434 10500 10444
rect 9660 10388 9716 10398
rect 9660 10294 9716 10332
rect 10444 10164 10500 10434
rect 7420 9986 7476 9996
rect 7980 10052 8036 10062
rect 7084 9940 7140 9950
rect 7868 9940 7924 9950
rect 7084 9826 7140 9884
rect 7644 9938 7924 9940
rect 7644 9886 7870 9938
rect 7922 9886 7924 9938
rect 7644 9884 7924 9886
rect 7084 9774 7086 9826
rect 7138 9774 7140 9826
rect 7084 9762 7140 9774
rect 7420 9828 7476 9838
rect 7420 9734 7476 9772
rect 7308 9210 7364 9222
rect 7308 9158 7310 9210
rect 7362 9158 7364 9210
rect 7196 9044 7252 9054
rect 6748 9042 7252 9044
rect 6748 8990 7198 9042
rect 7250 8990 7252 9042
rect 6748 8988 7252 8990
rect 7196 8484 7252 8988
rect 7308 9044 7364 9158
rect 7644 9098 7700 9884
rect 7868 9874 7924 9884
rect 7980 9811 8036 9996
rect 8988 10052 9044 10062
rect 7980 9759 7982 9811
rect 8034 9759 8036 9811
rect 7980 9747 8036 9759
rect 8204 9828 8260 9838
rect 8204 9734 8260 9772
rect 8988 9826 9044 9996
rect 8988 9774 8990 9826
rect 9042 9774 9044 9826
rect 7644 9046 7646 9098
rect 7698 9046 7700 9098
rect 7644 9034 7700 9046
rect 7868 9716 7924 9726
rect 7868 9042 7924 9660
rect 8708 9716 8764 9726
rect 8708 9622 8764 9660
rect 8988 9380 9044 9774
rect 9100 9828 9156 9838
rect 9100 9734 9156 9772
rect 8988 9314 9044 9324
rect 9772 9716 9828 9726
rect 7308 8978 7364 8988
rect 7868 8990 7870 9042
rect 7922 8990 7924 9042
rect 9772 9086 9828 9660
rect 9772 9034 9774 9086
rect 9826 9034 9828 9086
rect 9772 9022 9828 9034
rect 10108 9044 10164 9054
rect 7868 8978 7924 8990
rect 10108 8950 10164 8988
rect 10444 9042 10500 10108
rect 11508 10164 11564 10174
rect 11508 9938 11564 10108
rect 11508 9886 11510 9938
rect 11562 9886 11564 9938
rect 11508 9874 11564 9886
rect 10780 9828 10836 9838
rect 10780 9154 10836 9772
rect 10780 9102 10782 9154
rect 10834 9102 10836 9154
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 10444 8978 10500 8990
rect 10612 9044 10668 9054
rect 10612 8950 10668 8988
rect 10780 9044 10836 9102
rect 10780 8978 10836 8988
rect 10892 9380 10948 9390
rect 10892 9042 10948 9324
rect 10892 8990 10894 9042
rect 10946 8990 10948 9042
rect 10892 8978 10948 8990
rect 11788 9268 11844 9278
rect 11788 9042 11844 9212
rect 11788 8990 11790 9042
rect 11842 8990 11844 9042
rect 11788 8978 11844 8990
rect 12124 9044 12180 9054
rect 12124 8950 12180 8988
rect 9660 8930 9716 8942
rect 9660 8878 9662 8930
rect 9714 8878 9716 8930
rect 7532 8484 7588 8494
rect 7196 8482 7588 8484
rect 7196 8430 7534 8482
rect 7586 8430 7588 8482
rect 7196 8428 7588 8430
rect 7532 8418 7588 8428
rect 8204 8482 8260 8494
rect 8204 8430 8206 8482
rect 8258 8430 8260 8482
rect 7644 7588 7700 7598
rect 7644 6652 7700 7532
rect 8204 7252 8260 8430
rect 9660 8260 9716 8878
rect 11172 8818 11228 8830
rect 11172 8766 11174 8818
rect 11226 8766 11228 8818
rect 11172 8428 11228 8766
rect 12236 8428 12292 11452
rect 12460 10612 12516 12348
rect 12572 12178 12628 12190
rect 12572 12126 12574 12178
rect 12626 12126 12628 12178
rect 12572 11284 12628 12126
rect 12796 12066 12852 13356
rect 12908 12962 12964 14476
rect 13132 13748 13188 13758
rect 13132 13654 13188 13692
rect 13468 13412 13524 20132
rect 14588 18564 14644 24556
rect 14700 23266 14756 24668
rect 15036 24724 15092 24882
rect 15036 24658 15092 24668
rect 15260 24724 15316 26898
rect 15484 26628 15540 29372
rect 15708 29314 15764 30156
rect 16492 30154 16548 30166
rect 16492 30102 16494 30154
rect 16546 30102 16548 30154
rect 16492 29988 16548 30102
rect 16492 29922 16548 29932
rect 16716 30158 16718 30210
rect 16770 30158 16772 30210
rect 16716 29428 16772 30158
rect 16716 29362 16772 29372
rect 16828 30772 16884 30782
rect 15708 29262 15710 29314
rect 15762 29262 15764 29314
rect 15708 29250 15764 29262
rect 16212 29316 16268 29326
rect 16212 29222 16268 29260
rect 15372 26572 15540 26628
rect 16716 27748 16772 27758
rect 15372 26458 15428 26572
rect 15372 26406 15374 26458
rect 15426 26406 15428 26458
rect 15372 26394 15428 26406
rect 15260 24658 15316 24668
rect 16604 25172 16660 25182
rect 15092 24052 15148 24062
rect 15148 23996 15316 24052
rect 15092 23958 15148 23996
rect 14700 23214 14702 23266
rect 14754 23214 14756 23266
rect 14700 23202 14756 23214
rect 15260 23938 15316 23996
rect 15260 23886 15262 23938
rect 15314 23886 15316 23938
rect 15260 23604 15316 23886
rect 15036 23156 15092 23166
rect 14588 18498 14644 18508
rect 14812 23154 15092 23156
rect 14812 23102 15038 23154
rect 15090 23102 15092 23154
rect 14812 23100 15092 23102
rect 15260 23156 15316 23548
rect 15596 23716 15652 23726
rect 15484 23156 15540 23166
rect 15260 23154 15540 23156
rect 15260 23102 15486 23154
rect 15538 23102 15540 23154
rect 15260 23100 15540 23102
rect 14812 22260 14868 23100
rect 15036 23090 15092 23100
rect 15484 23090 15540 23100
rect 15316 22930 15372 22942
rect 15596 22932 15652 23660
rect 15876 23604 15932 23614
rect 15876 23378 15932 23548
rect 15876 23326 15878 23378
rect 15930 23326 15932 23378
rect 15876 23314 15932 23326
rect 16604 23378 16660 25116
rect 16604 23326 16606 23378
rect 16658 23326 16660 23378
rect 16604 23314 16660 23326
rect 15316 22878 15318 22930
rect 15370 22878 15372 22930
rect 15036 22484 15092 22494
rect 14924 22372 14980 22382
rect 14924 22278 14980 22316
rect 15036 22370 15092 22428
rect 15036 22318 15038 22370
rect 15090 22318 15092 22370
rect 15316 22372 15372 22878
rect 15036 22306 15092 22318
rect 15202 22314 15258 22326
rect 14700 18452 14756 18462
rect 14700 18358 14756 18396
rect 14812 18450 14868 22204
rect 15202 22262 15204 22314
rect 15256 22262 15258 22314
rect 15316 22306 15372 22316
rect 15484 22876 15652 22932
rect 16268 23154 16324 23166
rect 16268 23102 16270 23154
rect 16322 23102 16324 23154
rect 15202 22148 15258 22262
rect 15202 22082 15258 22092
rect 15484 21700 15540 22876
rect 15596 22484 15652 22494
rect 16268 22484 16324 23102
rect 15596 22482 16436 22484
rect 15596 22430 15598 22482
rect 15650 22430 16436 22482
rect 15596 22428 16436 22430
rect 15596 22418 15652 22428
rect 16380 22370 16436 22428
rect 16380 22318 16382 22370
rect 16434 22318 16436 22370
rect 16380 22306 16436 22318
rect 16604 22482 16660 22494
rect 16604 22430 16606 22482
rect 16658 22430 16660 22482
rect 16604 22370 16660 22430
rect 16604 22318 16606 22370
rect 16658 22318 16660 22370
rect 16604 22306 16660 22318
rect 16716 22484 16772 27692
rect 16100 22260 16156 22270
rect 16100 22166 16156 22204
rect 16604 22148 16660 22158
rect 15484 21634 15540 21644
rect 15932 21924 15988 21934
rect 15932 21586 15988 21868
rect 15932 21534 15934 21586
rect 15986 21534 15988 21586
rect 15932 21522 15988 21534
rect 16156 21700 16212 21710
rect 16156 21586 16212 21644
rect 16492 21588 16548 21598
rect 16156 21534 16158 21586
rect 16210 21534 16212 21586
rect 16156 21522 16212 21534
rect 16268 21586 16548 21588
rect 16268 21534 16494 21586
rect 16546 21534 16548 21586
rect 16268 21532 16548 21534
rect 15652 21364 15708 21374
rect 16268 21364 16324 21532
rect 16492 21522 16548 21532
rect 15596 21362 16324 21364
rect 15596 21310 15654 21362
rect 15706 21310 16324 21362
rect 16604 21418 16660 22092
rect 16716 21924 16772 22428
rect 16828 22484 16884 30716
rect 17556 30772 17612 30830
rect 17556 30706 17612 30716
rect 17108 30324 17164 30334
rect 17108 30266 17164 30268
rect 17108 30214 17110 30266
rect 17162 30214 17164 30266
rect 17108 30202 17164 30214
rect 16940 30100 16996 30110
rect 16940 30006 16996 30044
rect 17556 30100 17612 30110
rect 17556 30006 17612 30044
rect 17388 28532 17444 28542
rect 17388 27858 17444 28476
rect 17836 28084 17892 28094
rect 17500 28026 17556 28038
rect 17500 27974 17502 28026
rect 17554 27974 17556 28026
rect 17500 27972 17556 27974
rect 17500 27906 17556 27916
rect 17836 27914 17892 28028
rect 17388 27806 17390 27858
rect 17442 27806 17444 27858
rect 17836 27862 17838 27914
rect 17890 27862 17892 27914
rect 17836 27850 17892 27862
rect 17388 23716 17444 27806
rect 17388 23650 17444 23660
rect 17836 26292 17892 26302
rect 16996 22484 17052 22494
rect 16828 22482 17052 22484
rect 16828 22430 16830 22482
rect 16882 22430 16998 22482
rect 17050 22430 17052 22482
rect 16828 22428 17052 22430
rect 16828 22390 16884 22428
rect 16940 22418 17052 22428
rect 16716 21858 16772 21868
rect 16828 21588 16884 21598
rect 16828 21494 16884 21532
rect 16604 21366 16606 21418
rect 16658 21366 16660 21418
rect 16604 21354 16660 21366
rect 15596 21308 16324 21310
rect 15596 21298 15708 21308
rect 15596 18562 15652 21298
rect 15596 18510 15598 18562
rect 15650 18510 15652 18562
rect 14812 18398 14814 18450
rect 14866 18398 14868 18450
rect 14812 18386 14868 18398
rect 15204 18452 15260 18462
rect 15204 18358 15260 18396
rect 15484 18450 15540 18462
rect 15484 18398 15486 18450
rect 15538 18398 15540 18450
rect 14084 18340 14140 18350
rect 15036 18340 15092 18350
rect 14140 18284 14252 18340
rect 14084 18246 14140 18284
rect 14196 17778 14252 18284
rect 14420 18228 14476 18238
rect 14420 18226 14644 18228
rect 14420 18174 14422 18226
rect 14474 18174 14644 18226
rect 14420 18172 14644 18174
rect 14420 18162 14476 18172
rect 14196 17726 14198 17778
rect 14250 17726 14252 17778
rect 14196 17668 14252 17726
rect 14196 17602 14252 17612
rect 14476 17780 14532 17790
rect 14476 16882 14532 17724
rect 14476 16830 14478 16882
rect 14530 16830 14532 16882
rect 14028 15314 14084 15326
rect 14028 15262 14030 15314
rect 14082 15262 14084 15314
rect 13860 15204 13916 15214
rect 14028 15204 14084 15262
rect 13860 15202 14084 15204
rect 13860 15150 13862 15202
rect 13914 15150 14084 15202
rect 13860 15148 14084 15150
rect 13860 15138 13916 15148
rect 14028 14868 14084 15148
rect 14140 14868 14196 14878
rect 14028 14812 14140 14868
rect 13468 13346 13524 13356
rect 13580 14532 13636 14542
rect 13580 13746 13636 14476
rect 14140 14530 14196 14812
rect 14140 14478 14142 14530
rect 14194 14478 14196 14530
rect 14140 14466 14196 14478
rect 13580 13694 13582 13746
rect 13634 13694 13636 13746
rect 13580 13198 13636 13694
rect 13692 13860 13748 13870
rect 13692 13746 13748 13804
rect 14476 13860 14532 16830
rect 14588 16884 14644 18172
rect 14700 17668 14756 17678
rect 14700 17574 14756 17612
rect 15036 17666 15092 18284
rect 15484 18228 15540 18398
rect 15596 18452 15652 18510
rect 16324 19012 16380 19022
rect 15932 18450 15988 18462
rect 15596 18386 15652 18396
rect 15764 18394 15820 18406
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 15036 17602 15092 17614
rect 15260 18172 15540 18228
rect 15764 18342 15766 18394
rect 15818 18342 15820 18394
rect 15764 18340 15820 18342
rect 15260 17668 15316 18172
rect 15764 18116 15820 18284
rect 15484 18060 15820 18116
rect 15932 18398 15934 18450
rect 15986 18398 15988 18450
rect 15372 17780 15428 17818
rect 15372 17714 15428 17724
rect 15484 17622 15540 18060
rect 15260 17602 15316 17612
rect 15428 17610 15540 17622
rect 15428 17558 15430 17610
rect 15482 17558 15540 17610
rect 15428 17500 15540 17558
rect 15708 17668 15764 17678
rect 15932 17668 15988 18398
rect 16324 18450 16380 18956
rect 16324 18398 16326 18450
rect 16378 18398 16380 18450
rect 16324 18386 16380 18398
rect 16604 18452 16660 18462
rect 16604 18358 16660 18396
rect 16716 18450 16772 18462
rect 16716 18398 16718 18450
rect 16770 18398 16772 18450
rect 16716 18340 16772 18398
rect 16716 18274 16772 18284
rect 15708 17666 15988 17668
rect 15708 17614 15710 17666
rect 15762 17614 15988 17666
rect 15708 17612 15988 17614
rect 14700 16884 14756 16894
rect 14588 16882 14756 16884
rect 14588 16830 14702 16882
rect 14754 16830 14756 16882
rect 14588 16828 14756 16830
rect 14700 16818 14756 16828
rect 14980 16660 15036 16670
rect 14924 16658 15036 16660
rect 14924 16606 14982 16658
rect 15034 16606 15036 16658
rect 14924 16594 15036 16606
rect 14924 16098 14980 16594
rect 14924 16046 14926 16098
rect 14978 16046 14980 16098
rect 14924 16034 14980 16046
rect 15260 15876 15316 15886
rect 14812 15874 15316 15876
rect 14812 15822 15262 15874
rect 15314 15822 15316 15874
rect 14812 15820 15316 15822
rect 14812 15314 14868 15820
rect 15260 15810 15316 15820
rect 15708 15540 15764 17612
rect 16940 16100 16996 22418
rect 17724 22372 17780 22382
rect 17724 22278 17780 22316
rect 17556 22260 17612 22270
rect 17556 22166 17612 22204
rect 17836 20188 17892 26236
rect 17948 25172 18004 30940
rect 18060 27860 18116 27870
rect 18060 27766 18116 27804
rect 18172 26414 18228 31164
rect 18284 30996 18340 33294
rect 18396 33348 18506 33358
rect 18396 33292 18450 33348
rect 18450 33254 18506 33292
rect 19292 33348 19348 33358
rect 18284 30930 18340 30940
rect 18396 33124 18452 33134
rect 18284 30772 18340 30782
rect 18396 30772 18452 33068
rect 18844 31556 18900 31566
rect 18844 31038 18900 31500
rect 18844 30986 18846 31038
rect 18898 30986 18900 31038
rect 18844 30974 18900 30986
rect 19180 30996 19236 31006
rect 19180 30902 19236 30940
rect 18284 30770 18452 30772
rect 18284 30718 18286 30770
rect 18338 30718 18452 30770
rect 18284 30716 18452 30718
rect 18732 30882 18788 30894
rect 18732 30830 18734 30882
rect 18786 30830 18788 30882
rect 18284 30100 18340 30716
rect 18732 30324 18788 30830
rect 18732 30258 18788 30268
rect 18284 28756 18340 30044
rect 18284 28690 18340 28700
rect 19068 28642 19124 28654
rect 19068 28590 19070 28642
rect 19122 28590 19124 28642
rect 19068 28532 19124 28590
rect 19068 28466 19124 28476
rect 18788 28084 18844 28094
rect 18788 27990 18844 28028
rect 19292 28084 19348 33292
rect 19460 33348 19516 33358
rect 19460 33254 19516 33292
rect 21532 33124 21588 33852
rect 21644 33842 21700 33852
rect 22484 33908 22540 33918
rect 22484 33814 22540 33852
rect 23324 33908 23380 34078
rect 23324 33842 23380 33852
rect 21644 33572 21700 33582
rect 21644 33346 21700 33516
rect 22596 33572 22652 33582
rect 22596 33460 22652 33516
rect 23660 33572 23716 34302
rect 23660 33506 23716 33516
rect 24556 33570 24612 37996
rect 25004 37828 25060 37838
rect 25004 36594 25060 37772
rect 26348 37380 26404 37390
rect 26348 37322 26404 37324
rect 25452 37299 25508 37311
rect 25452 37247 25454 37299
rect 25506 37247 25508 37299
rect 25452 36708 25508 37247
rect 25900 37302 25956 37314
rect 25900 37268 25902 37302
rect 25954 37268 25956 37302
rect 26348 37270 26350 37322
rect 26402 37270 26404 37322
rect 26684 37378 26740 40236
rect 26796 40226 26852 40236
rect 28364 38834 28420 38846
rect 28364 38782 28366 38834
rect 28418 38782 28420 38834
rect 28028 38052 28084 38062
rect 26684 37326 26686 37378
rect 26738 37326 26740 37378
rect 26684 37314 26740 37326
rect 27804 37380 27860 37390
rect 26348 37258 26404 37270
rect 26504 37299 26560 37311
rect 25004 36542 25006 36594
rect 25058 36542 25060 36594
rect 25004 36530 25060 36542
rect 25116 36652 25508 36708
rect 25564 37156 25620 37166
rect 24836 36426 24892 36438
rect 24836 36374 24838 36426
rect 24890 36374 24892 36426
rect 24836 36372 24892 36374
rect 25116 36372 25172 36652
rect 24836 36316 25172 36372
rect 25228 36482 25284 36494
rect 25228 36430 25230 36482
rect 25282 36430 25284 36482
rect 24836 35812 24892 36316
rect 24556 33518 24558 33570
rect 24610 33518 24612 33570
rect 21644 33294 21646 33346
rect 21698 33294 21700 33346
rect 21644 33282 21700 33294
rect 22428 33458 22652 33460
rect 22428 33406 22598 33458
rect 22650 33406 22652 33458
rect 22428 33404 22652 33406
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 21196 32116 21252 32126
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20076 30996 20132 31006
rect 19964 30322 20020 30334
rect 19964 30270 19966 30322
rect 20018 30270 20020 30322
rect 19964 30100 20020 30270
rect 19964 30034 20020 30044
rect 20076 30166 20132 30940
rect 20076 30114 20078 30166
rect 20130 30114 20132 30166
rect 20076 29988 20132 30114
rect 20412 30210 20468 30222
rect 20412 30158 20414 30210
rect 20466 30158 20468 30210
rect 20412 30100 20468 30158
rect 20412 30034 20468 30044
rect 21084 30100 21140 30110
rect 20188 29988 20244 29998
rect 21084 29988 21140 30044
rect 20076 29932 20188 29988
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 29428 19572 29438
rect 19516 28754 19572 29372
rect 20188 28868 20244 29932
rect 21046 29932 21140 29988
rect 21046 29464 21102 29932
rect 20748 29426 20804 29438
rect 20748 29374 20750 29426
rect 20802 29374 20804 29426
rect 20468 29316 20524 29326
rect 20748 29316 20804 29374
rect 20860 29428 20916 29438
rect 21046 29412 21048 29464
rect 21100 29412 21102 29464
rect 21046 29400 21102 29412
rect 20860 29334 20916 29372
rect 20468 29314 20804 29316
rect 20468 29262 20470 29314
rect 20522 29262 20804 29314
rect 20468 29260 20804 29262
rect 20468 29250 20524 29260
rect 20188 28802 20244 28812
rect 20636 28868 20692 28878
rect 20636 28774 20692 28812
rect 19516 28702 19518 28754
rect 19570 28702 19572 28754
rect 19516 28690 19572 28702
rect 20300 28644 20356 28654
rect 20412 28644 20468 28654
rect 20300 28642 20412 28644
rect 19292 28018 19348 28028
rect 19404 28598 19460 28610
rect 19404 28546 19406 28598
rect 19458 28546 19460 28598
rect 20300 28590 20302 28642
rect 20354 28590 20412 28642
rect 20300 28588 20412 28590
rect 20300 28578 20356 28588
rect 18620 27860 18676 27870
rect 18508 26964 18564 26974
rect 18172 26404 18284 26414
rect 18172 26348 18228 26404
rect 18228 26310 18284 26348
rect 18508 26292 18564 26908
rect 18508 26198 18564 26236
rect 18620 26290 18676 27804
rect 19404 27748 19460 28546
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19404 27682 19460 27692
rect 18900 27636 18956 27646
rect 18900 26964 18956 27580
rect 18900 26870 18956 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19124 26404 19180 26414
rect 19124 26346 19180 26348
rect 18956 26292 19012 26302
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 18620 26068 18676 26238
rect 18508 26012 18676 26068
rect 18732 26290 19012 26292
rect 18732 26238 18958 26290
rect 19010 26238 19012 26290
rect 19124 26294 19126 26346
rect 19178 26294 19180 26346
rect 19124 26282 19180 26294
rect 19292 26290 19348 26302
rect 18732 26236 19012 26238
rect 18172 25732 18228 25742
rect 18172 25506 18228 25676
rect 18172 25454 18174 25506
rect 18226 25454 18228 25506
rect 18172 25442 18228 25454
rect 18396 25506 18452 25518
rect 18396 25454 18398 25506
rect 18450 25454 18452 25506
rect 17948 25106 18004 25116
rect 18396 25172 18452 25454
rect 18396 25106 18452 25116
rect 18508 23278 18564 26012
rect 18732 25742 18788 26236
rect 18956 26226 19012 26236
rect 19292 26238 19294 26290
rect 19346 26238 19348 26290
rect 19068 26180 19124 26190
rect 18676 25730 18788 25742
rect 18676 25678 18678 25730
rect 18730 25678 18788 25730
rect 18676 25676 18788 25678
rect 18844 26068 18900 26078
rect 18676 25666 18732 25676
rect 18508 23266 18620 23278
rect 18508 23214 18566 23266
rect 18618 23214 18620 23266
rect 18508 23212 18620 23214
rect 18564 23202 18620 23212
rect 18060 23154 18116 23166
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 18060 22596 18116 23102
rect 18284 23156 18340 23166
rect 18284 23154 18452 23156
rect 18284 23102 18286 23154
rect 18338 23102 18452 23154
rect 18284 23100 18452 23102
rect 18284 23090 18340 23100
rect 18060 22530 18116 22540
rect 17948 22484 18004 22494
rect 17948 22370 18004 22428
rect 17948 22318 17950 22370
rect 18002 22318 18004 22370
rect 17948 22306 18004 22318
rect 18228 22260 18284 22270
rect 18228 22166 18284 22204
rect 18396 22036 18452 23100
rect 18620 22596 18676 22606
rect 18620 22370 18676 22540
rect 18620 22318 18622 22370
rect 18674 22318 18676 22370
rect 18620 22306 18676 22318
rect 18396 21970 18452 21980
rect 17836 20132 18228 20188
rect 18172 19346 18228 20132
rect 18172 19294 18174 19346
rect 18226 19294 18228 19346
rect 18172 19282 18228 19294
rect 17780 19236 17836 19246
rect 17612 19180 17780 19236
rect 17388 18340 17444 18350
rect 17388 18228 17444 18284
rect 17500 18228 17556 18238
rect 17388 18226 17556 18228
rect 17388 18174 17502 18226
rect 17554 18174 17556 18226
rect 17388 18172 17556 18174
rect 17388 17666 17444 18172
rect 17500 18162 17556 18172
rect 17388 17614 17390 17666
rect 17442 17614 17444 17666
rect 17388 17602 17444 17614
rect 16940 16034 16996 16044
rect 17612 15550 17668 19180
rect 17780 19142 17836 19180
rect 18844 18676 18900 26012
rect 18956 22484 19012 22522
rect 18956 22418 19012 22428
rect 18956 22314 19012 22326
rect 18956 22262 18958 22314
rect 19010 22262 19012 22314
rect 18956 22036 19012 22262
rect 18956 21970 19012 21980
rect 19068 21476 19124 26124
rect 19180 25732 19236 25742
rect 19180 25506 19236 25676
rect 19180 25454 19182 25506
rect 19234 25454 19236 25506
rect 19180 25284 19236 25454
rect 19292 25618 19348 26238
rect 19404 26292 19460 26302
rect 19404 26290 19572 26292
rect 19404 26238 19406 26290
rect 19458 26238 19572 26290
rect 19404 26236 19572 26238
rect 19404 26226 19460 26236
rect 19292 25566 19294 25618
rect 19346 25566 19348 25618
rect 19292 25508 19348 25566
rect 19292 25442 19348 25452
rect 19180 25218 19236 25228
rect 19516 24610 19572 26236
rect 19684 26068 19740 26078
rect 19684 25974 19740 26012
rect 19852 25506 19908 25518
rect 19628 25450 19684 25462
rect 19628 25398 19630 25450
rect 19682 25398 19684 25450
rect 19628 25396 19684 25398
rect 19628 25330 19684 25340
rect 19852 25454 19854 25506
rect 19906 25454 19908 25506
rect 19852 25284 19908 25454
rect 20300 25396 20356 25406
rect 19852 25228 20244 25284
rect 19628 25172 19684 25182
rect 19628 24948 19684 25116
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 25228
rect 19628 24892 19946 24948
rect 19890 24760 19946 24892
rect 19890 24708 19892 24760
rect 19944 24708 19946 24760
rect 19890 24696 19946 24708
rect 20076 24892 20188 24948
rect 20076 24722 20132 24892
rect 20188 24882 20244 24892
rect 20076 24670 20078 24722
rect 20130 24670 20132 24722
rect 20076 24658 20132 24670
rect 20188 24724 20244 24734
rect 20300 24724 20356 25340
rect 20188 24722 20356 24724
rect 20188 24670 20190 24722
rect 20242 24670 20356 24722
rect 20188 24668 20356 24670
rect 20188 24658 20244 24668
rect 19516 24558 19518 24610
rect 19570 24558 19572 24610
rect 19516 24546 19572 24558
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20076 22596 20132 22606
rect 19292 22370 19348 22382
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 19292 21588 19348 22318
rect 19628 22370 19684 22382
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19460 22260 19516 22270
rect 19460 21810 19516 22204
rect 19628 22260 19684 22318
rect 19628 22194 19684 22204
rect 20076 22260 20132 22540
rect 20412 22484 20468 28588
rect 20748 26292 20804 29260
rect 20748 26236 21140 26292
rect 20412 22418 20468 22428
rect 20076 22148 20132 22204
rect 20076 22092 20244 22148
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22092
rect 19460 21758 19462 21810
rect 19514 21758 19516 21810
rect 19460 21746 19516 21758
rect 20076 21756 20244 21812
rect 19292 21522 19348 21532
rect 20076 21586 20132 21756
rect 20972 21700 21028 21710
rect 20076 21534 20078 21586
rect 20130 21534 20132 21586
rect 20076 21522 20132 21534
rect 20300 21588 20356 21598
rect 19068 21410 19124 21420
rect 19796 21476 19852 21486
rect 19796 21382 19852 21420
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20300 20188 20356 21532
rect 20300 20132 20804 20188
rect 20076 19234 20132 19246
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19012 20132 19182
rect 20076 18956 20244 19012
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18844 18620 20132 18676
rect 17836 18450 17892 18462
rect 17836 18398 17838 18450
rect 17890 18398 17892 18450
rect 17836 17892 17892 18398
rect 19964 18450 20020 18462
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19964 18340 20020 18398
rect 20076 18450 20132 18620
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 20076 18386 20132 18398
rect 19964 18274 20020 18284
rect 20188 18228 20244 18956
rect 20356 18452 20412 18462
rect 20636 18452 20692 18462
rect 20356 18450 20692 18452
rect 20356 18398 20358 18450
rect 20410 18398 20638 18450
rect 20690 18398 20692 18450
rect 20356 18396 20692 18398
rect 20356 18386 20412 18396
rect 20636 18386 20692 18396
rect 20188 18162 20244 18172
rect 17836 17826 17892 17836
rect 20748 17892 20804 20132
rect 20860 19236 20916 19246
rect 20860 19142 20916 19180
rect 20748 17826 20804 17836
rect 20860 18788 20916 18798
rect 20748 17668 20804 17678
rect 17724 17444 17780 17454
rect 17724 17350 17780 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20748 17108 20804 17612
rect 20860 17444 20916 18732
rect 20972 18564 21028 21644
rect 21084 18788 21140 26236
rect 21084 18722 21140 18732
rect 20972 18508 21140 18564
rect 20972 18228 21028 18238
rect 20972 18134 21028 18172
rect 21084 17556 21140 18508
rect 20860 17378 20916 17388
rect 21028 17500 21140 17556
rect 20748 17052 20916 17108
rect 20748 16884 20804 16894
rect 20748 16790 20804 16828
rect 20860 16882 20916 17052
rect 20860 16830 20862 16882
rect 20914 16830 20916 16882
rect 21028 16938 21084 17500
rect 21028 16886 21030 16938
rect 21082 16886 21084 16938
rect 21028 16874 21084 16886
rect 21196 17108 21252 32060
rect 21532 30772 21588 33068
rect 21980 33122 22036 33134
rect 21980 33070 21982 33122
rect 22034 33070 22036 33122
rect 21868 32562 21924 32574
rect 21868 32510 21870 32562
rect 21922 32510 21924 32562
rect 21868 31892 21924 32510
rect 21868 31826 21924 31836
rect 21980 32004 22036 33070
rect 21532 30706 21588 30716
rect 21476 30100 21532 30110
rect 21476 30006 21532 30044
rect 21980 30100 22036 31948
rect 22428 32116 22484 33404
rect 22596 33394 22652 33404
rect 23436 33348 23492 33358
rect 23268 33346 23492 33348
rect 23268 33294 23438 33346
rect 23490 33294 23492 33346
rect 23268 33292 23492 33294
rect 23268 33124 23324 33292
rect 23436 33282 23492 33292
rect 23660 33348 23716 33358
rect 23660 33254 23716 33292
rect 23940 33348 23996 33358
rect 24220 33348 24276 33358
rect 23940 33346 24276 33348
rect 23940 33294 23942 33346
rect 23994 33294 24222 33346
rect 24274 33294 24276 33346
rect 23940 33292 24276 33294
rect 23940 33282 23996 33292
rect 24220 33282 24276 33292
rect 23268 33030 23324 33068
rect 22652 32676 22708 32686
rect 22652 32562 22708 32620
rect 24556 32676 24612 33518
rect 24668 35756 24892 35812
rect 24668 33348 24724 35756
rect 25228 35140 25284 36430
rect 25564 36444 25620 37100
rect 25564 36392 25566 36444
rect 25618 36392 25620 36444
rect 25564 36380 25620 36392
rect 25340 35474 25396 35486
rect 25340 35422 25342 35474
rect 25394 35422 25396 35474
rect 25340 35140 25396 35422
rect 25228 35138 25396 35140
rect 25228 35086 25230 35138
rect 25282 35086 25396 35138
rect 25228 35084 25396 35086
rect 25228 35074 25284 35084
rect 24836 34916 24892 34926
rect 24836 34822 24892 34860
rect 25620 34916 25676 34926
rect 25620 34822 25676 34860
rect 25788 34914 25844 34926
rect 25788 34862 25790 34914
rect 25842 34862 25844 34914
rect 25788 34692 25844 34862
rect 25788 34626 25844 34636
rect 25900 34916 25956 37212
rect 26504 37247 26506 37299
rect 26558 37247 26560 37299
rect 26504 37156 26560 37247
rect 27580 37268 27636 37278
rect 27580 37174 27636 37212
rect 27804 37268 27860 37324
rect 27916 37268 27972 37278
rect 27804 37266 27972 37268
rect 27804 37214 27918 37266
rect 27970 37214 27972 37266
rect 27804 37212 27972 37214
rect 26504 37090 26560 37100
rect 26572 35476 26628 35486
rect 26572 35474 26740 35476
rect 26572 35422 26574 35474
rect 26626 35422 26740 35474
rect 26572 35420 26740 35422
rect 26572 35410 26628 35420
rect 24668 33282 24724 33292
rect 24556 32610 24612 32620
rect 22652 32510 22654 32562
rect 22706 32510 22708 32562
rect 22652 32498 22708 32510
rect 24556 32450 24612 32462
rect 24556 32398 24558 32450
rect 24610 32398 24612 32450
rect 22428 31778 22484 32060
rect 23324 32116 23380 32126
rect 23324 31948 23380 32060
rect 23324 31892 23436 31948
rect 23380 31890 23436 31892
rect 23380 31838 23382 31890
rect 23434 31838 23436 31890
rect 23380 31826 23436 31838
rect 22428 31726 22430 31778
rect 22482 31726 22484 31778
rect 22428 31714 22484 31726
rect 24556 31780 24612 32398
rect 25396 32450 25452 32462
rect 25396 32398 25398 32450
rect 25450 32398 25452 32450
rect 25396 31948 25452 32398
rect 25900 31948 25956 34860
rect 26684 34914 26740 35420
rect 26852 35252 26908 35262
rect 26852 35138 26908 35196
rect 26852 35086 26854 35138
rect 26906 35086 26908 35138
rect 26852 35074 26908 35086
rect 26684 34862 26686 34914
rect 26738 34862 26740 34914
rect 26684 34850 26740 34862
rect 27356 34916 27412 34926
rect 27356 34822 27412 34860
rect 27804 34914 27860 37212
rect 27916 37202 27972 37212
rect 28028 37098 28084 37996
rect 28364 38052 28420 38782
rect 28364 37986 28420 37996
rect 28028 37046 28030 37098
rect 28082 37046 28084 37098
rect 28028 37034 28084 37046
rect 28364 35364 28420 35374
rect 27804 34862 27806 34914
rect 27858 34862 27860 34914
rect 27804 34692 27860 34862
rect 28028 34916 28084 34926
rect 27804 34626 27860 34636
rect 27916 34802 27972 34814
rect 27916 34750 27918 34802
rect 27970 34750 27972 34802
rect 27804 34132 27860 34142
rect 27916 34132 27972 34750
rect 27804 34130 27972 34132
rect 27804 34078 27806 34130
rect 27858 34078 27972 34130
rect 27804 34076 27972 34078
rect 28028 34169 28084 34860
rect 28252 34914 28308 34926
rect 28252 34862 28254 34914
rect 28306 34862 28308 34914
rect 28252 34356 28308 34862
rect 28252 34290 28308 34300
rect 28364 34298 28420 35308
rect 28476 34914 28532 34926
rect 28476 34862 28478 34914
rect 28530 34862 28532 34914
rect 28476 34804 28532 34862
rect 28476 34738 28532 34748
rect 28364 34246 28366 34298
rect 28418 34246 28420 34298
rect 28364 34234 28420 34246
rect 28028 34117 28030 34169
rect 28082 34117 28084 34169
rect 27804 34066 27860 34076
rect 27300 34018 27356 34030
rect 27300 33966 27302 34018
rect 27354 33966 27356 34018
rect 27300 33572 27356 33966
rect 27300 33506 27356 33516
rect 24556 31714 24612 31724
rect 24668 31892 24724 31902
rect 22764 31556 22820 31566
rect 22652 31554 22820 31556
rect 22652 31502 22766 31554
rect 22818 31502 22820 31554
rect 22652 31500 22820 31502
rect 21980 29662 22036 30044
rect 22428 30212 22484 30222
rect 21980 29650 22092 29662
rect 21980 29598 22038 29650
rect 22090 29598 22092 29650
rect 21980 29596 22092 29598
rect 22036 29586 22092 29596
rect 21420 29204 21476 29214
rect 21420 29110 21476 29148
rect 21980 28642 22036 28654
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21756 27076 21812 27086
rect 21980 27076 22036 28590
rect 21812 27020 22036 27076
rect 21756 26982 21812 27020
rect 21420 26962 21476 26974
rect 21420 26910 21422 26962
rect 21474 26910 21476 26962
rect 21420 26292 21476 26910
rect 21420 25396 21476 26236
rect 21420 25330 21476 25340
rect 21868 24724 21924 24734
rect 21364 23268 21420 23278
rect 21364 23174 21420 23212
rect 21644 23268 21700 23278
rect 21644 23181 21700 23212
rect 21644 23129 21646 23181
rect 21698 23129 21700 23181
rect 21644 23117 21700 23129
rect 21868 20914 21924 24668
rect 22428 22932 22484 30156
rect 22652 27972 22708 31500
rect 22764 31490 22820 31500
rect 24108 29988 24164 29998
rect 22652 27906 22708 27916
rect 22764 28756 22820 28766
rect 22764 27300 22820 28700
rect 23884 28644 23940 28654
rect 23660 28642 23940 28644
rect 23660 28590 23886 28642
rect 23938 28590 23940 28642
rect 23660 28588 23940 28590
rect 23660 27748 23716 28588
rect 23884 28578 23940 28588
rect 23548 27692 23716 27748
rect 22596 27244 23044 27300
rect 22596 27186 22652 27244
rect 22596 27134 22598 27186
rect 22650 27134 22652 27186
rect 22596 27122 22652 27134
rect 22988 27036 23044 27244
rect 23548 27186 23604 27692
rect 23548 27134 23550 27186
rect 23602 27134 23604 27186
rect 23548 27122 23604 27134
rect 22876 27018 22932 27030
rect 22876 26966 22878 27018
rect 22930 26966 22932 27018
rect 22876 26628 22932 26966
rect 22708 26572 22932 26628
rect 22988 26984 22990 27036
rect 23042 26984 23044 27036
rect 22708 26514 22764 26572
rect 22708 26462 22710 26514
rect 22762 26462 22764 26514
rect 22708 26450 22764 26462
rect 22540 26292 22596 26302
rect 22540 25508 22596 26236
rect 22988 25844 23044 26984
rect 23716 27018 23772 27030
rect 23716 26966 23718 27018
rect 23770 26966 23772 27018
rect 23716 26404 23772 26966
rect 23716 26348 24052 26404
rect 22540 25442 22596 25452
rect 22764 25788 23044 25844
rect 22764 24500 22820 25788
rect 22988 25508 23044 25518
rect 22988 25414 23044 25452
rect 23864 25450 23920 25462
rect 23864 25398 23866 25450
rect 23918 25398 23920 25450
rect 23864 25060 23920 25398
rect 23996 25396 24052 26348
rect 24108 25844 24164 29932
rect 24668 28756 24724 31836
rect 25340 31892 25452 31948
rect 25676 31892 25956 31948
rect 27132 33348 27188 33358
rect 25340 31826 25396 31836
rect 25060 28756 25116 28766
rect 24668 28754 25116 28756
rect 24668 28702 25062 28754
rect 25114 28702 25116 28754
rect 24668 28700 25116 28702
rect 24668 28642 24724 28700
rect 25060 28690 25116 28700
rect 24668 28590 24670 28642
rect 24722 28590 24724 28642
rect 24668 28578 24724 28590
rect 25228 27860 25284 27870
rect 24724 27748 24780 27758
rect 24724 27654 24780 27692
rect 25004 27748 25060 27758
rect 24276 26180 24332 26190
rect 25004 26180 25060 27692
rect 25228 26180 25284 27804
rect 25564 27860 25620 27870
rect 25564 27766 25620 27804
rect 25676 27746 25732 31892
rect 25788 31780 25844 31790
rect 25788 31686 25844 31724
rect 25956 31556 26012 31566
rect 25956 31554 26516 31556
rect 25956 31502 25958 31554
rect 26010 31502 26516 31554
rect 25956 31500 26516 31502
rect 25956 31490 26012 31500
rect 26460 31050 26516 31500
rect 26460 30998 26462 31050
rect 26514 30998 26516 31050
rect 27132 31106 27188 33292
rect 27748 31892 27804 31902
rect 27748 31798 27804 31836
rect 28028 31220 28084 34117
rect 28476 34130 28532 34142
rect 28476 34078 28478 34130
rect 28530 34078 28532 34130
rect 28476 33572 28532 34078
rect 28476 32004 28532 33516
rect 28476 31938 28532 31948
rect 28588 32562 28644 40348
rect 29316 40404 29372 40414
rect 29316 40310 29372 40348
rect 29708 40404 29764 40414
rect 29708 40310 29764 40348
rect 32788 40404 32844 40910
rect 35980 40514 36036 41132
rect 36372 40962 36428 40974
rect 36372 40910 36374 40962
rect 36426 40910 36428 40962
rect 35980 40462 35982 40514
rect 36034 40462 36036 40514
rect 35980 40450 36036 40462
rect 36092 40516 36148 40526
rect 32788 40338 32844 40348
rect 33292 40404 33348 40414
rect 33292 40310 33348 40348
rect 30492 40292 30548 40302
rect 30268 40290 30548 40292
rect 30268 40238 30494 40290
rect 30546 40238 30548 40290
rect 30268 40236 30548 40238
rect 30268 39842 30324 40236
rect 30492 40226 30548 40236
rect 34076 40290 34132 40302
rect 34076 40238 34078 40290
rect 34130 40238 34132 40290
rect 30268 39790 30270 39842
rect 30322 39790 30324 39842
rect 30268 39778 30324 39790
rect 32844 39844 32900 39854
rect 32844 39750 32900 39788
rect 34076 39844 34132 40238
rect 36092 40180 36148 40460
rect 36372 40404 36428 40910
rect 39676 40628 39732 40638
rect 39676 40534 39732 40572
rect 40124 40628 40180 41945
rect 41132 41860 41188 41870
rect 41132 41766 41188 41804
rect 43708 41186 43764 45200
rect 40124 40562 40180 40572
rect 41804 41158 41860 41170
rect 41804 41106 41806 41158
rect 41858 41106 41860 41158
rect 43708 41134 43710 41186
rect 43762 41134 43764 41186
rect 43708 41122 43764 41134
rect 39004 40516 39060 40526
rect 39004 40422 39060 40460
rect 39340 40516 39396 40526
rect 36372 40292 36428 40348
rect 39340 40402 39396 40460
rect 40404 40404 40460 40414
rect 40796 40404 40852 40414
rect 39340 40350 39342 40402
rect 39394 40350 39396 40402
rect 39340 40338 39396 40350
rect 40348 40402 40852 40404
rect 40348 40350 40406 40402
rect 40458 40350 40798 40402
rect 40850 40350 40852 40402
rect 40348 40348 40852 40350
rect 40348 40338 40460 40348
rect 40796 40338 40852 40348
rect 36372 40236 36596 40292
rect 35980 40124 36148 40180
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34076 39778 34132 39788
rect 29036 39620 29092 39630
rect 28812 39618 29092 39620
rect 28812 39566 29038 39618
rect 29090 39566 29092 39618
rect 28812 39564 29092 39566
rect 28700 38849 28756 38861
rect 28700 38797 28702 38849
rect 28754 38797 28756 38849
rect 28700 37828 28756 38797
rect 28812 38722 28868 39564
rect 29036 39554 29092 39564
rect 29260 39618 29316 39630
rect 29260 39566 29262 39618
rect 29314 39566 29316 39618
rect 29148 39508 29204 39518
rect 28812 38670 28814 38722
rect 28866 38670 28868 38722
rect 28812 38658 28868 38670
rect 28924 38836 28980 38846
rect 28700 37156 28756 37772
rect 28700 37090 28756 37100
rect 28924 36260 28980 38780
rect 29036 38052 29092 38062
rect 29036 37958 29092 37996
rect 29148 37380 29204 39452
rect 29260 38836 29316 39566
rect 29540 39620 29596 39630
rect 29932 39620 29988 39630
rect 29540 39618 29988 39620
rect 29540 39566 29542 39618
rect 29594 39566 29934 39618
rect 29986 39566 29988 39618
rect 29540 39564 29988 39566
rect 29540 39554 29596 39564
rect 29932 39554 29988 39564
rect 32508 39618 32564 39630
rect 32508 39566 32510 39618
rect 32562 39566 32564 39618
rect 29260 38770 29316 38780
rect 29260 38108 29764 38164
rect 29260 38050 29316 38108
rect 29260 37998 29262 38050
rect 29314 37998 29316 38050
rect 29260 37986 29316 37998
rect 29708 38052 29764 38108
rect 29820 38052 29876 38062
rect 29708 38050 29988 38052
rect 29708 37998 29822 38050
rect 29874 37998 29988 38050
rect 29708 37996 29988 37998
rect 29820 37986 29876 37996
rect 29540 37940 29596 37950
rect 29540 37846 29596 37884
rect 29372 37380 29428 37390
rect 29148 37324 29316 37380
rect 28924 36204 29014 36260
rect 28958 35736 29014 36204
rect 28700 35698 28756 35710
rect 28700 35646 28702 35698
rect 28754 35646 28756 35698
rect 28700 34916 28756 35646
rect 28812 35698 28868 35710
rect 28812 35646 28814 35698
rect 28866 35646 28868 35698
rect 28812 35252 28868 35646
rect 28958 35684 28960 35736
rect 29012 35684 29014 35736
rect 28958 35364 29014 35684
rect 28958 35298 29014 35308
rect 28812 35186 28868 35196
rect 29260 35026 29316 37324
rect 29372 35586 29428 37324
rect 29372 35534 29374 35586
rect 29426 35534 29428 35586
rect 29372 35522 29428 35534
rect 29820 35698 29876 35710
rect 29820 35646 29822 35698
rect 29874 35646 29876 35698
rect 29260 34974 29262 35026
rect 29314 34974 29316 35026
rect 29260 34962 29316 34974
rect 29596 35252 29652 35262
rect 28700 34850 28756 34860
rect 29148 34916 29204 34926
rect 29148 34822 29204 34860
rect 29596 34858 29652 35196
rect 29596 34806 29598 34858
rect 29650 34806 29652 34858
rect 29372 34692 29428 34702
rect 29260 34356 29316 34366
rect 28588 32510 28590 32562
rect 28642 32510 28644 32562
rect 28364 31892 28420 31902
rect 28364 31778 28420 31836
rect 28588 31892 28644 32510
rect 28588 31826 28644 31836
rect 28700 33348 28756 33358
rect 28364 31726 28366 31778
rect 28418 31726 28420 31778
rect 28364 31714 28420 31726
rect 28196 31556 28252 31566
rect 28196 31462 28252 31500
rect 27132 31054 27134 31106
rect 27186 31054 27188 31106
rect 27132 31042 27188 31054
rect 27468 31164 28084 31220
rect 26460 30212 26516 30998
rect 27132 30436 27188 30446
rect 27468 30436 27524 31164
rect 28140 31050 28196 31062
rect 26460 30194 26572 30212
rect 26460 30156 26518 30194
rect 26516 30142 26518 30156
rect 26570 30142 26572 30194
rect 27132 30182 27188 30380
rect 26516 30130 26572 30142
rect 26684 30154 26740 30166
rect 26684 30102 26686 30154
rect 26738 30102 26740 30154
rect 26684 29988 26740 30102
rect 26908 30154 26964 30166
rect 26908 30102 26910 30154
rect 26962 30102 26964 30154
rect 26908 30100 26964 30102
rect 26908 30034 26964 30044
rect 27132 30130 27134 30182
rect 27186 30130 27188 30182
rect 27412 30380 27524 30436
rect 27580 30996 27636 31006
rect 27412 30210 27468 30380
rect 27412 30158 27414 30210
rect 27466 30158 27468 30210
rect 27412 30146 27468 30158
rect 26684 29922 26740 29932
rect 26908 29428 26964 29438
rect 26908 29426 27076 29428
rect 26908 29374 26910 29426
rect 26962 29374 27076 29426
rect 26908 29372 27076 29374
rect 26908 29362 26964 29372
rect 26460 28642 26516 28654
rect 26460 28590 26462 28642
rect 26514 28590 26516 28642
rect 25676 27694 25678 27746
rect 25730 27694 25732 27746
rect 25676 27682 25732 27694
rect 25900 27885 25956 27897
rect 25900 27833 25902 27885
rect 25954 27833 25956 27885
rect 25900 27748 25956 27833
rect 25900 27682 25956 27692
rect 26236 27860 26292 27870
rect 26460 27860 26516 28590
rect 27020 28644 27076 29372
rect 27132 28980 27188 30130
rect 27244 29204 27300 29214
rect 27580 29204 27636 30940
rect 28140 30998 28142 31050
rect 28194 30998 28196 31050
rect 28140 30100 28196 30998
rect 28476 31050 28532 31062
rect 28476 30998 28478 31050
rect 28530 30998 28532 31050
rect 28476 30436 28532 30998
rect 28700 30996 28756 33292
rect 28700 30930 28756 30940
rect 29148 31750 29204 31762
rect 29148 31698 29150 31750
rect 29202 31698 29204 31750
rect 29148 31556 29204 31698
rect 28476 30370 28532 30380
rect 29148 30324 29204 31500
rect 29148 30258 29204 30268
rect 27804 29204 27860 29214
rect 27244 29202 27860 29204
rect 27244 29150 27246 29202
rect 27298 29150 27806 29202
rect 27858 29150 27860 29202
rect 27244 29148 27860 29150
rect 27244 29138 27300 29148
rect 27804 29138 27860 29148
rect 27132 28924 27300 28980
rect 27244 28810 27300 28924
rect 27244 28758 27246 28810
rect 27298 28758 27300 28810
rect 27244 28746 27300 28758
rect 27020 28550 27076 28588
rect 26236 27858 26516 27860
rect 26236 27806 26238 27858
rect 26290 27806 26516 27858
rect 26236 27804 26516 27806
rect 26572 27860 26628 27870
rect 26236 26964 26292 27804
rect 26572 27766 26628 27804
rect 28140 27242 28196 30044
rect 29260 29986 29316 34300
rect 29372 33514 29428 34636
rect 29372 33462 29374 33514
rect 29426 33462 29428 33514
rect 29372 33450 29428 33462
rect 29484 33348 29540 33358
rect 29484 33254 29540 33292
rect 29372 32564 29428 32574
rect 29596 32564 29652 34806
rect 29820 34914 29876 35646
rect 29932 35530 29988 37996
rect 30156 37828 30212 37838
rect 30156 37734 30212 37772
rect 32508 37380 32564 39566
rect 35980 38836 36036 40124
rect 36148 39396 36204 39406
rect 36540 39396 36596 40236
rect 37100 40290 37156 40302
rect 37100 40238 37102 40290
rect 37154 40238 37156 40290
rect 37100 39844 37156 40238
rect 37212 39844 37268 39854
rect 37100 39842 37268 39844
rect 37100 39790 37214 39842
rect 37266 39790 37268 39842
rect 37100 39788 37268 39790
rect 37212 39778 37268 39788
rect 36876 39620 36932 39630
rect 36148 39394 36596 39396
rect 36148 39342 36150 39394
rect 36202 39342 36596 39394
rect 36148 39340 36596 39342
rect 36148 39330 36204 39340
rect 36390 38871 36446 38883
rect 36092 38836 36148 38846
rect 35980 38834 36148 38836
rect 35980 38782 36094 38834
rect 36146 38782 36148 38834
rect 35980 38780 36148 38782
rect 36092 38770 36148 38780
rect 36204 38834 36260 38846
rect 36204 38782 36206 38834
rect 36258 38782 36260 38834
rect 35812 38724 35868 38734
rect 35812 38630 35868 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 32508 37314 32564 37324
rect 32956 37828 33012 37838
rect 32956 36594 33012 37772
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 32956 36542 32958 36594
rect 33010 36542 33012 36594
rect 32956 36530 33012 36542
rect 33740 36482 33796 36494
rect 33740 36430 33742 36482
rect 33794 36430 33796 36482
rect 31052 36372 31108 36382
rect 30828 36370 31108 36372
rect 30828 36318 31054 36370
rect 31106 36318 31108 36370
rect 30828 36316 31108 36318
rect 29932 35478 29934 35530
rect 29986 35478 29988 35530
rect 29932 35466 29988 35478
rect 30156 35698 30212 35710
rect 30156 35646 30158 35698
rect 30210 35646 30212 35698
rect 29820 34862 29822 34914
rect 29874 34862 29876 34914
rect 29820 34356 29876 34862
rect 29820 34290 29876 34300
rect 30156 34914 30212 35646
rect 30156 34862 30158 34914
rect 30210 34862 30212 34914
rect 30156 34804 30212 34862
rect 30156 34242 30212 34748
rect 30156 34190 30158 34242
rect 30210 34190 30212 34242
rect 30156 34178 30212 34190
rect 30828 34186 30884 36316
rect 31052 36306 31108 36316
rect 33740 36260 33796 36430
rect 34132 36260 34188 36270
rect 33740 36194 33796 36204
rect 34076 36204 34132 36260
rect 34076 36166 34188 36204
rect 33964 35700 34020 35710
rect 34076 35700 34132 36166
rect 33964 35698 34132 35700
rect 33964 35646 33966 35698
rect 34018 35646 34132 35698
rect 33964 35644 34132 35646
rect 33964 35634 34020 35644
rect 30604 34158 30660 34170
rect 30604 34106 30606 34158
rect 30658 34106 30660 34158
rect 30828 34134 30830 34186
rect 30882 34134 30884 34186
rect 30828 34122 30884 34134
rect 29988 34074 30044 34086
rect 29988 34022 29990 34074
rect 30042 34022 30044 34074
rect 29988 33908 30044 34022
rect 29988 33842 30044 33852
rect 30604 33460 30660 34106
rect 30604 33394 30660 33404
rect 32508 33908 32564 33918
rect 29820 33348 29876 33358
rect 29820 33254 29876 33292
rect 31276 33348 31332 33358
rect 31276 32674 31332 33292
rect 32508 33346 32564 33852
rect 32508 33294 32510 33346
rect 32562 33294 32564 33346
rect 32508 33282 32564 33294
rect 31276 32622 31278 32674
rect 31330 32622 31332 32674
rect 31276 32610 31332 32622
rect 32844 33122 32900 33134
rect 32844 33070 32846 33122
rect 32898 33070 32900 33122
rect 29372 32562 29652 32564
rect 29372 32510 29374 32562
rect 29426 32510 29652 32562
rect 29372 32508 29652 32510
rect 29372 32498 29428 32508
rect 31892 32450 31948 32462
rect 31892 32398 31894 32450
rect 31946 32398 31948 32450
rect 31892 32116 31948 32398
rect 31836 32060 31948 32116
rect 30492 32002 30548 32014
rect 30492 31950 30494 32002
rect 30546 31950 30548 32002
rect 30492 31948 30548 31950
rect 30156 31892 30548 31948
rect 31836 31892 31892 32060
rect 32844 32004 32900 33070
rect 32844 31938 32900 31948
rect 30156 31826 30212 31836
rect 31836 31826 31892 31836
rect 33460 31892 33516 31902
rect 33516 31836 33684 31892
rect 33460 31798 33516 31836
rect 33628 31778 33684 31836
rect 33628 31726 33630 31778
rect 33682 31726 33684 31778
rect 33628 31714 33684 31726
rect 32564 31556 32620 31566
rect 32564 31218 32620 31500
rect 32564 31166 32566 31218
rect 32618 31166 32620 31218
rect 32564 31154 32620 31166
rect 33068 31556 33124 31566
rect 33068 31021 33124 31500
rect 33068 30969 33070 31021
rect 33122 30969 33124 31021
rect 33068 30957 33124 30969
rect 34076 30882 34132 35644
rect 34748 35586 34804 35598
rect 34748 35534 34750 35586
rect 34802 35534 34804 35586
rect 34748 34244 34804 35534
rect 36204 35364 36260 38782
rect 36390 38819 36392 38871
rect 36444 38819 36446 38871
rect 36390 38724 36446 38819
rect 36390 38388 36446 38668
rect 36390 38332 36484 38388
rect 36428 36036 36484 38332
rect 36540 36260 36596 39340
rect 36764 39618 36932 39620
rect 36764 39566 36878 39618
rect 36930 39566 36932 39618
rect 36764 39564 36932 39566
rect 36764 38722 36820 39564
rect 36876 39554 36932 39564
rect 39340 39620 39396 39630
rect 36764 38670 36766 38722
rect 36818 38670 36820 38722
rect 36764 38658 36820 38670
rect 39340 38668 39396 39564
rect 40348 38668 40404 40338
rect 41580 40292 41636 40302
rect 41020 40290 41636 40292
rect 41020 40238 41582 40290
rect 41634 40238 41636 40290
rect 41020 40236 41636 40238
rect 41020 39842 41076 40236
rect 41580 40226 41636 40236
rect 41020 39790 41022 39842
rect 41074 39790 41076 39842
rect 41020 39778 41076 39790
rect 41804 39844 41860 41106
rect 43484 40290 43540 40302
rect 43484 40238 43486 40290
rect 43538 40238 43540 40290
rect 41804 39778 41860 39788
rect 42588 39844 42644 39854
rect 42588 39750 42644 39788
rect 39228 38612 39396 38668
rect 39676 38612 40404 38668
rect 40684 39618 40740 39630
rect 40684 39566 40686 39618
rect 40738 39566 40740 39618
rect 36540 36194 36596 36204
rect 37156 36260 37212 36270
rect 37156 36166 37212 36204
rect 36428 35980 36596 36036
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35756 35308 36260 35364
rect 36428 35700 36484 35710
rect 34748 34178 34804 34188
rect 35644 34158 35700 34170
rect 35644 34106 35646 34158
rect 35698 34106 35700 34158
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34636 32004 34692 32014
rect 34412 31778 34468 31790
rect 34412 31726 34414 31778
rect 34466 31726 34468 31778
rect 34412 31108 34468 31726
rect 34412 31042 34468 31052
rect 34076 30830 34078 30882
rect 34130 30830 34132 30882
rect 29260 29934 29262 29986
rect 29314 29934 29316 29986
rect 29260 29922 29316 29934
rect 29820 29986 29876 29998
rect 29820 29934 29822 29986
rect 29874 29934 29876 29986
rect 29036 29204 29092 29214
rect 29036 29202 29204 29204
rect 29036 29150 29038 29202
rect 29090 29150 29204 29202
rect 29036 29148 29204 29150
rect 29036 29138 29092 29148
rect 29148 28642 29204 29148
rect 29820 28878 29876 29934
rect 33628 29426 33684 29438
rect 33628 29374 33630 29426
rect 33682 29374 33684 29426
rect 33292 29202 33348 29214
rect 33292 29150 33294 29202
rect 33346 29150 33348 29202
rect 29820 28866 29932 28878
rect 29820 28814 29878 28866
rect 29930 28814 29932 28866
rect 29820 28812 29932 28814
rect 29876 28802 29932 28812
rect 31388 28868 31444 28878
rect 29148 28590 29150 28642
rect 29202 28590 29204 28642
rect 29596 28642 29652 28654
rect 29148 28578 29204 28590
rect 29316 28586 29372 28598
rect 29316 28534 29318 28586
rect 29370 28534 29372 28586
rect 29596 28590 29598 28642
rect 29650 28590 29652 28642
rect 29316 28084 29372 28534
rect 29148 28028 29372 28084
rect 29484 28530 29540 28542
rect 29484 28478 29486 28530
rect 29538 28478 29540 28530
rect 29484 28084 29540 28478
rect 29596 28196 29652 28590
rect 31388 28642 31444 28812
rect 33292 28754 33348 29150
rect 33628 29204 33684 29374
rect 33964 29204 34020 29214
rect 33628 29202 34020 29204
rect 33628 29150 33966 29202
rect 34018 29150 34020 29202
rect 33628 29148 34020 29150
rect 33964 29138 34020 29148
rect 33292 28702 33294 28754
rect 33346 28702 33348 28754
rect 33292 28690 33348 28702
rect 31388 28590 31390 28642
rect 31442 28590 31444 28642
rect 29596 28140 29876 28196
rect 29820 28084 29876 28140
rect 29484 28028 29764 28084
rect 29820 28028 29988 28084
rect 28140 27190 28142 27242
rect 28194 27190 28196 27242
rect 28140 27178 28196 27190
rect 28924 27858 28980 27870
rect 28924 27806 28926 27858
rect 28978 27806 28980 27858
rect 28252 27076 28308 27086
rect 28252 26982 28308 27020
rect 28588 27076 28644 27086
rect 28924 27076 28980 27806
rect 29036 27860 29092 27870
rect 29148 27860 29204 28028
rect 29092 27804 29204 27860
rect 29260 27858 29316 27870
rect 29260 27806 29262 27858
rect 29314 27806 29316 27858
rect 29036 27690 29092 27804
rect 29036 27638 29038 27690
rect 29090 27638 29092 27690
rect 29036 27626 29092 27638
rect 29260 27300 29316 27806
rect 29708 27690 29764 28028
rect 29708 27638 29710 27690
rect 29762 27638 29764 27690
rect 29708 27626 29764 27638
rect 29820 27858 29876 27870
rect 29820 27806 29822 27858
rect 29874 27806 29876 27858
rect 29820 27300 29876 27806
rect 29260 27244 29876 27300
rect 28588 27074 28980 27076
rect 28588 27022 28590 27074
rect 28642 27022 28980 27074
rect 28588 27020 28980 27022
rect 29596 27074 29652 27086
rect 29596 27022 29598 27074
rect 29650 27022 29652 27074
rect 28588 27010 28644 27020
rect 26236 26898 26292 26908
rect 28364 26964 28420 26974
rect 24276 26178 25060 26180
rect 24276 26126 24278 26178
rect 24330 26126 25060 26178
rect 24276 26124 25060 26126
rect 24276 26114 24332 26124
rect 24108 25778 24164 25788
rect 24108 25620 24164 25630
rect 24108 25618 24948 25620
rect 24108 25566 24110 25618
rect 24162 25566 24948 25618
rect 24108 25564 24948 25566
rect 24108 25554 24164 25564
rect 24892 25506 24948 25564
rect 24892 25454 24894 25506
rect 24946 25454 24948 25506
rect 24892 25442 24948 25454
rect 25004 25506 25060 26124
rect 25004 25454 25006 25506
rect 25058 25454 25060 25506
rect 25172 26124 25284 26180
rect 28252 26740 28308 26750
rect 28252 26290 28308 26684
rect 28252 26238 28254 26290
rect 28306 26238 28308 26290
rect 25172 25562 25228 26124
rect 25172 25510 25174 25562
rect 25226 25510 25228 25562
rect 25172 25498 25228 25510
rect 25340 25506 25396 25518
rect 25004 25442 25060 25454
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 24612 25396 24668 25406
rect 23996 25394 24668 25396
rect 23996 25342 24614 25394
rect 24666 25342 24668 25394
rect 23996 25340 24668 25342
rect 24612 25330 24668 25340
rect 25340 25396 25396 25454
rect 25340 25330 25396 25340
rect 25844 25396 25900 25406
rect 25844 25302 25900 25340
rect 23772 25004 23920 25060
rect 24108 25172 24164 25182
rect 23436 24948 23492 24958
rect 23436 24854 23492 24892
rect 23772 24948 23828 25004
rect 22932 24724 22988 24734
rect 23100 24724 23156 24734
rect 22988 24722 23156 24724
rect 22988 24670 23102 24722
rect 23154 24670 23156 24722
rect 22988 24668 23156 24670
rect 22932 24630 22988 24668
rect 23100 24658 23156 24668
rect 23772 24722 23828 24892
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 23772 24658 23828 24670
rect 23940 24500 23996 24510
rect 22764 24444 22988 24500
rect 22932 24050 22988 24444
rect 22932 23998 22934 24050
rect 22986 23998 22988 24050
rect 22932 23940 22988 23998
rect 23772 24498 24052 24500
rect 23772 24446 23942 24498
rect 23994 24446 24052 24498
rect 23772 24444 24052 24446
rect 22932 23874 22988 23884
rect 23548 23940 23604 23950
rect 23548 23846 23604 23884
rect 23772 23938 23828 24444
rect 23940 24434 24052 24444
rect 23772 23886 23774 23938
rect 23826 23886 23828 23938
rect 23996 23994 24052 24434
rect 23996 23942 23998 23994
rect 24050 23942 24052 23994
rect 23996 23930 24052 23942
rect 23772 23874 23828 23886
rect 24108 23900 24164 25116
rect 25284 24500 25340 24510
rect 25284 24052 25340 24444
rect 24108 23848 24110 23900
rect 24162 23848 24164 23900
rect 23268 23826 23324 23838
rect 24108 23836 24164 23848
rect 24836 24050 25340 24052
rect 24836 23998 25286 24050
rect 25338 23998 25340 24050
rect 24836 23996 25340 23998
rect 24836 23994 24892 23996
rect 24836 23942 24838 23994
rect 24890 23942 24892 23994
rect 25284 23986 25340 23996
rect 24668 23828 24724 23838
rect 23268 23774 23270 23826
rect 23322 23774 23324 23826
rect 23268 23268 23324 23774
rect 24556 23826 24724 23828
rect 24556 23774 24670 23826
rect 24722 23774 24724 23826
rect 24556 23772 24724 23774
rect 23268 23202 23324 23212
rect 23772 23268 23828 23278
rect 22652 22932 22708 22942
rect 22428 22930 22708 22932
rect 22428 22878 22654 22930
rect 22706 22878 22708 22930
rect 22428 22876 22708 22878
rect 21868 20862 21870 20914
rect 21922 20862 21924 20914
rect 21868 20132 21924 20862
rect 21868 20066 21924 20076
rect 21588 18340 21644 18350
rect 21532 18284 21588 18340
rect 21532 18246 21644 18284
rect 21364 17892 21420 17902
rect 21364 17798 21420 17836
rect 21196 16882 21252 17052
rect 20468 16660 20524 16670
rect 20188 16658 20524 16660
rect 20188 16606 20470 16658
rect 20522 16606 20524 16658
rect 20188 16604 20524 16606
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 15708 15474 15764 15484
rect 17556 15538 17668 15550
rect 17556 15486 17558 15538
rect 17610 15486 17668 15538
rect 17556 15484 17668 15486
rect 14812 15262 14814 15314
rect 14866 15262 14868 15314
rect 14812 15250 14868 15262
rect 14700 15204 14756 15214
rect 14700 14644 14756 15148
rect 14700 14502 14756 14588
rect 14700 14450 14702 14502
rect 14754 14450 14756 14502
rect 14700 14438 14756 14450
rect 15036 15204 15092 15214
rect 14476 13794 14532 13804
rect 14812 13914 14868 13926
rect 14812 13862 14814 13914
rect 14866 13862 14868 13914
rect 13692 13694 13694 13746
rect 13746 13694 13748 13746
rect 13692 13682 13748 13694
rect 13860 13746 13916 13758
rect 13860 13694 13862 13746
rect 13914 13694 13916 13746
rect 13860 13636 13916 13694
rect 13860 13570 13916 13580
rect 14028 13748 14084 13758
rect 14028 13412 14084 13692
rect 14700 13748 14756 13758
rect 14700 13654 14756 13692
rect 14364 13636 14420 13646
rect 14252 13524 14308 13534
rect 14252 13430 14308 13468
rect 13524 13186 13636 13198
rect 13524 13134 13526 13186
rect 13578 13134 13636 13186
rect 13524 13132 13636 13134
rect 13692 13356 14084 13412
rect 13524 13122 13580 13132
rect 12908 12910 12910 12962
rect 12962 12910 12964 12962
rect 12908 12898 12964 12910
rect 13692 12962 13748 13356
rect 13692 12910 13694 12962
rect 13746 12910 13748 12962
rect 13692 12898 13748 12910
rect 14084 12740 14140 12750
rect 13692 12738 14140 12740
rect 13692 12686 14086 12738
rect 14138 12686 14140 12738
rect 13692 12684 14140 12686
rect 12796 12014 12798 12066
rect 12850 12014 12852 12066
rect 12796 12002 12852 12014
rect 12908 12205 12964 12217
rect 12908 12153 12910 12205
rect 12962 12153 12964 12205
rect 12908 11508 12964 12153
rect 13244 12180 13300 12190
rect 13244 12086 13300 12124
rect 13580 12180 13636 12190
rect 13580 12086 13636 12124
rect 12908 11442 12964 11452
rect 12572 11228 13020 11284
rect 12964 10834 13020 11228
rect 12964 10782 12966 10834
rect 13018 10782 13020 10834
rect 12964 10770 13020 10782
rect 12684 10612 12740 10622
rect 12460 10610 12740 10612
rect 12460 10558 12686 10610
rect 12738 10558 12740 10610
rect 12460 10556 12740 10558
rect 12348 10386 12404 10398
rect 12348 10334 12350 10386
rect 12402 10334 12404 10386
rect 12348 9380 12404 10334
rect 12348 9314 12404 9324
rect 12460 9268 12516 10556
rect 12684 10546 12740 10556
rect 13132 10610 13188 10622
rect 13132 10558 13134 10610
rect 13186 10558 13188 10610
rect 13132 9940 13188 10558
rect 13132 9874 13188 9884
rect 13468 9940 13524 9950
rect 12460 9202 12516 9212
rect 11004 8372 11228 8428
rect 12124 8372 12292 8428
rect 12348 9156 12404 9166
rect 12348 9098 12404 9100
rect 12348 9046 12350 9098
rect 12402 9046 12404 9098
rect 13300 9156 13356 9166
rect 13300 9098 13356 9100
rect 12348 8428 12404 9046
rect 12796 9044 12852 9054
rect 13132 9044 13188 9054
rect 12796 9042 13188 9044
rect 12796 8990 12798 9042
rect 12850 8990 13134 9042
rect 13186 8990 13188 9042
rect 13300 9046 13302 9098
rect 13354 9046 13356 9098
rect 13468 9154 13524 9884
rect 13468 9102 13470 9154
rect 13522 9102 13524 9154
rect 13468 9090 13524 9102
rect 13580 9268 13636 9278
rect 13300 9034 13356 9046
rect 13580 9042 13636 9212
rect 12796 8988 13188 8990
rect 12796 8978 12852 8988
rect 12572 8930 12628 8942
rect 12572 8878 12574 8930
rect 12626 8878 12628 8930
rect 12348 8372 12516 8428
rect 9660 8194 9716 8204
rect 10668 8260 10724 8270
rect 10668 8166 10724 8204
rect 11004 8243 11060 8372
rect 11004 8191 11006 8243
rect 11058 8191 11060 8243
rect 11004 8179 11060 8191
rect 10892 8090 10948 8102
rect 10892 8038 10894 8090
rect 10946 8038 10948 8090
rect 8204 7196 8428 7252
rect 8372 6746 8428 7196
rect 7980 6692 8036 6702
rect 7644 6600 7646 6652
rect 7698 6600 7700 6652
rect 7644 5684 7700 6600
rect 7756 6690 8036 6692
rect 7756 6638 7982 6690
rect 8034 6638 8036 6690
rect 8372 6694 8374 6746
rect 8426 6694 8428 6746
rect 8372 6682 8428 6694
rect 7756 6636 8036 6638
rect 7756 5908 7812 6636
rect 7980 6626 8036 6636
rect 8204 6578 8260 6590
rect 8204 6526 8206 6578
rect 8258 6526 8260 6578
rect 8204 6244 8260 6526
rect 8204 6188 8708 6244
rect 7756 5814 7812 5852
rect 7868 5906 7924 5918
rect 7868 5854 7870 5906
rect 7922 5854 7924 5906
rect 7868 5684 7924 5854
rect 8148 5908 8204 5918
rect 8428 5908 8484 5918
rect 8148 5906 8484 5908
rect 8148 5854 8150 5906
rect 8202 5854 8430 5906
rect 8482 5854 8484 5906
rect 8148 5852 8484 5854
rect 8148 5842 8204 5852
rect 8428 5842 8484 5852
rect 8652 5906 8708 6188
rect 8652 5854 8654 5906
rect 8706 5854 8708 5906
rect 8652 5842 8708 5854
rect 9604 5908 9660 5918
rect 9212 5796 9268 5806
rect 7644 5628 7924 5684
rect 8428 5684 8484 5694
rect 5852 5058 5908 5068
rect 6524 5124 6580 5134
rect 6524 5030 6580 5068
rect 7308 5124 7364 5134
rect 7308 5122 7588 5124
rect 7308 5070 7310 5122
rect 7362 5070 7588 5122
rect 7308 5068 7588 5070
rect 7308 5058 7364 5068
rect 7532 4562 7588 5068
rect 8428 4900 8484 5628
rect 8932 5684 8988 5694
rect 8932 5590 8988 5628
rect 9212 5234 9268 5740
rect 9604 5738 9660 5852
rect 9772 5908 9828 5918
rect 9772 5814 9828 5852
rect 9604 5686 9606 5738
rect 9658 5686 9660 5738
rect 9604 5674 9660 5686
rect 9212 5182 9214 5234
rect 9266 5182 9268 5234
rect 9212 5170 9268 5182
rect 9828 5236 9884 5246
rect 9828 5142 9884 5180
rect 10108 5236 10164 5246
rect 10108 5122 10164 5180
rect 10892 5234 10948 8038
rect 12124 6074 12180 8372
rect 12460 6692 12516 8372
rect 12572 7588 12628 8878
rect 12572 7522 12628 7532
rect 12684 6692 12740 6702
rect 13020 6692 13076 6702
rect 12460 6690 12740 6692
rect 12460 6638 12686 6690
rect 12738 6638 12740 6690
rect 12460 6636 12740 6638
rect 12684 6626 12740 6636
rect 12796 6690 13076 6692
rect 12796 6638 13022 6690
rect 13074 6638 13076 6690
rect 12796 6636 13076 6638
rect 12124 6022 12126 6074
rect 12178 6022 12180 6074
rect 12124 6010 12180 6022
rect 12460 5945 12516 5957
rect 12012 5908 12068 5918
rect 12012 5814 12068 5852
rect 12460 5908 12462 5945
rect 12514 5908 12516 5945
rect 12460 5842 12516 5852
rect 12684 5908 12740 5918
rect 12796 5908 12852 6636
rect 13020 6626 13076 6636
rect 12684 5906 12852 5908
rect 12684 5854 12686 5906
rect 12738 5854 12852 5906
rect 12684 5852 12852 5854
rect 12684 5842 12740 5852
rect 10892 5182 10894 5234
rect 10946 5182 10948 5234
rect 10892 5170 10948 5182
rect 12796 5234 12852 5852
rect 13132 5908 13188 8988
rect 13580 8990 13582 9042
rect 13634 8990 13636 9042
rect 13580 8978 13636 8990
rect 13692 8428 13748 12684
rect 14084 12674 14140 12684
rect 14364 10164 14420 13580
rect 14812 12180 14868 13862
rect 15036 13790 15092 15148
rect 16716 15204 16772 15214
rect 17556 15148 17612 15484
rect 16716 15110 16772 15148
rect 17500 15092 17612 15148
rect 15372 14868 15428 14878
rect 15372 14754 15428 14812
rect 15372 14702 15374 14754
rect 15426 14702 15428 14754
rect 15372 14690 15428 14702
rect 17500 14868 17556 15092
rect 17332 14644 17388 14654
rect 17332 14550 17388 14588
rect 15036 13738 15038 13790
rect 15090 13738 15092 13790
rect 15036 13726 15092 13738
rect 15652 13972 15708 13982
rect 15652 13524 15708 13916
rect 15652 13458 15708 13468
rect 17500 13086 17556 14812
rect 19628 14308 19684 14318
rect 19628 13792 19684 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 16604
rect 20468 16594 20524 16604
rect 20860 16324 20916 16830
rect 21196 16830 21198 16882
rect 21250 16830 21252 16882
rect 21196 16818 21252 16830
rect 21532 16324 21588 18246
rect 21644 17666 21700 17678
rect 21644 17614 21646 17666
rect 21698 17614 21700 17666
rect 21644 17332 21700 17614
rect 21868 17668 21924 17678
rect 21868 17574 21924 17612
rect 22260 17668 22316 17678
rect 22260 17574 22316 17612
rect 21644 17276 21924 17332
rect 21700 17108 21756 17118
rect 21700 17014 21756 17052
rect 21756 16884 21812 16894
rect 21868 16884 21924 17276
rect 22204 17108 22260 17118
rect 22204 17014 22260 17052
rect 21812 16882 21924 16884
rect 21812 16830 21870 16882
rect 21922 16830 21924 16882
rect 21812 16828 21924 16830
rect 20860 16268 21476 16324
rect 21420 16110 21476 16268
rect 21588 16268 21700 16324
rect 21532 16258 21588 16268
rect 21420 16098 21532 16110
rect 21420 16046 21478 16098
rect 21530 16046 21532 16098
rect 21420 16044 21532 16046
rect 21476 16034 21532 16044
rect 20356 14308 20412 14318
rect 20356 14214 20412 14252
rect 20188 13906 20244 13916
rect 20300 13860 20356 13870
rect 19740 13792 19796 13802
rect 19628 13790 19796 13792
rect 19628 13738 19742 13790
rect 19794 13738 19796 13790
rect 19628 13736 19796 13738
rect 19740 13726 19796 13736
rect 20076 13748 20132 13758
rect 20076 13654 20132 13692
rect 20300 13746 20356 13804
rect 21084 13860 21140 13870
rect 20300 13694 20302 13746
rect 20354 13694 20356 13746
rect 19628 13636 19684 13646
rect 18508 13634 19684 13636
rect 18508 13582 19630 13634
rect 19682 13582 19684 13634
rect 18508 13580 19684 13582
rect 17500 13076 17612 13086
rect 17500 13074 17780 13076
rect 17500 13022 17558 13074
rect 17610 13022 17780 13074
rect 17500 13020 17780 13022
rect 17500 13010 17612 13020
rect 16884 12180 16940 12190
rect 17388 12180 17444 12190
rect 17500 12180 17556 13010
rect 17724 12962 17780 13020
rect 18508 13074 18564 13580
rect 19628 13570 19684 13580
rect 20300 13524 20356 13694
rect 18508 13022 18510 13074
rect 18562 13022 18564 13074
rect 18508 13010 18564 13022
rect 20076 13468 20356 13524
rect 20524 13748 20580 13758
rect 17724 12910 17726 12962
rect 17778 12910 17780 12962
rect 17724 12898 17780 12910
rect 20076 12740 20132 13468
rect 20412 13076 20468 13086
rect 20524 13076 20580 13692
rect 21084 13746 21140 13804
rect 21084 13694 21086 13746
rect 21138 13694 21140 13746
rect 21084 13682 21140 13694
rect 21308 13748 21364 13758
rect 21308 13654 21364 13692
rect 21644 13748 21700 16268
rect 21644 13682 21700 13692
rect 20804 13524 20860 13534
rect 21588 13524 21644 13534
rect 20412 13074 20580 13076
rect 20412 13022 20414 13074
rect 20466 13022 20580 13074
rect 20412 13020 20580 13022
rect 20636 13522 21364 13524
rect 20636 13470 20806 13522
rect 20858 13470 21364 13522
rect 20636 13468 21364 13470
rect 20412 13010 20468 13020
rect 20076 12684 20244 12740
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20188 12404 20244 12684
rect 20076 12348 20244 12404
rect 20076 12290 20132 12348
rect 20076 12238 20078 12290
rect 20130 12238 20132 12290
rect 20076 12226 20132 12238
rect 14812 12114 14868 12124
rect 16828 12178 17556 12180
rect 16828 12126 16886 12178
rect 16938 12126 17390 12178
rect 17442 12126 17556 12178
rect 16828 12124 17556 12126
rect 20636 12178 20692 13468
rect 20804 13458 20860 13468
rect 21308 12962 21364 13468
rect 21308 12910 21310 12962
rect 21362 12910 21364 12962
rect 21308 12898 21364 12910
rect 21420 13522 21644 13524
rect 21420 13470 21590 13522
rect 21642 13470 21644 13522
rect 21420 13468 21644 13470
rect 21420 12404 21476 13468
rect 21588 13458 21644 13468
rect 20636 12126 20638 12178
rect 20690 12126 20692 12178
rect 16828 12114 16940 12124
rect 17388 12114 17444 12124
rect 20636 12114 20692 12126
rect 20748 12348 21476 12404
rect 21532 13300 21588 13310
rect 21756 13300 21812 16828
rect 21868 16818 21924 16828
rect 22652 16212 22708 22876
rect 23772 22370 23828 23212
rect 24556 23044 24612 23772
rect 24668 23762 24724 23772
rect 24836 23380 24892 23942
rect 28252 23940 28308 26238
rect 28364 26178 28420 26908
rect 28364 26126 28366 26178
rect 28418 26126 28420 26178
rect 28364 26114 28420 26126
rect 28588 26317 28644 26329
rect 28588 26265 28590 26317
rect 28642 26265 28644 26317
rect 28588 26068 28644 26265
rect 28588 26002 28644 26012
rect 28700 25172 28756 27020
rect 28924 26292 28980 26302
rect 29484 26292 29540 26302
rect 28924 25732 28980 26236
rect 28924 25666 28980 25676
rect 29260 26290 29540 26292
rect 29260 26238 29486 26290
rect 29538 26238 29540 26290
rect 29260 26236 29540 26238
rect 29260 25508 29316 26236
rect 29484 26226 29540 26236
rect 29596 26292 29652 27022
rect 29708 26852 29764 27244
rect 29932 27186 29988 28028
rect 29932 27134 29934 27186
rect 29986 27134 29988 27186
rect 29932 27122 29988 27134
rect 30044 27858 30100 27870
rect 30044 27806 30046 27858
rect 30098 27806 30100 27858
rect 29932 27018 29988 27030
rect 29932 26966 29934 27018
rect 29986 26966 29988 27018
rect 29932 26964 29988 26966
rect 29932 26898 29988 26908
rect 29708 26786 29764 26796
rect 30044 26628 30100 27806
rect 30268 27074 30324 27086
rect 30268 27022 30270 27074
rect 30322 27022 30324 27074
rect 30268 26740 30324 27022
rect 30268 26674 30324 26684
rect 30492 26964 30548 26974
rect 30044 26572 30212 26628
rect 29596 26226 29652 26236
rect 30156 26068 30212 26572
rect 30360 26290 30416 26302
rect 30360 26238 30362 26290
rect 30414 26238 30416 26290
rect 30360 26180 30416 26238
rect 30360 26114 30416 26124
rect 30156 26002 30212 26012
rect 30492 25956 30548 26908
rect 30604 26852 30660 26862
rect 30604 26402 30660 26796
rect 30604 26350 30606 26402
rect 30658 26350 30660 26402
rect 30604 26338 30660 26350
rect 31220 26180 31276 26190
rect 31220 26086 31276 26124
rect 30380 25900 30548 25956
rect 30716 26068 30772 26078
rect 29708 25508 29764 25518
rect 29260 25506 29764 25508
rect 29260 25454 29710 25506
rect 29762 25454 29764 25506
rect 29260 25452 29764 25454
rect 28476 25116 28756 25172
rect 28252 23884 28420 23940
rect 23772 22318 23774 22370
rect 23826 22318 23828 22370
rect 23772 22306 23828 22318
rect 23996 22988 24612 23044
rect 24780 23324 24892 23380
rect 23996 22370 24052 22988
rect 23996 22318 23998 22370
rect 24050 22318 24052 22370
rect 23996 22306 24052 22318
rect 24276 22260 24332 22270
rect 24108 22258 24332 22260
rect 24108 22206 24278 22258
rect 24330 22206 24332 22258
rect 24108 22204 24332 22206
rect 24108 21924 24164 22204
rect 24276 22194 24332 22204
rect 23772 21868 24164 21924
rect 23772 21586 23828 21868
rect 23772 21534 23774 21586
rect 23826 21534 23828 21586
rect 23772 21522 23828 21534
rect 23436 21364 23492 21374
rect 23436 21362 23828 21364
rect 23436 21310 23438 21362
rect 23490 21310 23828 21362
rect 23436 21308 23828 21310
rect 23436 21298 23492 21308
rect 23772 20914 23828 21308
rect 23772 20862 23774 20914
rect 23826 20862 23828 20914
rect 23772 20850 23828 20862
rect 24556 20804 24612 20814
rect 24556 20710 24612 20748
rect 24780 20188 24836 23324
rect 27356 22370 27412 22382
rect 27356 22318 27358 22370
rect 27410 22318 27412 22370
rect 27356 22260 27412 22318
rect 27356 22194 27412 22204
rect 28232 22314 28288 22326
rect 28232 22262 28234 22314
rect 28286 22262 28288 22314
rect 28232 21812 28288 22262
rect 28364 22260 28420 23884
rect 28476 22594 28532 25116
rect 29708 24052 29764 25452
rect 28476 22542 28478 22594
rect 28530 22542 28532 22594
rect 28476 22530 28532 22542
rect 28588 23996 29764 24052
rect 28364 22194 28420 22204
rect 28232 21746 28288 21756
rect 24948 20804 25004 20814
rect 24948 20580 25004 20748
rect 24948 20578 25172 20580
rect 24948 20526 24950 20578
rect 25002 20526 25172 20578
rect 24948 20524 25172 20526
rect 24948 20514 25004 20524
rect 24780 20132 24948 20188
rect 24444 18340 24500 18350
rect 24444 17780 24500 18284
rect 22652 14644 22708 16156
rect 23884 16324 23940 16334
rect 23044 16100 23100 16110
rect 23212 16100 23268 16110
rect 23100 16098 23268 16100
rect 23100 16046 23214 16098
rect 23266 16046 23268 16098
rect 23100 16044 23268 16046
rect 23044 16006 23100 16044
rect 23212 16034 23268 16044
rect 23548 15874 23604 15886
rect 23548 15822 23550 15874
rect 23602 15822 23604 15874
rect 23548 15316 23604 15822
rect 23884 15538 23940 16268
rect 23884 15486 23886 15538
rect 23938 15486 23940 15538
rect 23884 15474 23940 15486
rect 23548 15222 23604 15260
rect 22652 14578 22708 14588
rect 24444 15202 24500 17724
rect 24892 16222 24948 20132
rect 25116 20020 25172 20524
rect 27804 20132 27860 20142
rect 27804 20038 27860 20076
rect 24892 16210 25004 16222
rect 24892 16158 24950 16210
rect 25002 16158 25004 16210
rect 24892 16146 25004 16158
rect 24780 15316 24836 15326
rect 24892 15316 24948 16146
rect 24780 15314 25060 15316
rect 24780 15262 24782 15314
rect 24834 15262 25060 15314
rect 24780 15260 25060 15262
rect 24780 15250 24836 15260
rect 24444 15150 24446 15202
rect 24498 15150 24500 15202
rect 24444 14532 24500 15150
rect 25004 15148 25060 15260
rect 25116 15314 25172 19964
rect 25900 19906 25956 19918
rect 25900 19854 25902 19906
rect 25954 19854 25956 19906
rect 25900 19458 25956 19854
rect 25900 19406 25902 19458
rect 25954 19406 25956 19458
rect 25900 19394 25956 19406
rect 28364 19796 28420 19806
rect 28588 19796 28644 23996
rect 30380 23266 30436 25900
rect 30584 25508 30640 25518
rect 30584 25414 30640 25452
rect 30380 23214 30382 23266
rect 30434 23214 30436 23266
rect 30380 23202 30436 23214
rect 29260 23156 29316 23166
rect 29036 23154 29316 23156
rect 29036 23102 29262 23154
rect 29314 23102 29316 23154
rect 29036 23100 29316 23102
rect 29036 22372 29092 23100
rect 29260 23090 29316 23100
rect 30136 23156 30192 23166
rect 30136 23062 30192 23100
rect 30492 22596 30548 22606
rect 30716 22596 30772 26012
rect 30828 25732 30884 25742
rect 30828 25638 30884 25676
rect 30492 22594 30772 22596
rect 30492 22542 30494 22594
rect 30546 22542 30772 22594
rect 30492 22540 30772 22542
rect 30492 22530 30548 22540
rect 29372 22372 29428 22382
rect 30248 22372 30304 22382
rect 29036 22370 29540 22372
rect 29036 22318 29374 22370
rect 29426 22318 29540 22370
rect 29036 22316 29540 22318
rect 29372 22306 29428 22316
rect 29036 21812 29092 21822
rect 28812 21700 28868 21710
rect 28812 21642 28868 21644
rect 28812 21590 28814 21642
rect 28866 21590 28868 21642
rect 28812 21578 28868 21590
rect 29036 21616 29092 21756
rect 29484 21698 29540 22316
rect 30248 22278 30304 22316
rect 29484 21646 29486 21698
rect 29538 21646 29540 21698
rect 29484 21634 29540 21646
rect 31276 22260 31332 22270
rect 29036 21564 29038 21616
rect 29090 21564 29092 21616
rect 29036 21028 29092 21564
rect 29204 21530 29260 21542
rect 29204 21478 29206 21530
rect 29258 21478 29260 21530
rect 29204 21028 29260 21478
rect 29540 21028 29596 21038
rect 29204 20972 29428 21028
rect 29036 20962 29092 20972
rect 29036 20802 29092 20814
rect 29036 20750 29038 20802
rect 29090 20750 29092 20802
rect 29036 20188 29092 20750
rect 29260 20804 29316 20814
rect 29260 20710 29316 20748
rect 28700 20132 29092 20188
rect 29372 20188 29428 20972
rect 29540 20934 29596 20972
rect 29372 20132 29652 20188
rect 28700 20018 28756 20076
rect 29092 20020 29148 20030
rect 28700 19966 28702 20018
rect 28754 19966 28756 20018
rect 28700 19954 28756 19966
rect 29036 19964 29092 20020
rect 28364 19794 28644 19796
rect 28364 19742 28366 19794
rect 28418 19742 28644 19794
rect 28364 19740 28644 19742
rect 29036 19926 29148 19964
rect 26236 19234 26292 19246
rect 26236 19182 26238 19234
rect 26290 19182 26292 19234
rect 26236 18900 26292 19182
rect 26236 18844 26628 18900
rect 26572 18618 26628 18844
rect 26572 18566 26574 18618
rect 26626 18566 26628 18618
rect 28140 18676 28196 18686
rect 26572 18554 26628 18566
rect 26908 18564 26964 18574
rect 26908 18506 26964 18508
rect 26460 18450 26516 18462
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 26908 18454 26910 18506
rect 26962 18454 26964 18506
rect 27692 18564 27748 18574
rect 26908 18442 26964 18454
rect 27132 18450 27188 18462
rect 26180 18340 26236 18350
rect 26180 18246 26236 18284
rect 26460 18340 26516 18398
rect 26460 18274 26516 18284
rect 27132 18398 27134 18450
rect 27186 18398 27188 18450
rect 27132 18340 27188 18398
rect 27132 18274 27188 18284
rect 27692 18338 27748 18508
rect 27692 18286 27694 18338
rect 27746 18286 27748 18338
rect 27692 18274 27748 18286
rect 27804 18465 27860 18477
rect 27804 18452 27806 18465
rect 27858 18452 27860 18465
rect 27412 17444 27468 17454
rect 27412 17350 27468 17388
rect 27804 17444 27860 18396
rect 28140 18450 28196 18620
rect 28364 18676 28420 19740
rect 28364 18610 28420 18620
rect 28924 18676 28980 18686
rect 28140 18398 28142 18450
rect 28194 18398 28196 18450
rect 28140 18386 28196 18398
rect 28756 18452 28812 18462
rect 28756 18116 28812 18396
rect 28924 18450 28980 18620
rect 28924 18398 28926 18450
rect 28978 18398 28980 18450
rect 28924 18386 28980 18398
rect 28756 18050 28812 18060
rect 27804 17378 27860 17388
rect 28028 17220 28084 17230
rect 28028 16882 28084 17164
rect 28476 16996 28532 17006
rect 28364 16884 28420 16894
rect 28028 16830 28030 16882
rect 28082 16830 28084 16882
rect 25116 15262 25118 15314
rect 25170 15262 25172 15314
rect 25116 15250 25172 15262
rect 27468 16772 27524 16782
rect 25900 15202 25956 15214
rect 25900 15150 25902 15202
rect 25954 15150 25956 15202
rect 25004 15092 25284 15148
rect 24444 14466 24500 14476
rect 25228 14644 25284 15092
rect 25620 14644 25676 14654
rect 25228 14642 25676 14644
rect 25228 14590 25622 14642
rect 25674 14590 25676 14642
rect 25228 14588 25676 14590
rect 25228 14530 25284 14588
rect 25620 14578 25676 14588
rect 25900 14644 25956 15150
rect 25900 14578 25956 14588
rect 27020 14644 27076 14654
rect 27020 14550 27076 14588
rect 25228 14478 25230 14530
rect 25282 14478 25284 14530
rect 27468 14530 27524 16716
rect 27860 16212 27916 16222
rect 27860 16118 27916 16156
rect 27804 15428 27860 15438
rect 28028 15428 28084 16830
rect 28140 16828 28364 16884
rect 28140 16098 28196 16828
rect 28364 16790 28420 16828
rect 28476 16660 28532 16940
rect 28868 16882 28924 16894
rect 28868 16830 28870 16882
rect 28922 16830 28924 16882
rect 28868 16772 28924 16830
rect 28868 16706 28924 16716
rect 28140 16046 28142 16098
rect 28194 16046 28196 16098
rect 28140 16034 28196 16046
rect 28252 16604 28532 16660
rect 28252 16098 28308 16604
rect 28252 16046 28254 16098
rect 28306 16046 28308 16098
rect 28252 16034 28308 16046
rect 29036 16324 29092 19926
rect 29148 18564 29204 18574
rect 29148 18450 29204 18508
rect 29148 18398 29150 18450
rect 29202 18398 29204 18450
rect 29148 18386 29204 18398
rect 29260 18452 29316 18462
rect 29148 18228 29204 18238
rect 29148 16996 29204 18172
rect 29148 16882 29204 16940
rect 29148 16830 29150 16882
rect 29202 16830 29204 16882
rect 29148 16818 29204 16830
rect 29260 16884 29316 18396
rect 29428 18340 29484 18350
rect 29428 18246 29484 18284
rect 29596 17220 29652 20132
rect 31052 19796 31108 19806
rect 31052 19124 31108 19740
rect 31032 19068 31108 19124
rect 31032 18506 31088 19068
rect 30156 18452 30212 18490
rect 31032 18454 31034 18506
rect 31086 18454 31088 18506
rect 31032 18442 31088 18454
rect 31276 18450 31332 22204
rect 31388 21700 31444 28590
rect 34076 28644 34132 30830
rect 34412 29202 34468 29214
rect 34412 29150 34414 29202
rect 34466 29150 34468 29202
rect 34412 28866 34468 29150
rect 34412 28814 34414 28866
rect 34466 28814 34468 28866
rect 34412 28802 34468 28814
rect 34076 28642 34300 28644
rect 34076 28590 34078 28642
rect 34130 28590 34300 28642
rect 34076 28588 34300 28590
rect 34076 28578 34132 28588
rect 34244 28082 34300 28588
rect 34244 28030 34246 28082
rect 34298 28030 34300 28082
rect 34244 28018 34300 28030
rect 34300 26852 34356 26862
rect 33964 26292 34020 26302
rect 33964 26198 34020 26236
rect 34076 26180 34132 26190
rect 32060 25508 32116 25518
rect 31948 23156 32004 23166
rect 31948 22594 32004 23100
rect 31948 22542 31950 22594
rect 32002 22542 32004 22594
rect 31948 22530 32004 22542
rect 31388 21634 31444 21644
rect 32060 21028 32116 25452
rect 32396 25396 32452 25406
rect 32191 22314 32247 22326
rect 32191 22262 32193 22314
rect 32245 22262 32247 22314
rect 32191 22260 32247 22262
rect 32191 22194 32247 22204
rect 32060 20972 32228 21028
rect 32060 20804 32116 20814
rect 32060 20244 32116 20748
rect 32060 20018 32116 20188
rect 32172 20188 32228 20972
rect 32396 20188 32452 25340
rect 33068 22372 33124 22382
rect 33404 22372 33460 22382
rect 32956 22370 33460 22372
rect 32956 22318 33070 22370
rect 33122 22318 33406 22370
rect 33458 22318 33460 22370
rect 32956 22316 33460 22318
rect 32172 20132 32284 20188
rect 32396 20132 32564 20188
rect 32060 19966 32062 20018
rect 32114 19966 32116 20018
rect 32060 19954 32116 19966
rect 32228 19794 32284 20132
rect 32228 19742 32230 19794
rect 32282 19742 32284 19794
rect 32228 19684 32284 19742
rect 32228 19618 32284 19628
rect 30156 18386 30212 18396
rect 31276 18398 31278 18450
rect 31330 18398 31332 18450
rect 31276 18386 31332 18398
rect 29596 17154 29652 17164
rect 31836 17668 31892 17678
rect 30156 16996 30212 17006
rect 29260 16790 29316 16828
rect 30044 16884 30100 16894
rect 28532 15988 28588 15998
rect 27804 15426 28084 15428
rect 27804 15374 27806 15426
rect 27858 15374 28084 15426
rect 27804 15372 28084 15374
rect 28364 15986 28588 15988
rect 28364 15934 28534 15986
rect 28586 15934 28588 15986
rect 28364 15932 28588 15934
rect 27804 15362 27860 15372
rect 28364 15314 28420 15932
rect 28532 15922 28588 15932
rect 28364 15262 28366 15314
rect 28418 15262 28420 15314
rect 28364 15250 28420 15262
rect 28588 15316 28644 15326
rect 25228 14466 25284 14478
rect 27132 14486 27188 14498
rect 27132 14434 27134 14486
rect 27186 14434 27188 14486
rect 27468 14478 27470 14530
rect 27522 14478 27524 14530
rect 27468 14466 27524 14478
rect 28140 15204 28196 15214
rect 28140 14654 28196 15148
rect 28364 15146 28420 15158
rect 28364 15094 28366 15146
rect 28418 15094 28420 15146
rect 28140 14642 28252 14654
rect 28140 14590 28198 14642
rect 28250 14590 28252 14642
rect 28140 14578 28252 14590
rect 24892 14308 24948 14318
rect 24892 14214 24948 14252
rect 27132 13970 27188 14434
rect 27132 13918 27134 13970
rect 27186 13918 27188 13970
rect 27132 13906 27188 13918
rect 27244 14308 27300 14318
rect 13860 8818 13916 8830
rect 13860 8766 13862 8818
rect 13914 8766 13916 8818
rect 13860 8428 13916 8766
rect 14364 8428 14420 10108
rect 13580 8372 13748 8428
rect 13804 8372 13916 8428
rect 14140 8372 14420 8428
rect 16324 8372 16380 8382
rect 16828 8372 16884 12114
rect 18172 12066 18228 12078
rect 18172 12014 18174 12066
rect 18226 12014 18228 12066
rect 18172 11508 18228 12014
rect 20524 12010 20580 12022
rect 20524 11958 20526 12010
rect 20578 11958 20580 12010
rect 19852 11844 19908 11854
rect 18172 11442 18228 11452
rect 19740 11508 19796 11518
rect 19740 11414 19796 11452
rect 19852 11379 19908 11788
rect 20524 11844 20580 11958
rect 20524 11778 20580 11788
rect 20748 11508 20804 12348
rect 19852 11327 19854 11379
rect 19906 11327 19908 11379
rect 19852 11315 19908 11327
rect 20188 11452 20804 11508
rect 20972 12178 21028 12190
rect 20972 12126 20974 12178
rect 21026 12126 21028 12178
rect 20972 12068 21028 12126
rect 21532 12078 21588 13244
rect 21644 13244 21812 13300
rect 21644 12794 21700 13244
rect 21980 12964 22036 12974
rect 21980 12962 22148 12964
rect 21644 12742 21646 12794
rect 21698 12742 21700 12794
rect 21644 12730 21700 12742
rect 21756 12906 21812 12918
rect 21756 12854 21758 12906
rect 21810 12854 21812 12906
rect 21980 12910 21982 12962
rect 22034 12910 22148 12962
rect 21980 12908 22148 12910
rect 21980 12898 22036 12908
rect 21476 12068 21588 12078
rect 20972 12066 21588 12068
rect 20972 12014 21478 12066
rect 21530 12014 21588 12066
rect 20972 12012 21588 12014
rect 20188 11394 20244 11452
rect 20188 11342 20190 11394
rect 20242 11342 20244 11394
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 11342
rect 19964 9212 20244 9268
rect 20972 9268 21028 12012
rect 21476 12002 21532 12012
rect 21756 10724 21812 12854
rect 21756 10658 21812 10668
rect 21980 10612 22036 10622
rect 19964 9086 20020 9212
rect 13468 8260 13524 8270
rect 13468 8166 13524 8204
rect 13132 5842 13188 5852
rect 12796 5182 12798 5234
rect 12850 5182 12852 5234
rect 12796 5170 12852 5182
rect 13580 5246 13636 8372
rect 13804 8260 13860 8372
rect 13804 8194 13860 8204
rect 14140 8260 14196 8372
rect 16324 8370 16884 8372
rect 16324 8318 16326 8370
rect 16378 8318 16884 8370
rect 16324 8316 16884 8318
rect 19180 9044 19236 9054
rect 19180 8370 19236 8988
rect 19740 9044 19796 9054
rect 19740 8950 19796 8988
rect 19964 9034 19966 9086
rect 20018 9034 20020 9086
rect 19964 8484 20020 9034
rect 20188 9044 20244 9054
rect 19964 8418 20020 8428
rect 20076 8930 20132 8942
rect 20076 8878 20078 8930
rect 20130 8878 20132 8930
rect 19180 8318 19182 8370
rect 19234 8318 19236 8370
rect 16324 8306 16380 8316
rect 14756 8260 14812 8270
rect 14140 8258 14812 8260
rect 14140 8206 14142 8258
rect 14194 8206 14758 8258
rect 14810 8206 14812 8258
rect 14140 8204 14812 8206
rect 14140 8194 14196 8204
rect 14756 8194 14812 8204
rect 16492 8258 16548 8316
rect 16492 8206 16494 8258
rect 16546 8206 16548 8258
rect 16492 8194 16548 8206
rect 14252 8090 14308 8102
rect 14252 8038 14254 8090
rect 14306 8038 14308 8090
rect 14140 7588 14196 7598
rect 14140 7474 14196 7532
rect 14140 7422 14142 7474
rect 14194 7422 14196 7474
rect 14140 7410 14196 7422
rect 14252 7476 14308 8038
rect 14364 7476 14420 7486
rect 14252 7474 14420 7476
rect 14252 7422 14366 7474
rect 14418 7422 14420 7474
rect 14252 7420 14420 7422
rect 14364 7410 14420 7420
rect 14644 7250 14700 7262
rect 14644 7198 14646 7250
rect 14698 7198 14700 7250
rect 14140 6690 14196 6702
rect 14140 6638 14142 6690
rect 14194 6638 14196 6690
rect 14028 5908 14084 5918
rect 13804 5682 13860 5694
rect 13804 5630 13806 5682
rect 13858 5630 13860 5682
rect 13580 5236 13692 5246
rect 13636 5234 13692 5236
rect 13636 5182 13638 5234
rect 13690 5182 13692 5234
rect 13636 5180 13692 5182
rect 13580 5170 13692 5180
rect 13804 5236 13860 5630
rect 13804 5170 13860 5180
rect 14028 5234 14084 5852
rect 14140 5906 14196 6638
rect 14644 6690 14700 7198
rect 14644 6638 14646 6690
rect 14698 6638 14700 6690
rect 14644 6626 14700 6638
rect 14140 5854 14142 5906
rect 14194 5854 14196 5906
rect 14140 5842 14196 5854
rect 14028 5182 14030 5234
rect 14082 5182 14084 5234
rect 14028 5170 14084 5182
rect 15932 5236 15988 5246
rect 13580 5142 13636 5170
rect 15932 5142 15988 5180
rect 16716 5236 16772 8316
rect 19180 8306 19236 8318
rect 19740 8372 19796 8382
rect 17276 8260 17332 8270
rect 17276 8258 17556 8260
rect 17276 8206 17278 8258
rect 17330 8206 17556 8258
rect 17276 8204 17556 8206
rect 17276 8194 17332 8204
rect 17500 7812 17556 8204
rect 19740 8258 19796 8316
rect 19740 8206 19742 8258
rect 19794 8206 19796 8258
rect 19740 8194 19796 8206
rect 20076 8219 20132 8878
rect 20076 8167 20078 8219
rect 20130 8167 20132 8219
rect 20076 8155 20132 8167
rect 19740 8090 19796 8102
rect 18396 8036 18452 8046
rect 17500 7756 18116 7812
rect 18060 7698 18116 7756
rect 18060 7646 18062 7698
rect 18114 7646 18116 7698
rect 18060 7634 18116 7646
rect 18396 7474 18452 7980
rect 19740 8038 19742 8090
rect 19794 8038 19796 8090
rect 19740 8036 19796 8038
rect 19740 7970 19796 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 18396 7422 18398 7474
rect 18450 7422 18452 7474
rect 18396 7410 18452 7422
rect 20188 7474 20244 8988
rect 20804 8930 20860 8942
rect 20804 8878 20806 8930
rect 20858 8878 20860 8930
rect 20804 8596 20860 8878
rect 20804 8372 20860 8540
rect 20804 8306 20860 8316
rect 20300 8260 20356 8270
rect 20300 8258 20580 8260
rect 20300 8206 20302 8258
rect 20354 8206 20580 8258
rect 20300 8204 20580 8206
rect 20300 8194 20356 8204
rect 20188 7422 20190 7474
rect 20242 7422 20244 7474
rect 20188 7410 20244 7422
rect 20300 8036 20356 8046
rect 20300 7474 20356 7980
rect 20524 7598 20580 8204
rect 20524 7588 20636 7598
rect 20524 7586 20804 7588
rect 20524 7534 20582 7586
rect 20634 7534 20804 7586
rect 20524 7532 20804 7534
rect 20580 7522 20636 7532
rect 20300 7422 20302 7474
rect 20354 7422 20356 7474
rect 20300 7410 20356 7422
rect 20356 6468 20412 6478
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19740 6132 19796 6142
rect 19740 5906 19796 6076
rect 20356 6132 20412 6412
rect 20356 6066 20412 6076
rect 20748 6132 20804 7532
rect 20972 6468 21028 9212
rect 21868 10610 22036 10612
rect 21868 10558 21982 10610
rect 22034 10558 22036 10610
rect 21868 10556 22036 10558
rect 21868 9044 21924 10556
rect 21980 10546 22036 10556
rect 21868 8708 21924 8988
rect 21756 8652 21924 8708
rect 21644 8372 21700 8382
rect 21644 8278 21700 8316
rect 21308 8258 21364 8270
rect 21308 8206 21310 8258
rect 21362 8206 21364 8258
rect 21308 7476 21364 8206
rect 21756 8219 21812 8652
rect 21980 8260 22036 8270
rect 21756 8167 21758 8219
rect 21810 8167 21812 8219
rect 21756 8155 21812 8167
rect 21868 8258 22036 8260
rect 21868 8206 21982 8258
rect 22034 8206 22036 8258
rect 21868 8204 22036 8206
rect 21644 7476 21700 7486
rect 21308 7474 21700 7476
rect 21308 7422 21646 7474
rect 21698 7422 21700 7474
rect 21308 7420 21700 7422
rect 21644 6468 21700 7420
rect 21868 7474 21924 8204
rect 21980 8194 22036 8204
rect 22092 7598 22148 12908
rect 25754 10836 25810 10846
rect 24612 10778 24668 10790
rect 22484 10724 22540 10734
rect 22484 10630 22540 10668
rect 24612 10726 24614 10778
rect 24666 10726 24668 10778
rect 22204 10612 22260 10622
rect 22204 10518 22260 10556
rect 23772 10612 23828 10622
rect 23772 9938 23828 10556
rect 24444 10612 24500 10622
rect 24444 10518 24500 10556
rect 24612 10612 24668 10726
rect 25754 10648 25810 10780
rect 26516 10836 26572 10846
rect 26516 10742 26572 10780
rect 25754 10596 25756 10648
rect 25808 10596 25810 10648
rect 25754 10584 25810 10596
rect 25900 10610 25956 10622
rect 24612 10546 24668 10556
rect 25900 10558 25902 10610
rect 25954 10558 25956 10610
rect 25340 10388 25396 10398
rect 25340 10386 25508 10388
rect 25340 10334 25342 10386
rect 25394 10334 25508 10386
rect 25340 10332 25508 10334
rect 25340 10322 25396 10332
rect 23772 9886 23774 9938
rect 23826 9886 23828 9938
rect 23772 9874 23828 9886
rect 24444 9716 24500 9726
rect 24220 8372 24276 8382
rect 22316 8260 22372 8270
rect 22316 8166 22372 8204
rect 24220 8258 24276 8316
rect 24220 8206 24222 8258
rect 24274 8206 24276 8258
rect 24220 8194 24276 8206
rect 24444 8258 24500 9660
rect 25452 9156 25508 10332
rect 25676 9828 25732 9838
rect 25396 9100 25508 9156
rect 25564 9826 25732 9828
rect 25564 9774 25678 9826
rect 25730 9774 25732 9826
rect 25564 9772 25732 9774
rect 25564 9210 25620 9772
rect 25676 9762 25732 9772
rect 25900 9828 25956 10558
rect 26012 10612 26068 10622
rect 26012 10518 26068 10556
rect 26684 10612 26740 10622
rect 26572 9940 26628 9950
rect 25564 9158 25566 9210
rect 25618 9158 25620 9210
rect 25564 9146 25620 9158
rect 25396 9098 25452 9100
rect 25396 9046 25398 9098
rect 25450 9046 25452 9098
rect 25396 9034 25452 9046
rect 25676 9044 25732 9054
rect 25676 8950 25732 8988
rect 25900 8484 25956 9772
rect 26460 9828 26516 9838
rect 26572 9828 26628 9884
rect 26460 9826 26628 9828
rect 26460 9774 26462 9826
rect 26514 9774 26628 9826
rect 26460 9772 26628 9774
rect 26460 9762 26516 9772
rect 25900 8418 25956 8428
rect 26572 8942 26628 9772
rect 26684 9826 26740 10556
rect 27132 9938 27188 9950
rect 27132 9886 27134 9938
rect 27186 9886 27188 9938
rect 26684 9774 26686 9826
rect 26738 9774 26740 9826
rect 26684 9762 26740 9774
rect 27020 9828 27076 9838
rect 27020 9759 27022 9772
rect 27074 9759 27076 9772
rect 27020 9734 27076 9759
rect 27132 9044 27188 9886
rect 26572 8930 26684 8942
rect 26572 8878 26630 8930
rect 26682 8878 26684 8930
rect 26572 8866 26684 8878
rect 24444 8206 24446 8258
rect 24498 8206 24500 8258
rect 24444 8194 24500 8206
rect 23940 8148 23996 8158
rect 23772 8146 23996 8148
rect 23772 8094 23942 8146
rect 23994 8094 23996 8146
rect 23772 8092 23996 8094
rect 22092 7586 22204 7598
rect 22092 7534 22150 7586
rect 22202 7534 22204 7586
rect 22092 7532 22204 7534
rect 22148 7522 22204 7532
rect 21868 7422 21870 7474
rect 21922 7422 21924 7474
rect 21868 6914 21924 7422
rect 21868 6862 21870 6914
rect 21922 6862 21924 6914
rect 21868 6850 21924 6862
rect 22428 6914 22484 6926
rect 22428 6862 22430 6914
rect 22482 6862 22484 6914
rect 20972 6402 21028 6412
rect 21420 6412 21700 6468
rect 20748 6076 21364 6132
rect 19740 5854 19742 5906
rect 19794 5854 19796 5906
rect 19740 5842 19796 5854
rect 19964 5908 20020 5918
rect 19964 5814 20020 5852
rect 20468 5908 20524 5918
rect 20468 5814 20524 5852
rect 20748 5906 20804 6076
rect 20748 5854 20750 5906
rect 20802 5854 20804 5906
rect 20748 5842 20804 5854
rect 20860 5908 20916 5918
rect 21084 5908 21140 5918
rect 20860 5906 21140 5908
rect 20860 5854 20862 5906
rect 20914 5854 21086 5906
rect 21138 5854 21140 5906
rect 20860 5852 21140 5854
rect 20076 5738 20132 5750
rect 20076 5686 20078 5738
rect 20130 5686 20132 5738
rect 10108 5070 10110 5122
rect 10162 5070 10164 5122
rect 10108 5058 10164 5070
rect 16716 5124 16772 5180
rect 17444 5236 17500 5246
rect 17500 5180 17668 5236
rect 17444 5142 17500 5180
rect 16716 5122 16940 5124
rect 16716 5070 16718 5122
rect 16770 5070 16940 5122
rect 16716 5068 16940 5070
rect 16716 5058 16772 5068
rect 7532 4510 7534 4562
rect 7586 4510 7588 4562
rect 7532 4498 7588 4510
rect 8204 4844 8484 4900
rect 7868 4340 7924 4350
rect 8204 4340 8260 4844
rect 16884 4562 16940 5068
rect 17612 5122 17668 5180
rect 17612 5070 17614 5122
rect 17666 5070 17668 5122
rect 17612 5058 17668 5070
rect 18396 5122 18452 5134
rect 18396 5070 18398 5122
rect 18450 5070 18452 5122
rect 16884 4510 16886 4562
rect 16938 4510 16940 4562
rect 16884 4498 16940 4510
rect 7868 4338 8260 4340
rect 7868 4286 7870 4338
rect 7922 4286 8260 4338
rect 7868 4284 8260 4286
rect 7868 4274 7924 4284
rect 18396 4228 18452 5070
rect 20076 4900 20132 5686
rect 20412 5684 20468 5694
rect 20300 5236 20356 5246
rect 20300 5142 20356 5180
rect 20076 4844 20244 4900
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20188 4564 20244 4844
rect 20076 4508 20244 4564
rect 20076 4382 20132 4508
rect 20076 4330 20078 4382
rect 20130 4330 20132 4382
rect 20076 4318 20132 4330
rect 20412 4338 20468 5628
rect 20860 5236 20916 5852
rect 21084 5684 21140 5852
rect 21308 5906 21364 6076
rect 21308 5854 21310 5906
rect 21362 5854 21364 5906
rect 21308 5842 21364 5854
rect 21420 5684 21476 6412
rect 22428 5906 22484 6862
rect 22428 5854 22430 5906
rect 22482 5854 22484 5906
rect 21084 5628 21476 5684
rect 21588 5684 21644 5694
rect 21588 5590 21644 5628
rect 22428 5236 22484 5854
rect 22540 5906 22596 5918
rect 22540 5854 22542 5906
rect 22594 5854 22596 5906
rect 22540 5684 22596 5854
rect 22820 5908 22876 5918
rect 22820 5814 22876 5852
rect 23548 5908 23604 5918
rect 23548 5814 23604 5852
rect 23772 5906 23828 8092
rect 23940 8082 23996 8092
rect 23772 5854 23774 5906
rect 23826 5854 23828 5906
rect 23772 5842 23828 5854
rect 24052 5684 24108 5694
rect 22540 5618 22596 5628
rect 23884 5682 24108 5684
rect 23884 5630 24054 5682
rect 24106 5630 24108 5682
rect 23884 5628 24108 5630
rect 23212 5236 23268 5246
rect 22428 5234 23268 5236
rect 22428 5182 23214 5234
rect 23266 5182 23268 5234
rect 22428 5180 23268 5182
rect 20860 5170 20916 5180
rect 23212 5170 23268 5180
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 23884 4338 23940 5628
rect 24052 5618 24108 5628
rect 25116 5124 25172 5134
rect 24892 5122 25172 5124
rect 24892 5070 25118 5122
rect 25170 5070 25172 5122
rect 24892 5068 25172 5070
rect 24892 4676 24948 5068
rect 25116 5058 25172 5068
rect 25900 5124 25956 5134
rect 26292 5124 26348 5134
rect 26572 5124 26628 8866
rect 27132 6356 27188 8988
rect 27132 6290 27188 6300
rect 27244 8596 27300 14252
rect 27468 13522 27524 13534
rect 27468 13470 27470 13522
rect 27522 13470 27524 13522
rect 27468 10610 27524 13470
rect 28140 13522 28196 14578
rect 28364 13970 28420 15094
rect 28364 13918 28366 13970
rect 28418 13918 28420 13970
rect 28364 13906 28420 13918
rect 28140 13470 28142 13522
rect 28194 13470 28196 13522
rect 28140 13458 28196 13470
rect 27916 11396 27972 11406
rect 27916 11394 28084 11396
rect 27916 11342 27918 11394
rect 27970 11342 28084 11394
rect 27916 11340 28084 11342
rect 27916 11330 27972 11340
rect 27468 10558 27470 10610
rect 27522 10558 27524 10610
rect 27468 9940 27524 10558
rect 27468 9874 27524 9884
rect 27804 10388 27860 10398
rect 27580 9826 27636 9838
rect 27580 9774 27582 9826
rect 27634 9774 27636 9826
rect 27412 9268 27468 9278
rect 27580 9268 27636 9774
rect 27804 9826 27860 10332
rect 28028 10062 28084 11340
rect 28252 11170 28308 11182
rect 28252 11118 28254 11170
rect 28306 11118 28308 11170
rect 28252 10610 28308 11118
rect 28588 10836 28644 15260
rect 29036 15314 29092 16268
rect 29148 16212 29204 16222
rect 29148 16070 29204 16156
rect 29148 16018 29150 16070
rect 29202 16018 29204 16070
rect 29148 15876 29204 16018
rect 29148 15810 29204 15820
rect 29036 15262 29038 15314
rect 29090 15262 29092 15314
rect 29036 15204 29092 15262
rect 29708 15540 29764 15550
rect 29708 15314 29764 15484
rect 29708 15262 29710 15314
rect 29762 15262 29764 15314
rect 29036 15138 29092 15148
rect 29540 15204 29596 15214
rect 29540 14642 29596 15148
rect 29540 14590 29542 14642
rect 29594 14590 29596 14642
rect 29540 14578 29596 14590
rect 28252 10558 28254 10610
rect 28306 10558 28308 10610
rect 28252 10546 28308 10558
rect 28476 10780 28644 10836
rect 29708 10836 29764 15262
rect 29876 15428 29932 15438
rect 29876 15370 29932 15372
rect 29876 15318 29878 15370
rect 29930 15318 29932 15370
rect 30044 15426 30100 16828
rect 30156 16548 30212 16940
rect 31164 16772 31220 16782
rect 30940 16660 30996 16670
rect 30156 16492 30324 16548
rect 30156 16324 30212 16334
rect 30156 16230 30212 16268
rect 30268 16100 30324 16492
rect 30044 15374 30046 15426
rect 30098 15374 30100 15426
rect 30044 15362 30100 15374
rect 30156 16044 30324 16100
rect 29876 14756 29932 15318
rect 30156 15314 30212 16044
rect 30940 15428 30996 16604
rect 30156 15262 30158 15314
rect 30210 15262 30212 15314
rect 30156 15250 30212 15262
rect 30436 15316 30492 15326
rect 30436 15222 30492 15260
rect 30940 15314 30996 15372
rect 30940 15262 30942 15314
rect 30994 15262 30996 15314
rect 31164 15358 31220 16716
rect 31164 15306 31166 15358
rect 31218 15306 31220 15358
rect 31164 15294 31220 15306
rect 31612 15314 31668 15326
rect 30940 15250 30996 15262
rect 31612 15262 31614 15314
rect 31666 15262 31668 15314
rect 31276 15204 31332 15214
rect 31612 15204 31668 15262
rect 31276 15202 31668 15204
rect 31276 15150 31278 15202
rect 31330 15150 31668 15202
rect 31276 15148 31668 15150
rect 31276 15138 31332 15148
rect 29876 14700 30100 14756
rect 30044 14642 30100 14700
rect 30044 14590 30046 14642
rect 30098 14590 30100 14642
rect 30044 14578 30100 14590
rect 28476 10276 28532 10780
rect 29708 10770 29764 10780
rect 30604 10612 30660 10622
rect 30380 10610 30660 10612
rect 30380 10558 30606 10610
rect 30658 10558 30660 10610
rect 30380 10556 30660 10558
rect 30156 10500 30212 10510
rect 30380 10500 30436 10556
rect 30604 10546 30660 10556
rect 31480 10612 31536 10622
rect 31480 10518 31536 10556
rect 30156 10498 30436 10500
rect 30156 10446 30158 10498
rect 30210 10446 30436 10498
rect 30156 10444 30436 10446
rect 28476 10220 28644 10276
rect 28028 10050 28140 10062
rect 28028 9998 28086 10050
rect 28138 9998 28140 10050
rect 28028 9996 28140 9998
rect 28084 9986 28140 9996
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9762 27860 9774
rect 28588 9716 28644 10220
rect 30156 10164 30212 10444
rect 31724 10388 31780 10398
rect 31724 10294 31780 10332
rect 30156 10098 30212 10108
rect 30940 10164 30996 10174
rect 31836 10164 31892 17612
rect 32508 15550 32564 20132
rect 32956 16660 33012 22316
rect 33068 22306 33124 22316
rect 33404 22306 33460 22316
rect 34076 21812 34132 26124
rect 34300 26066 34356 26796
rect 34300 26014 34302 26066
rect 34354 26014 34356 26066
rect 34300 25396 34356 26014
rect 34300 25330 34356 25340
rect 34636 26292 34692 31948
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34972 30212 35028 30222
rect 34806 28644 34862 28654
rect 34806 28550 34862 28588
rect 34972 28642 35028 30156
rect 35644 30212 35700 34106
rect 35756 31948 35812 35308
rect 36428 34914 36484 35644
rect 36428 34862 36430 34914
rect 36482 34862 36484 34914
rect 36428 34850 36484 34862
rect 36260 34690 36316 34702
rect 36260 34638 36262 34690
rect 36314 34638 36316 34690
rect 36260 34580 36316 34638
rect 35868 34524 36316 34580
rect 35868 34130 35924 34524
rect 36092 34244 36148 34254
rect 36092 34150 36148 34188
rect 35868 34078 35870 34130
rect 35922 34078 35924 34130
rect 35868 34066 35924 34078
rect 36260 34074 36316 34086
rect 36260 34022 36262 34074
rect 36314 34022 36316 34074
rect 36260 33460 36316 34022
rect 36260 33404 36372 33460
rect 36316 32686 36372 33404
rect 36316 32674 36428 32686
rect 36316 32622 36374 32674
rect 36426 32622 36428 32674
rect 36316 32620 36428 32622
rect 36372 32610 36428 32620
rect 35756 31892 36148 31948
rect 35980 31108 36036 31118
rect 35980 31014 36036 31052
rect 35812 30938 35868 30950
rect 35812 30886 35814 30938
rect 35866 30886 35868 30938
rect 35812 30436 35868 30886
rect 35812 30380 36036 30436
rect 35644 30146 35700 30156
rect 35532 30100 35588 30110
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34972 28590 34974 28642
rect 35026 28590 35028 28642
rect 34972 28578 35028 28590
rect 35084 28868 35140 28878
rect 35532 28868 35588 30044
rect 35084 28642 35140 28812
rect 35420 28812 35588 28868
rect 35420 28644 35476 28812
rect 35084 28590 35086 28642
rect 35138 28590 35140 28642
rect 35084 28578 35140 28590
rect 35196 28642 35476 28644
rect 35196 28590 35422 28642
rect 35474 28590 35476 28642
rect 35868 28756 35924 28766
rect 35868 28642 35924 28700
rect 35196 28588 35476 28590
rect 35196 28094 35252 28588
rect 35420 28578 35476 28588
rect 35588 28586 35644 28598
rect 35140 28082 35252 28094
rect 35140 28030 35142 28082
rect 35194 28030 35252 28082
rect 35140 28028 35252 28030
rect 35588 28534 35590 28586
rect 35642 28534 35644 28586
rect 35868 28590 35870 28642
rect 35922 28590 35924 28642
rect 35868 28578 35924 28590
rect 35588 28084 35644 28534
rect 35756 28530 35812 28542
rect 35756 28478 35758 28530
rect 35810 28478 35812 28530
rect 35756 28420 35812 28478
rect 35756 28364 35924 28420
rect 35588 28028 35812 28084
rect 35140 28018 35196 28028
rect 35644 27748 35700 27758
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35532 27300 35588 27310
rect 35196 27074 35252 27086
rect 35196 27022 35198 27074
rect 35250 27022 35252 27074
rect 35532 27074 35588 27244
rect 34916 26852 34972 26862
rect 34916 26758 34972 26796
rect 35196 26852 35252 27022
rect 35196 26786 35252 26796
rect 35364 27018 35420 27030
rect 35364 26966 35366 27018
rect 35418 26966 35420 27018
rect 35532 27022 35534 27074
rect 35586 27022 35588 27074
rect 35532 27010 35588 27022
rect 35644 27074 35700 27692
rect 35644 27022 35646 27074
rect 35698 27022 35700 27074
rect 35644 27010 35700 27022
rect 35364 26404 35420 26966
rect 35364 26348 35588 26404
rect 34636 24724 34692 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25508 35588 26348
rect 35532 25442 35588 25452
rect 34748 24724 34804 24734
rect 34636 24722 34804 24724
rect 34636 24670 34750 24722
rect 34802 24670 34804 24722
rect 34636 24668 34804 24670
rect 35756 24724 35812 28028
rect 35868 27524 35924 28364
rect 35868 27458 35924 27468
rect 35980 27310 36036 30380
rect 36092 28756 36148 31892
rect 36316 31780 36372 31790
rect 36316 31686 36372 31724
rect 36204 31556 36260 31566
rect 36204 30994 36260 31500
rect 36204 30942 36206 30994
rect 36258 30942 36260 30994
rect 36204 30930 36260 30942
rect 36428 31022 36484 31034
rect 36428 30970 36430 31022
rect 36482 30970 36484 31022
rect 36428 30212 36484 30970
rect 36428 30146 36484 30156
rect 36540 29204 36596 35980
rect 37100 35812 37156 35822
rect 36652 35700 36708 35710
rect 37100 35700 37156 35756
rect 38892 35812 38948 35822
rect 36652 35606 36708 35644
rect 36876 35698 37156 35700
rect 36876 35646 37102 35698
rect 37154 35646 37156 35698
rect 36876 35644 37156 35646
rect 36876 35364 36932 35644
rect 37100 35634 37156 35644
rect 37976 35700 38032 35710
rect 37976 35606 38032 35644
rect 38892 35700 38948 35756
rect 39116 35700 39172 35710
rect 38892 35698 39172 35700
rect 38892 35646 39118 35698
rect 39170 35646 39172 35698
rect 38892 35644 39172 35646
rect 38892 35598 38948 35644
rect 39116 35634 39172 35644
rect 39228 35700 39284 38612
rect 39676 38050 39732 38612
rect 40460 38052 40516 38062
rect 39676 37998 39678 38050
rect 39730 37998 39732 38050
rect 39508 37828 39564 37838
rect 39676 37828 39732 37998
rect 39508 37826 39732 37828
rect 39508 37774 39510 37826
rect 39562 37774 39732 37826
rect 39508 37772 39732 37774
rect 39508 37762 39564 37772
rect 39676 36260 39732 37772
rect 40124 38050 40516 38052
rect 40124 37998 40462 38050
rect 40514 37998 40516 38050
rect 40124 37996 40516 37998
rect 40124 36594 40180 37996
rect 40460 37986 40516 37996
rect 40124 36542 40126 36594
rect 40178 36542 40180 36594
rect 40124 36530 40180 36542
rect 39676 36194 39732 36204
rect 39956 36426 40012 36438
rect 39956 36374 39958 36426
rect 40010 36374 40012 36426
rect 40572 36426 40628 36438
rect 39956 35924 40012 36374
rect 39228 35634 39284 35644
rect 39788 35868 40012 35924
rect 40124 36372 40180 36382
rect 38836 35586 38948 35598
rect 38836 35534 38838 35586
rect 38890 35534 38948 35586
rect 38836 35532 38948 35534
rect 38220 35474 38276 35486
rect 38220 35422 38222 35474
rect 38274 35422 38276 35474
rect 36876 35308 37156 35364
rect 37100 35038 37156 35308
rect 37100 35026 37212 35038
rect 37100 34974 37158 35026
rect 37210 34974 37212 35026
rect 37100 34972 37212 34974
rect 37156 34962 37212 34972
rect 38220 34916 38276 35422
rect 38836 35364 38892 35532
rect 38836 35308 39060 35364
rect 38220 34850 38276 34860
rect 38444 34914 38500 34926
rect 38444 34862 38446 34914
rect 38498 34862 38500 34914
rect 38892 34916 38948 34926
rect 36764 32676 36820 32686
rect 36764 32582 36820 32620
rect 36652 32562 36708 32574
rect 36652 32510 36654 32562
rect 36706 32510 36708 32562
rect 37100 32564 37156 32574
rect 36652 32452 36708 32510
rect 36652 32386 36708 32396
rect 36932 32506 36988 32518
rect 36932 32454 36934 32506
rect 36986 32454 36988 32506
rect 37100 32470 37156 32508
rect 37324 32562 37380 32574
rect 37324 32510 37326 32562
rect 37378 32510 37380 32562
rect 36932 31948 36988 32454
rect 37324 32004 37380 32510
rect 37660 32564 37716 32574
rect 37660 32470 37716 32508
rect 38444 32564 38500 34862
rect 38612 34858 38668 34870
rect 38612 34806 38614 34858
rect 38666 34806 38668 34858
rect 38892 34822 38948 34860
rect 38612 34692 38668 34806
rect 38612 34626 38668 34636
rect 38780 34804 38836 34814
rect 38444 32498 38500 32508
rect 36932 31892 37044 31948
rect 37324 31938 37380 31948
rect 36876 31780 36932 31790
rect 36876 31686 36932 31724
rect 36988 31566 37044 31892
rect 36988 31556 37100 31566
rect 36988 31500 37044 31556
rect 37044 31462 37100 31500
rect 36540 29138 36596 29148
rect 36092 28700 36372 28756
rect 36148 28532 36204 28542
rect 36148 28438 36204 28476
rect 35924 27298 36036 27310
rect 35924 27246 35926 27298
rect 35978 27246 36036 27298
rect 35924 27244 36036 27246
rect 35924 27234 35980 27244
rect 35756 24668 36036 24724
rect 34748 24658 34804 24668
rect 34412 24500 34468 24510
rect 34412 24406 34468 24444
rect 35644 24500 35700 24510
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35476 23714 35532 23726
rect 35476 23662 35478 23714
rect 35530 23662 35532 23714
rect 35476 23492 35532 23662
rect 35476 23426 35532 23436
rect 35644 23156 35700 24444
rect 35812 24498 35868 24510
rect 35812 24446 35814 24498
rect 35866 24446 35868 24498
rect 35812 24162 35868 24446
rect 35812 24110 35814 24162
rect 35866 24110 35868 24162
rect 35812 24098 35868 24110
rect 35532 23100 35700 23156
rect 34860 22932 34916 22942
rect 34524 22484 34580 22494
rect 34524 22390 34580 22428
rect 34280 22372 34336 22382
rect 34280 22278 34336 22316
rect 34860 22370 34916 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34860 22318 34862 22370
rect 34914 22318 34916 22370
rect 34860 22260 34916 22318
rect 34188 21812 34244 21822
rect 34076 21810 34244 21812
rect 34076 21758 34190 21810
rect 34242 21758 34244 21810
rect 34076 21756 34244 21758
rect 34188 21746 34244 21756
rect 33292 21700 33348 21710
rect 33124 20186 33180 20198
rect 33124 20134 33126 20186
rect 33178 20134 33180 20186
rect 33124 20132 33180 20134
rect 33124 19796 33180 20076
rect 33292 20018 33348 21644
rect 34860 21698 34916 22204
rect 35028 22372 35084 22382
rect 35028 22202 35084 22316
rect 35028 22150 35030 22202
rect 35082 22150 35084 22202
rect 35028 22138 35084 22150
rect 34860 21646 34862 21698
rect 34914 21646 34916 21698
rect 34860 21634 34916 21646
rect 33292 19966 33294 20018
rect 33346 19966 33348 20018
rect 33292 19954 33348 19966
rect 33404 21588 33460 21598
rect 33404 20244 33460 21532
rect 34524 21588 34580 21598
rect 34524 21494 34580 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35532 21028 35588 23100
rect 35980 22932 36036 24668
rect 36316 24498 36372 28700
rect 37100 28644 37156 28654
rect 37100 28082 37156 28588
rect 38780 28644 38836 34748
rect 39004 30100 39060 35308
rect 39788 35252 39844 35868
rect 40124 35812 40180 36316
rect 39992 35756 40180 35812
rect 40572 36374 40574 36426
rect 40626 36374 40628 36426
rect 39992 35754 40048 35756
rect 39992 35702 39994 35754
rect 40046 35702 40048 35754
rect 39992 35690 40048 35702
rect 39172 35196 39844 35252
rect 40236 35474 40292 35486
rect 40236 35422 40238 35474
rect 40290 35422 40292 35474
rect 39172 35138 39228 35196
rect 39172 35086 39174 35138
rect 39226 35086 39228 35138
rect 39172 35074 39228 35086
rect 39340 35028 39396 35038
rect 39340 31556 39396 34972
rect 39676 34914 39732 34926
rect 39676 34862 39678 34914
rect 39730 34862 39732 34914
rect 40124 34916 40180 34926
rect 40236 34916 40292 35422
rect 40572 35028 40628 36374
rect 40572 34962 40628 34972
rect 40124 34914 40292 34916
rect 39676 32564 39732 34862
rect 39844 34858 39900 34870
rect 39844 34806 39846 34858
rect 39898 34806 39900 34858
rect 40124 34862 40126 34914
rect 40178 34862 40292 34914
rect 40124 34860 40292 34862
rect 40404 34916 40460 34926
rect 40124 34850 40180 34860
rect 40404 34822 40460 34860
rect 39844 34804 39900 34806
rect 39676 32498 39732 32508
rect 39788 34748 39900 34804
rect 40012 34804 40068 34814
rect 39788 34692 39844 34748
rect 40012 34710 40068 34748
rect 39004 30034 39060 30044
rect 39228 31554 39396 31556
rect 39228 31502 39342 31554
rect 39394 31502 39396 31554
rect 39228 31500 39396 31502
rect 39228 30210 39284 31500
rect 39340 31490 39396 31500
rect 39228 30158 39230 30210
rect 39282 30158 39284 30210
rect 39228 28866 39284 30158
rect 39228 28814 39230 28866
rect 39282 28814 39284 28866
rect 39228 28802 39284 28814
rect 39340 30212 39396 30222
rect 39788 30212 39844 34636
rect 40292 31554 40348 31566
rect 40292 31502 40294 31554
rect 40346 31502 40348 31554
rect 40292 31218 40348 31502
rect 40292 31166 40294 31218
rect 40346 31166 40348 31218
rect 40292 31154 40348 31166
rect 40684 30660 40740 39566
rect 42924 39620 42980 39630
rect 42924 39526 42980 39564
rect 43316 39620 43372 39630
rect 43484 39620 43540 40238
rect 43372 39564 43540 39620
rect 43316 39526 43372 39564
rect 42364 37938 42420 37950
rect 42364 37886 42366 37938
rect 42418 37886 42420 37938
rect 41132 37266 41188 37278
rect 41132 37214 41134 37266
rect 41186 37214 41188 37266
rect 40964 37044 41020 37054
rect 40796 37042 41020 37044
rect 40796 36990 40966 37042
rect 41018 36990 41020 37042
rect 40796 36988 41020 36990
rect 40796 36538 40852 36988
rect 40964 36978 41020 36988
rect 40796 36486 40798 36538
rect 40850 36486 40852 36538
rect 40796 36474 40852 36486
rect 41132 36932 41188 37214
rect 41132 36372 41188 36876
rect 42364 36932 42420 37886
rect 42364 36866 42420 36876
rect 41132 36306 41188 36316
rect 41300 36260 41356 36270
rect 41132 35700 41188 35710
rect 41300 35700 41356 36204
rect 41132 35698 41356 35700
rect 41132 35646 41134 35698
rect 41186 35646 41356 35698
rect 41132 35644 41356 35646
rect 41132 35140 41188 35644
rect 41916 35588 41972 35598
rect 40796 35084 41188 35140
rect 41244 35586 41972 35588
rect 41244 35534 41918 35586
rect 41970 35534 41972 35586
rect 41244 35532 41972 35534
rect 40796 31556 40852 35084
rect 40964 34916 41020 34926
rect 40964 34822 41020 34860
rect 41132 34916 41188 34926
rect 41244 34916 41300 35532
rect 41916 35522 41972 35532
rect 43820 35586 43876 35598
rect 43820 35534 43822 35586
rect 43874 35534 43876 35586
rect 42812 35364 42868 35374
rect 41580 35028 41636 35038
rect 41132 34914 41300 34916
rect 41132 34862 41134 34914
rect 41186 34862 41300 34914
rect 41132 34860 41300 34862
rect 41356 34914 41412 34926
rect 41356 34862 41358 34914
rect 41410 34862 41412 34914
rect 41132 34850 41188 34860
rect 41356 34692 41412 34862
rect 41356 33236 41412 34636
rect 41076 33180 41412 33236
rect 41580 34886 41636 34972
rect 41580 34834 41582 34886
rect 41634 34834 41636 34886
rect 42812 34914 42868 35308
rect 43820 35364 43876 35534
rect 43820 35298 43876 35308
rect 42812 34862 42814 34914
rect 42866 34862 42868 34914
rect 42812 34850 42868 34862
rect 41076 32618 41132 33180
rect 40908 32564 40964 32574
rect 41076 32566 41078 32618
rect 41130 32566 41132 32618
rect 41076 32554 41132 32566
rect 41244 32676 41300 32686
rect 40908 32470 40964 32508
rect 40964 31556 41020 31566
rect 41244 31556 41300 32620
rect 40796 31554 41076 31556
rect 40796 31502 40966 31554
rect 41018 31502 41076 31554
rect 40796 31500 41076 31502
rect 40964 31490 41076 31500
rect 41244 31490 41300 31500
rect 41356 32562 41412 32574
rect 41580 32564 41636 34834
rect 42644 34692 42700 34702
rect 42644 34598 42700 34636
rect 41356 32510 41358 32562
rect 41410 32510 41412 32562
rect 41356 32452 41412 32510
rect 40348 30604 40740 30660
rect 41020 30996 41076 31490
rect 41132 30996 41188 31006
rect 41020 30994 41188 30996
rect 41020 30942 41134 30994
rect 41186 30942 41188 30994
rect 41020 30940 41188 30942
rect 40348 30548 40404 30604
rect 40012 30492 40404 30548
rect 39900 30436 39956 30446
rect 40012 30436 40068 30492
rect 39900 30434 40068 30436
rect 39900 30382 39902 30434
rect 39954 30382 40068 30434
rect 39900 30380 40068 30382
rect 39900 30370 39956 30380
rect 40348 30212 40404 30222
rect 38780 28578 38836 28588
rect 39004 28644 39060 28654
rect 37100 28030 37102 28082
rect 37154 28030 37156 28082
rect 37100 28018 37156 28030
rect 37940 27972 37996 27982
rect 37996 27916 38164 27972
rect 37940 27878 37996 27916
rect 36764 27858 36820 27870
rect 36764 27806 36766 27858
rect 36818 27806 36820 27858
rect 36596 27748 36652 27758
rect 36764 27748 36820 27806
rect 38108 27858 38164 27916
rect 38108 27806 38110 27858
rect 38162 27806 38164 27858
rect 38108 27794 38164 27806
rect 38444 27860 38500 27870
rect 38444 27766 38500 27804
rect 36540 27746 36820 27748
rect 36540 27694 36598 27746
rect 36650 27694 36820 27746
rect 36540 27692 36820 27694
rect 37884 27748 37940 27758
rect 36540 27682 36652 27692
rect 36540 26974 36596 27682
rect 36484 26964 36596 26974
rect 36540 26908 36596 26964
rect 36652 27524 36708 27534
rect 36652 27076 36708 27468
rect 37212 27300 37268 27310
rect 37212 27206 37268 27244
rect 37884 27298 37940 27692
rect 39004 27636 39060 28588
rect 39116 28084 39172 28094
rect 39340 28084 39396 30156
rect 39508 30154 39564 30166
rect 39788 30156 39956 30212
rect 39508 30102 39510 30154
rect 39562 30102 39564 30154
rect 39508 29540 39564 30102
rect 39508 29484 39844 29540
rect 39676 28866 39732 28878
rect 39676 28814 39678 28866
rect 39730 28814 39732 28866
rect 39116 28082 39396 28084
rect 39116 28030 39118 28082
rect 39170 28030 39396 28082
rect 39116 28028 39396 28030
rect 39452 28418 39508 28430
rect 39452 28366 39454 28418
rect 39506 28366 39508 28418
rect 39116 28018 39172 28028
rect 39452 27858 39508 28366
rect 39452 27806 39454 27858
rect 39506 27806 39508 27858
rect 39452 27794 39508 27806
rect 39004 27580 39620 27636
rect 39452 27412 39508 27422
rect 37884 27246 37886 27298
rect 37938 27246 37940 27298
rect 37884 27234 37940 27246
rect 38780 27244 39340 27300
rect 36484 26870 36540 26908
rect 36540 26516 36596 26526
rect 36652 26516 36708 27020
rect 36540 26514 36708 26516
rect 36540 26462 36542 26514
rect 36594 26462 36708 26514
rect 36540 26460 36708 26462
rect 36876 27074 36932 27086
rect 36876 27022 36878 27074
rect 36930 27022 36932 27074
rect 36540 26450 36596 26460
rect 36876 26292 36932 27022
rect 37548 27074 37604 27086
rect 37548 27022 37550 27074
rect 37602 27022 37604 27074
rect 37324 26964 37380 26974
rect 37548 26964 37604 27022
rect 37380 26908 37604 26964
rect 37100 26292 37156 26302
rect 36876 26290 37044 26292
rect 36876 26238 36878 26290
rect 36930 26238 37044 26290
rect 36876 26236 37044 26238
rect 36876 26226 36932 26236
rect 36316 24446 36318 24498
rect 36370 24446 36372 24498
rect 36316 24434 36372 24446
rect 35980 22866 36036 22876
rect 36092 23938 36148 23950
rect 36092 23886 36094 23938
rect 36146 23886 36148 23938
rect 36092 23492 36148 23886
rect 36316 23940 36372 23950
rect 36316 23846 36372 23884
rect 36988 23938 37044 26236
rect 37100 26198 37156 26236
rect 36988 23886 36990 23938
rect 37042 23886 37044 23938
rect 36092 22596 36148 23436
rect 36708 23044 36764 23054
rect 36708 22950 36764 22988
rect 36092 22530 36148 22540
rect 35980 22372 36036 22382
rect 35420 20972 35588 21028
rect 35644 22314 35700 22326
rect 35644 22262 35646 22314
rect 35698 22262 35700 22314
rect 35980 22278 36036 22316
rect 36372 22372 36428 22382
rect 36372 22278 36428 22316
rect 35420 20188 35476 20972
rect 35644 20916 35700 22262
rect 36204 22258 36260 22270
rect 36204 22206 36206 22258
rect 36258 22206 36260 22258
rect 36204 21924 36260 22206
rect 36204 21868 36820 21924
rect 36764 21586 36820 21868
rect 36764 21534 36766 21586
rect 36818 21534 36820 21586
rect 36764 21522 36820 21534
rect 33124 19730 33180 19740
rect 33404 18562 33460 20188
rect 35364 20132 35476 20188
rect 35532 20860 35700 20916
rect 35364 20130 35420 20132
rect 35364 20078 35366 20130
rect 35418 20078 35420 20130
rect 35364 20020 35420 20078
rect 35364 19954 35420 19964
rect 34972 19684 35028 19694
rect 34972 19290 35028 19628
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34972 19238 34974 19290
rect 35026 19238 35028 19290
rect 34972 19226 35028 19238
rect 35532 19460 35588 20860
rect 36092 20356 36148 20366
rect 35980 20244 36036 20254
rect 35812 20132 35868 20142
rect 35812 20074 35868 20076
rect 35644 20020 35700 20030
rect 35812 20022 35814 20074
rect 35866 20022 35868 20074
rect 35980 20130 36036 20188
rect 35980 20078 35982 20130
rect 36034 20078 36036 20130
rect 35980 20066 36036 20078
rect 35812 20010 35868 20022
rect 36092 20018 36148 20300
rect 35644 19926 35700 19964
rect 36092 19966 36094 20018
rect 36146 19966 36148 20018
rect 36092 19954 36148 19966
rect 36372 19796 36428 19806
rect 35532 19236 35588 19404
rect 35252 19180 35588 19236
rect 35812 19794 36428 19796
rect 35812 19742 36374 19794
rect 36426 19742 36428 19794
rect 35812 19740 36428 19742
rect 35812 19290 35868 19740
rect 36372 19730 36428 19740
rect 35812 19238 35814 19290
rect 35866 19238 35868 19290
rect 35812 19226 35868 19238
rect 35252 19178 35308 19180
rect 35252 19126 35254 19178
rect 35306 19126 35308 19178
rect 35252 19114 35308 19126
rect 35644 19124 35700 19134
rect 35532 19122 35700 19124
rect 35532 19070 35646 19122
rect 35698 19070 35700 19122
rect 35532 19068 35700 19070
rect 35532 18676 35588 19068
rect 35644 19058 35700 19068
rect 33404 18510 33406 18562
rect 33458 18510 33460 18562
rect 33404 18498 33460 18510
rect 35308 18620 35588 18676
rect 35308 18450 35364 18620
rect 35308 18398 35310 18450
rect 35362 18398 35364 18450
rect 35308 18386 35364 18398
rect 35644 18452 35700 18462
rect 34076 18116 34132 18126
rect 33684 17668 33740 17678
rect 33404 17638 33460 17650
rect 33404 17586 33406 17638
rect 33458 17586 33460 17638
rect 33124 17444 33180 17454
rect 33404 17444 33460 17586
rect 33124 17442 33460 17444
rect 33124 17390 33126 17442
rect 33178 17390 33460 17442
rect 33124 17388 33460 17390
rect 33124 17378 33180 17388
rect 32956 16594 33012 16604
rect 33404 15876 33460 17388
rect 33684 17108 33740 17612
rect 33684 17106 33908 17108
rect 33684 17054 33686 17106
rect 33738 17054 33908 17106
rect 33684 17052 33908 17054
rect 33684 17042 33740 17052
rect 33852 16882 33908 17052
rect 33852 16830 33854 16882
rect 33906 16830 33908 16882
rect 33852 16818 33908 16830
rect 33404 15810 33460 15820
rect 32508 15540 32620 15550
rect 32564 15538 32620 15540
rect 32564 15486 32566 15538
rect 32618 15486 32620 15538
rect 32564 15484 32620 15486
rect 32508 15474 32620 15484
rect 32508 15446 32564 15474
rect 31948 15329 32004 15341
rect 31948 15316 31950 15329
rect 32002 15316 32004 15329
rect 31948 15237 32004 15260
rect 32060 15202 32116 15214
rect 32060 15150 32062 15202
rect 32114 15150 32116 15202
rect 31948 14644 32004 14654
rect 32060 14644 32116 15150
rect 31948 14642 32116 14644
rect 31948 14590 31950 14642
rect 32002 14590 32116 14642
rect 31948 14588 32116 14590
rect 32732 15204 32788 15214
rect 34076 15204 34132 18060
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35644 17666 35700 18396
rect 36092 18452 36148 18462
rect 36092 18358 36148 18396
rect 36484 18452 36540 18462
rect 36484 18358 36540 18396
rect 35644 17614 35646 17666
rect 35698 17614 35700 17666
rect 35644 17602 35700 17614
rect 36988 17666 37044 23886
rect 37100 24106 37156 24118
rect 37100 24054 37102 24106
rect 37154 24054 37156 24106
rect 37100 23940 37156 24054
rect 37100 23874 37156 23884
rect 37324 23938 37380 26908
rect 37436 26068 37492 26078
rect 37436 25974 37492 26012
rect 37324 23886 37326 23938
rect 37378 23886 37380 23938
rect 36988 17614 36990 17666
rect 37042 17614 37044 17666
rect 34188 17108 34244 17118
rect 34188 17014 34244 17052
rect 36988 17108 37044 17614
rect 36988 17042 37044 17052
rect 37100 23044 37156 23054
rect 37324 23044 37380 23886
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 37996 23716 38052 23726
rect 37996 23622 38052 23660
rect 37156 22988 37380 23044
rect 37100 16996 37156 22988
rect 37548 21586 37604 21598
rect 37548 21534 37550 21586
rect 37602 21534 37604 21586
rect 37548 21476 37604 21534
rect 37940 21476 37996 21486
rect 37548 21474 37996 21476
rect 37548 21422 37942 21474
rect 37994 21422 37996 21474
rect 37548 21420 37996 21422
rect 37548 20132 37604 21420
rect 37940 21410 37996 21420
rect 37548 18452 37604 20076
rect 37548 18386 37604 18396
rect 38668 20244 38724 20254
rect 38668 18450 38724 20188
rect 38668 18398 38670 18450
rect 38722 18398 38724 18450
rect 38668 18386 38724 18398
rect 37324 18340 37380 18350
rect 37324 17890 37380 18284
rect 38668 18228 38724 18238
rect 37324 17838 37326 17890
rect 37378 17838 37380 17890
rect 37324 17826 37380 17838
rect 37996 17892 38052 17902
rect 38556 17892 38612 17902
rect 37996 17890 38612 17892
rect 37996 17838 37998 17890
rect 38050 17838 38558 17890
rect 38610 17838 38612 17890
rect 37996 17836 38612 17838
rect 37996 17826 38052 17836
rect 37660 17666 37716 17678
rect 37660 17614 37662 17666
rect 37714 17614 37716 17666
rect 37100 16930 37156 16940
rect 37492 16996 37548 17006
rect 37660 16996 37716 17614
rect 37548 16940 37716 16996
rect 37492 16902 37548 16940
rect 38332 16772 38388 16782
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 37996 15652 38052 15662
rect 34412 15372 34692 15428
rect 34244 15204 34300 15214
rect 34412 15204 34468 15372
rect 34636 15358 34692 15372
rect 34636 15306 34638 15358
rect 34690 15306 34692 15358
rect 34636 15294 34692 15306
rect 34972 15316 35028 15326
rect 34972 15222 35028 15260
rect 36316 15316 36372 15326
rect 34076 15202 34468 15204
rect 34076 15150 34246 15202
rect 34298 15150 34468 15202
rect 34076 15148 34468 15150
rect 34524 15204 34580 15214
rect 34524 15202 34804 15204
rect 34524 15150 34526 15202
rect 34578 15150 34804 15202
rect 34524 15148 34804 15150
rect 32732 14644 32788 15148
rect 34244 15138 34300 15148
rect 34524 15138 34580 15148
rect 33124 14644 33180 14654
rect 32732 14642 33180 14644
rect 32732 14590 33126 14642
rect 33178 14590 33180 14642
rect 32732 14588 33180 14590
rect 31948 14578 32004 14588
rect 32732 14530 32788 14588
rect 33124 14578 33180 14588
rect 32732 14478 32734 14530
rect 32786 14478 32788 14530
rect 32732 14466 32788 14478
rect 33796 14532 33852 14542
rect 33796 14438 33852 14476
rect 34076 14532 34132 14542
rect 34076 14438 34132 14476
rect 34188 14503 34468 14532
rect 34188 14476 34414 14503
rect 33628 13748 33684 13758
rect 33628 13654 33684 13692
rect 34188 13076 34244 14476
rect 34412 14451 34414 14476
rect 34466 14451 34468 14503
rect 34748 14530 34804 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34748 14478 34750 14530
rect 34802 14478 34804 14530
rect 34748 14466 34804 14478
rect 34412 14439 34468 14451
rect 34188 13010 34244 13020
rect 34300 14362 34356 14374
rect 34300 14310 34302 14362
rect 34354 14310 34356 14362
rect 34300 12962 34356 14310
rect 36316 13858 36372 15260
rect 37996 15314 38052 15596
rect 38332 15428 38388 16716
rect 38332 15334 38388 15372
rect 37996 15262 37998 15314
rect 38050 15262 38052 15314
rect 37996 15250 38052 15262
rect 38164 15316 38220 15326
rect 38164 15222 38220 15260
rect 38444 15314 38500 17836
rect 38556 17826 38612 17836
rect 38668 16772 38724 18172
rect 38668 16706 38724 16716
rect 38780 15540 38836 27244
rect 39284 27130 39340 27244
rect 39116 27074 39172 27086
rect 39116 27022 39118 27074
rect 39170 27022 39172 27074
rect 39284 27078 39286 27130
rect 39338 27078 39340 27130
rect 39284 27066 39340 27078
rect 39452 27076 39508 27356
rect 39116 26068 39172 27022
rect 39452 26982 39508 27020
rect 39564 27074 39620 27580
rect 39564 27022 39566 27074
rect 39618 27022 39620 27074
rect 39564 27010 39620 27022
rect 39676 27076 39732 28814
rect 39788 27310 39844 29484
rect 39900 27524 39956 30156
rect 40236 30210 40404 30212
rect 40236 30158 40350 30210
rect 40402 30158 40404 30210
rect 40236 30156 40404 30158
rect 40236 30100 40292 30156
rect 40348 30146 40404 30156
rect 40068 29316 40124 29326
rect 40236 29316 40292 30044
rect 41020 29876 41076 30940
rect 41132 30930 41188 30940
rect 41224 30212 41280 30250
rect 41224 30146 41280 30156
rect 41356 29988 41412 32396
rect 41468 32508 41636 32564
rect 41468 31750 41524 32508
rect 41636 32340 41692 32350
rect 41636 32338 41972 32340
rect 41636 32286 41638 32338
rect 41690 32286 41972 32338
rect 41636 32284 41972 32286
rect 41636 32274 41692 32284
rect 41916 31892 41972 32284
rect 41916 31836 42140 31892
rect 42084 31834 42140 31836
rect 41468 31698 41470 31750
rect 41522 31698 41524 31750
rect 41692 31780 41748 31790
rect 42084 31782 42086 31834
rect 42138 31782 42140 31834
rect 41692 31778 41860 31780
rect 41692 31726 41694 31778
rect 41746 31726 41860 31778
rect 42084 31770 42140 31782
rect 41692 31724 41860 31726
rect 41692 31714 41748 31724
rect 41468 30324 41524 31698
rect 41692 31556 41748 31566
rect 41468 30268 41636 30324
rect 40068 29314 40292 29316
rect 40068 29262 40070 29314
rect 40122 29262 40292 29314
rect 40068 29260 40292 29262
rect 40068 29250 40124 29260
rect 39900 27458 39956 27468
rect 40124 28418 40180 28430
rect 40124 28366 40126 28418
rect 40178 28366 40180 28418
rect 39788 27298 39900 27310
rect 39788 27246 39846 27298
rect 39898 27246 39900 27298
rect 39788 27244 39900 27246
rect 39844 27234 39900 27244
rect 39676 27010 39732 27020
rect 40124 27074 40180 28366
rect 40236 27188 40292 29260
rect 40796 29820 41076 29876
rect 41244 29932 41412 29988
rect 41468 30098 41524 30110
rect 41468 30046 41470 30098
rect 41522 30046 41524 30098
rect 40684 28420 40740 28430
rect 40460 28418 40740 28420
rect 40460 28366 40686 28418
rect 40738 28366 40740 28418
rect 40460 28364 40740 28366
rect 40460 27298 40516 28364
rect 40684 28354 40740 28364
rect 40460 27246 40462 27298
rect 40514 27246 40516 27298
rect 40460 27234 40516 27246
rect 40236 27132 40348 27188
rect 40124 27022 40126 27074
rect 40178 27022 40180 27074
rect 39788 26964 39844 26974
rect 39116 24500 39172 26012
rect 39676 26852 39844 26908
rect 40012 26964 40068 26974
rect 38892 24444 39172 24500
rect 39228 24724 39284 24734
rect 38892 18116 38948 24444
rect 39228 23716 39284 24668
rect 39676 23828 39732 26852
rect 40012 23940 40068 26908
rect 40124 24724 40180 27022
rect 40292 26964 40348 27132
rect 40236 26908 40348 26964
rect 40236 26180 40292 26908
rect 40404 26292 40460 26302
rect 40796 26292 40852 29820
rect 41076 28420 41132 28430
rect 40908 27860 40964 27870
rect 40908 27188 40964 27804
rect 41076 27802 41132 28364
rect 41076 27750 41078 27802
rect 41130 27750 41132 27802
rect 41076 27300 41132 27750
rect 41244 27970 41300 29932
rect 41468 28532 41524 30046
rect 41244 27918 41246 27970
rect 41298 27918 41300 27970
rect 41244 27748 41300 27918
rect 41356 28476 41524 28532
rect 41356 27858 41412 28476
rect 41580 28420 41636 30268
rect 41356 27806 41358 27858
rect 41410 27806 41412 27858
rect 41356 27794 41412 27806
rect 41468 28418 41636 28420
rect 41468 28366 41582 28418
rect 41634 28366 41636 28418
rect 41468 28364 41636 28366
rect 41244 27682 41300 27692
rect 41076 27234 41132 27244
rect 40908 27122 40964 27132
rect 41468 27076 41524 28364
rect 41580 28354 41636 28364
rect 41692 28420 41748 31500
rect 41804 30772 41860 31724
rect 41916 31666 41972 31678
rect 41916 31614 41918 31666
rect 41970 31614 41972 31666
rect 41916 30994 41972 31614
rect 41916 30942 41918 30994
rect 41970 30942 41972 30994
rect 41916 30930 41972 30942
rect 42140 30884 42196 30894
rect 41804 30716 42028 30772
rect 41972 30434 42028 30716
rect 41972 30382 41974 30434
rect 42026 30382 42028 30434
rect 41972 30370 42028 30382
rect 42140 30212 42196 30828
rect 43820 30884 43876 30894
rect 43820 30790 43876 30828
rect 42140 30118 42196 30156
rect 41692 28354 41748 28364
rect 41636 27636 41692 27646
rect 41636 27634 42028 27636
rect 41636 27582 41638 27634
rect 41690 27582 42028 27634
rect 41636 27580 42028 27582
rect 41636 27570 41692 27580
rect 41972 27130 42028 27580
rect 41412 27020 41524 27076
rect 41580 27074 41636 27086
rect 41580 27022 41582 27074
rect 41634 27022 41636 27074
rect 41972 27078 41974 27130
rect 42026 27078 42028 27130
rect 41972 27066 42028 27078
rect 41412 27018 41468 27020
rect 41412 26966 41414 27018
rect 41466 26966 41468 27018
rect 41412 26954 41468 26966
rect 41132 26292 41188 26302
rect 40404 26290 41188 26292
rect 40404 26238 40406 26290
rect 40458 26238 41134 26290
rect 41186 26238 41188 26290
rect 40404 26236 41188 26238
rect 40404 26226 40460 26236
rect 41132 26226 41188 26236
rect 40236 26114 40292 26124
rect 40124 24658 40180 24668
rect 41244 25284 41300 25294
rect 40404 23940 40460 23950
rect 40012 23938 40460 23940
rect 40012 23886 40014 23938
rect 40066 23886 40406 23938
rect 40458 23886 40460 23938
rect 40012 23884 40460 23886
rect 40012 23874 40068 23884
rect 40404 23874 40460 23884
rect 39060 22372 39116 22382
rect 39060 22278 39116 22316
rect 39116 20356 39172 20366
rect 39116 18788 39172 20300
rect 39228 19236 39284 23660
rect 39564 23772 39732 23828
rect 39564 23154 39620 23772
rect 39844 23716 39900 23726
rect 39564 23102 39566 23154
rect 39618 23102 39620 23154
rect 39564 23090 39620 23102
rect 39676 23714 39900 23716
rect 39676 23662 39846 23714
rect 39898 23662 39900 23714
rect 39676 23660 39900 23662
rect 39676 22932 39732 23660
rect 39844 23650 39900 23660
rect 39620 22876 39732 22932
rect 39788 23154 39844 23166
rect 39788 23102 39790 23154
rect 39842 23102 39844 23154
rect 39620 22426 39676 22876
rect 39340 22370 39396 22382
rect 39340 22318 39342 22370
rect 39394 22318 39396 22370
rect 39620 22374 39622 22426
rect 39674 22374 39676 22426
rect 39620 22362 39676 22374
rect 39788 22370 39844 23102
rect 39340 21700 39396 22318
rect 39788 22318 39790 22370
rect 39842 22318 39844 22370
rect 39452 22258 39508 22270
rect 39788 22260 39844 22318
rect 39452 22206 39454 22258
rect 39506 22206 39508 22258
rect 39452 21812 39508 22206
rect 39452 21746 39508 21756
rect 39564 22204 39844 22260
rect 40908 22370 40964 22382
rect 40908 22318 40910 22370
rect 40962 22318 40964 22370
rect 39340 21634 39396 21644
rect 39564 21588 39620 22204
rect 40740 22148 40796 22158
rect 40908 22148 40964 22318
rect 41244 22260 41300 25228
rect 41580 25284 41636 27022
rect 41804 26962 41860 26974
rect 41804 26910 41806 26962
rect 41858 26910 41860 26962
rect 41804 26292 41860 26910
rect 41916 26292 41972 26302
rect 41804 26290 41972 26292
rect 41804 26238 41918 26290
rect 41970 26238 41972 26290
rect 41804 26236 41972 26238
rect 41916 26226 41972 26236
rect 43820 26178 43876 26190
rect 43820 26126 43822 26178
rect 43874 26126 43876 26178
rect 42812 25508 42868 25518
rect 42812 25414 42868 25452
rect 43820 25508 43876 26126
rect 43820 25442 43876 25452
rect 41580 25218 41636 25228
rect 42644 25284 42700 25294
rect 42644 25190 42700 25228
rect 41692 22372 41748 22382
rect 40684 22146 40964 22148
rect 40684 22094 40742 22146
rect 40794 22094 40964 22146
rect 40684 22092 40964 22094
rect 41076 22204 41300 22260
rect 41468 22370 41748 22372
rect 41468 22318 41694 22370
rect 41746 22318 41748 22370
rect 41468 22316 41748 22318
rect 40684 22082 40796 22092
rect 39900 21812 39956 21822
rect 39900 21586 39956 21756
rect 39564 21494 39620 21532
rect 39732 21530 39788 21542
rect 39732 21478 39734 21530
rect 39786 21478 39788 21530
rect 39732 21364 39788 21478
rect 39732 21298 39788 21308
rect 39900 21534 39902 21586
rect 39954 21534 39956 21586
rect 39900 20244 39956 21534
rect 40012 21700 40068 21710
rect 40012 21586 40068 21644
rect 40012 21534 40014 21586
rect 40066 21534 40068 21586
rect 40012 20356 40068 21534
rect 40292 21364 40348 21374
rect 40012 20290 40068 20300
rect 40236 21362 40348 21364
rect 40236 21310 40294 21362
rect 40346 21310 40348 21362
rect 40236 21298 40348 21310
rect 39900 20178 39956 20188
rect 40236 19684 40292 21298
rect 40684 20188 40740 22082
rect 41076 21642 41132 22204
rect 40908 21588 40964 21598
rect 41076 21590 41078 21642
rect 41130 21590 41132 21642
rect 41244 21812 41300 21822
rect 41244 21698 41300 21756
rect 41244 21646 41246 21698
rect 41298 21646 41300 21698
rect 41244 21634 41300 21646
rect 41356 21700 41412 21710
rect 41076 21578 41132 21590
rect 41356 21586 41412 21644
rect 40908 21494 40964 21532
rect 41356 21534 41358 21586
rect 41410 21534 41412 21586
rect 41356 21522 41412 21534
rect 41244 21364 41300 21374
rect 41244 20802 41300 21308
rect 41468 20914 41524 22316
rect 41692 22306 41748 22316
rect 43596 22260 43652 22270
rect 42812 22258 43652 22260
rect 42812 22206 43598 22258
rect 43650 22206 43652 22258
rect 42812 22204 43652 22206
rect 42812 21586 42868 22204
rect 43596 22194 43652 22204
rect 42812 21534 42814 21586
rect 42866 21534 42868 21586
rect 42812 21522 42868 21534
rect 41468 20862 41470 20914
rect 41522 20862 41524 20914
rect 41468 20850 41524 20862
rect 41636 21362 41692 21374
rect 41636 21310 41638 21362
rect 41690 21310 41692 21362
rect 41636 20858 41692 21310
rect 42644 21364 42700 21374
rect 42644 21270 42700 21308
rect 40236 19618 40292 19628
rect 40572 20132 40740 20188
rect 40908 20746 40964 20758
rect 40908 20694 40910 20746
rect 40962 20694 40964 20746
rect 41244 20750 41246 20802
rect 41298 20750 41300 20802
rect 41636 20806 41638 20858
rect 41690 20806 41692 20858
rect 41636 20794 41692 20806
rect 41244 20738 41300 20750
rect 39564 19460 39620 19470
rect 39564 19366 39620 19404
rect 39228 19234 39508 19236
rect 39228 19182 39230 19234
rect 39282 19182 39508 19234
rect 39228 19180 39508 19182
rect 39228 19170 39284 19180
rect 39452 18788 39508 19180
rect 39116 18732 39284 18788
rect 39452 18732 39620 18788
rect 39004 18450 39060 18462
rect 39004 18398 39006 18450
rect 39058 18398 39060 18450
rect 39004 18340 39060 18398
rect 39004 18274 39060 18284
rect 39116 18450 39172 18462
rect 39116 18398 39118 18450
rect 39170 18398 39172 18450
rect 38892 18060 39060 18116
rect 39004 16882 39060 18060
rect 39116 17890 39172 18398
rect 39228 18452 39284 18732
rect 39452 18452 39508 18462
rect 39228 18450 39508 18452
rect 39228 18398 39454 18450
rect 39506 18398 39508 18450
rect 39228 18396 39508 18398
rect 39452 18386 39508 18396
rect 39116 17838 39118 17890
rect 39170 17838 39172 17890
rect 39116 17826 39172 17838
rect 39340 18228 39396 18238
rect 39340 17556 39396 18172
rect 39004 16830 39006 16882
rect 39058 16830 39060 16882
rect 39172 17500 39396 17556
rect 39452 17890 39508 17902
rect 39452 17838 39454 17890
rect 39506 17838 39508 17890
rect 39172 16938 39228 17500
rect 39172 16886 39174 16938
rect 39226 16886 39228 16938
rect 39172 16874 39228 16886
rect 39340 16882 39396 16894
rect 39004 15652 39060 16830
rect 39340 16830 39342 16882
rect 39394 16830 39396 16882
rect 39340 16772 39396 16830
rect 39452 16882 39508 17838
rect 39452 16830 39454 16882
rect 39506 16830 39508 16882
rect 39452 16818 39508 16830
rect 39340 16706 39396 16716
rect 39564 16098 39620 18732
rect 40572 17892 40628 20076
rect 40740 19684 40796 19694
rect 40740 19290 40796 19628
rect 40908 19460 40964 20694
rect 40908 19394 40964 19404
rect 41356 19460 41412 19470
rect 40740 19238 40742 19290
rect 40794 19238 40796 19290
rect 40740 19226 40796 19238
rect 41132 19234 41188 19246
rect 41132 19182 41134 19234
rect 41186 19182 41188 19234
rect 40908 19122 40964 19134
rect 40908 19070 40910 19122
rect 40962 19070 40964 19122
rect 40908 18228 40964 19070
rect 41132 18686 41188 19182
rect 41356 19206 41412 19404
rect 41356 19154 41358 19206
rect 41410 19154 41412 19206
rect 41356 19142 41412 19154
rect 41132 18674 41244 18686
rect 41132 18622 41190 18674
rect 41242 18622 41244 18674
rect 41132 18620 41244 18622
rect 41188 18610 41244 18620
rect 41020 18452 41076 18462
rect 41020 18358 41076 18396
rect 43596 18452 43652 18462
rect 40908 18172 41748 18228
rect 40348 17836 40796 17892
rect 39732 16660 39788 16670
rect 39732 16658 40180 16660
rect 39732 16606 39734 16658
rect 39786 16606 40180 16658
rect 39732 16604 40180 16606
rect 39732 16594 39788 16604
rect 39564 16046 39566 16098
rect 39618 16046 39620 16098
rect 39564 16034 39620 16046
rect 39228 15876 39284 15886
rect 39228 15874 39732 15876
rect 39228 15822 39230 15874
rect 39282 15822 39732 15874
rect 39228 15820 39732 15822
rect 39228 15810 39284 15820
rect 39004 15586 39060 15596
rect 39340 15652 39396 15662
rect 38780 15474 38836 15484
rect 39004 15428 39060 15438
rect 38444 15262 38446 15314
rect 38498 15262 38500 15314
rect 38444 15204 38500 15262
rect 38724 15316 38780 15326
rect 38724 15222 38780 15260
rect 38444 15138 38500 15148
rect 38892 15204 38948 15214
rect 38892 14530 38948 15148
rect 38892 14478 38894 14530
rect 38946 14478 38948 14530
rect 38892 14466 38948 14478
rect 39004 14530 39060 15372
rect 39004 14478 39006 14530
rect 39058 14478 39060 14530
rect 39340 14530 39396 15596
rect 39564 15540 39620 15550
rect 39564 15314 39620 15484
rect 39564 15262 39566 15314
rect 39618 15262 39620 15314
rect 39564 15250 39620 15262
rect 39676 15314 39732 15820
rect 39676 15262 39678 15314
rect 39730 15262 39732 15314
rect 39004 14466 39060 14478
rect 39172 14474 39228 14486
rect 36316 13806 36318 13858
rect 36370 13806 36372 13858
rect 36316 13794 36372 13806
rect 36932 14420 36988 14430
rect 36932 13970 36988 14364
rect 38612 14420 38668 14430
rect 39172 14422 39174 14474
rect 39226 14422 39228 14474
rect 39340 14478 39342 14530
rect 39394 14478 39396 14530
rect 39340 14466 39396 14478
rect 38612 14418 38836 14420
rect 38612 14366 38614 14418
rect 38666 14366 38836 14418
rect 38612 14364 38836 14366
rect 38612 14354 38668 14364
rect 36932 13918 36934 13970
rect 36986 13918 36988 13970
rect 36932 13748 36988 13918
rect 36876 13692 36932 13748
rect 36876 13682 36988 13692
rect 34412 13636 34468 13646
rect 34412 13634 34692 13636
rect 34412 13582 34414 13634
rect 34466 13582 34692 13634
rect 34412 13580 34692 13582
rect 34412 13570 34468 13580
rect 34636 13186 34692 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34636 13134 34638 13186
rect 34690 13134 34692 13186
rect 34636 13122 34692 13134
rect 34300 12910 34302 12962
rect 34354 12910 34356 12962
rect 34300 12898 34356 12910
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 36708 10836 36764 10846
rect 36876 10836 36932 13682
rect 38220 13076 38276 13086
rect 38220 12982 38276 13020
rect 38668 12962 38724 12974
rect 38332 12918 38388 12930
rect 38332 12866 38334 12918
rect 38386 12866 38388 12918
rect 38332 12180 38388 12866
rect 38668 12910 38670 12962
rect 38722 12910 38724 12962
rect 38668 12180 38724 12910
rect 38780 12292 38836 14364
rect 39172 13860 39228 14422
rect 39676 13860 39732 15262
rect 39822 15351 39878 15363
rect 39822 15316 39824 15351
rect 39876 15316 39878 15351
rect 39822 15250 39878 15260
rect 39172 13804 39284 13860
rect 39676 13804 40068 13860
rect 39228 12964 39284 13804
rect 39228 12898 39284 12908
rect 39900 12964 39956 12974
rect 39900 12870 39956 12908
rect 40012 12962 40068 13804
rect 40012 12910 40014 12962
rect 40066 12910 40068 12962
rect 38780 12236 39210 12292
rect 39154 12216 39210 12236
rect 38668 12124 39060 12180
rect 39154 12164 39156 12216
rect 39208 12164 39210 12216
rect 39154 12152 39210 12164
rect 39340 12180 39396 12190
rect 38332 12114 38388 12124
rect 38780 11956 38836 11966
rect 39004 11956 39060 12124
rect 39340 12086 39396 12124
rect 39452 12180 39508 12190
rect 40012 12180 40068 12910
rect 40124 12974 40180 16604
rect 40236 15092 40292 15102
rect 40236 14998 40292 15036
rect 40348 14654 40404 17836
rect 40740 17780 40796 17836
rect 40740 17778 40964 17780
rect 40740 17726 40742 17778
rect 40794 17726 40964 17778
rect 40740 17724 40964 17726
rect 40740 17714 40796 17724
rect 40908 17666 40964 17724
rect 41692 17778 41748 18172
rect 41692 17726 41694 17778
rect 41746 17726 41748 17778
rect 41692 17714 41748 17726
rect 43596 17778 43652 18396
rect 43596 17726 43598 17778
rect 43650 17726 43652 17778
rect 43596 17714 43652 17726
rect 40908 17614 40910 17666
rect 40962 17614 40964 17666
rect 40908 17602 40964 17614
rect 43820 15540 43876 15550
rect 40292 14642 40404 14654
rect 40292 14590 40294 14642
rect 40346 14590 40404 14642
rect 40292 14578 40404 14590
rect 40348 14532 40404 14578
rect 40348 14466 40404 14476
rect 40460 15092 40516 15102
rect 41020 15092 41076 15102
rect 40460 14530 40516 15036
rect 40796 15090 41076 15092
rect 40796 15038 41022 15090
rect 41074 15038 41076 15090
rect 40796 15036 41076 15038
rect 40796 14754 40852 15036
rect 41020 15026 41076 15036
rect 41916 15090 41972 15102
rect 41916 15038 41918 15090
rect 41970 15038 41972 15090
rect 40796 14702 40798 14754
rect 40850 14702 40852 14754
rect 40796 14690 40852 14702
rect 41916 14642 41972 15038
rect 41916 14590 41918 14642
rect 41970 14590 41972 14642
rect 41916 14578 41972 14590
rect 43820 14642 43876 15484
rect 43820 14590 43822 14642
rect 43874 14590 43876 14642
rect 43820 14578 43876 14590
rect 41132 14532 41188 14542
rect 40460 14478 40462 14530
rect 40514 14478 40516 14530
rect 40460 14466 40516 14478
rect 41020 14476 41132 14532
rect 40572 13074 40628 13086
rect 40572 13022 40574 13074
rect 40626 13022 40628 13074
rect 40124 12962 40234 12974
rect 40124 12910 40180 12962
rect 40232 12910 40234 12962
rect 40124 12908 40234 12910
rect 40178 12898 40234 12908
rect 39452 12178 39620 12180
rect 39452 12126 39454 12178
rect 39506 12126 39620 12178
rect 39452 12124 39620 12126
rect 39452 11956 39508 12124
rect 38780 11954 38948 11956
rect 38780 11902 38782 11954
rect 38834 11902 38948 11954
rect 38780 11900 38948 11902
rect 39004 11900 39508 11956
rect 38780 11890 38836 11900
rect 38892 11394 38948 11900
rect 38892 11342 38894 11394
rect 38946 11342 38948 11394
rect 38892 11330 38948 11342
rect 38556 11172 38612 11182
rect 36708 10834 36932 10836
rect 36708 10782 36710 10834
rect 36762 10782 36932 10834
rect 36708 10780 36932 10782
rect 36708 10770 36764 10780
rect 30548 9940 30604 9950
rect 30548 9846 30604 9884
rect 30940 9826 30996 10108
rect 31724 10108 31892 10164
rect 32172 10612 32228 10622
rect 30940 9774 30942 9826
rect 30994 9774 30996 9826
rect 31612 9826 31668 9838
rect 30940 9762 30996 9774
rect 31388 9770 31444 9782
rect 28588 9650 28644 9660
rect 31388 9718 31390 9770
rect 31442 9718 31444 9770
rect 27468 9212 27636 9268
rect 27412 9174 27468 9212
rect 31388 9044 31444 9718
rect 31388 8978 31444 8988
rect 31612 9774 31614 9826
rect 31666 9774 31668 9826
rect 27244 6142 27300 8540
rect 31612 6916 31668 9774
rect 31724 9658 31780 10108
rect 31724 9606 31726 9658
rect 31778 9606 31780 9658
rect 32060 9826 32116 9838
rect 32060 9774 32062 9826
rect 32114 9774 32116 9826
rect 32060 9716 32116 9774
rect 32060 9650 32116 9660
rect 32172 9660 32228 10556
rect 32956 10612 33012 10622
rect 33180 10612 33236 10622
rect 32956 10518 33012 10556
rect 33068 10610 33236 10612
rect 33068 10558 33182 10610
rect 33234 10558 33236 10610
rect 33068 10556 33236 10558
rect 33068 10164 33124 10556
rect 33180 10546 33236 10556
rect 36876 10610 36932 10780
rect 36876 10558 36878 10610
rect 36930 10558 36932 10610
rect 33460 10388 33516 10398
rect 33460 10386 33572 10388
rect 33460 10334 33462 10386
rect 33514 10334 33572 10386
rect 33460 10322 33572 10334
rect 32564 10108 33124 10164
rect 32564 10050 32620 10108
rect 32564 9998 32566 10050
rect 32618 9998 32620 10050
rect 32564 9986 32620 9998
rect 33516 9940 33572 10322
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 36876 10052 36932 10558
rect 37660 11170 38612 11172
rect 37660 11118 38558 11170
rect 38610 11118 38612 11170
rect 37660 11116 38612 11118
rect 37660 10610 37716 11116
rect 38556 11106 38612 11116
rect 39564 10722 39620 12124
rect 40012 12114 40068 12124
rect 40572 12180 40628 13022
rect 40572 12114 40628 12124
rect 40852 11508 40908 11518
rect 41020 11508 41076 14476
rect 41132 14438 41188 14476
rect 43708 12964 43764 12974
rect 41132 12180 41188 12190
rect 41132 12086 41188 12124
rect 41468 11956 41524 11966
rect 41468 11954 41860 11956
rect 41468 11902 41470 11954
rect 41522 11902 41860 11954
rect 41468 11900 41860 11902
rect 41468 11890 41524 11900
rect 40852 11506 41076 11508
rect 40852 11454 40854 11506
rect 40906 11454 41076 11506
rect 40852 11452 41076 11454
rect 40852 11442 40908 11452
rect 41020 11394 41076 11452
rect 41804 11506 41860 11900
rect 41804 11454 41806 11506
rect 41858 11454 41860 11506
rect 41804 11442 41860 11454
rect 43708 11506 43764 12908
rect 43708 11454 43710 11506
rect 43762 11454 43764 11506
rect 43708 11442 43764 11454
rect 41020 11342 41022 11394
rect 41074 11342 41076 11394
rect 41020 11330 41076 11342
rect 39564 10670 39566 10722
rect 39618 10670 39620 10722
rect 39564 10658 39620 10670
rect 37660 10558 37662 10610
rect 37714 10558 37716 10610
rect 37660 10546 37716 10558
rect 36876 9996 37212 10052
rect 33516 9884 33796 9940
rect 32284 9828 32340 9838
rect 32284 9826 33180 9828
rect 32284 9774 32286 9826
rect 32338 9774 33180 9826
rect 32284 9772 33180 9774
rect 32284 9762 32340 9772
rect 31724 9594 31780 9606
rect 32172 9604 32340 9660
rect 31220 6860 31668 6916
rect 32172 9044 32228 9054
rect 30828 6692 30884 6702
rect 30828 6598 30884 6636
rect 30940 6690 30996 6702
rect 30940 6638 30942 6690
rect 30994 6638 30996 6690
rect 27188 6132 27300 6142
rect 27188 6130 27244 6132
rect 27188 6078 27190 6130
rect 27242 6078 27244 6130
rect 27188 6076 27244 6078
rect 27188 6066 27300 6076
rect 27244 6038 27300 6066
rect 27580 6356 27636 6366
rect 27580 5950 27636 6300
rect 29596 6356 29652 6366
rect 28252 6132 28308 6142
rect 27580 5898 27582 5950
rect 27634 5898 27636 5950
rect 27580 5886 27636 5898
rect 27916 6020 27972 6030
rect 27916 5906 27972 5964
rect 27916 5854 27918 5906
rect 27970 5854 27972 5906
rect 27916 5842 27972 5854
rect 28252 5906 28308 6076
rect 28252 5854 28254 5906
rect 28306 5854 28308 5906
rect 28252 5842 28308 5854
rect 28476 6074 28532 6086
rect 28476 6022 28478 6074
rect 28530 6022 28532 6074
rect 27468 5796 27524 5806
rect 27468 5702 27524 5740
rect 25900 5122 26628 5124
rect 25900 5070 25902 5122
rect 25954 5070 26294 5122
rect 26346 5070 26628 5122
rect 25900 5068 26628 5070
rect 28476 5122 28532 6022
rect 29484 6020 29540 6030
rect 28588 5933 28644 5945
rect 28588 5881 28590 5933
rect 28642 5881 28644 5933
rect 28588 5796 28644 5881
rect 28588 5730 28644 5740
rect 28924 5906 28980 5918
rect 28924 5854 28926 5906
rect 28978 5854 28980 5906
rect 28924 5796 28980 5854
rect 28924 5730 28980 5740
rect 29484 5906 29540 5964
rect 29484 5854 29486 5906
rect 29538 5854 29540 5906
rect 28476 5070 28478 5122
rect 28530 5070 28532 5122
rect 25900 5058 25956 5068
rect 24220 4620 24948 4676
rect 24220 4562 24276 4620
rect 24220 4510 24222 4562
rect 24274 4510 24276 4562
rect 24220 4498 24276 4510
rect 23884 4286 23886 4338
rect 23938 4286 23940 4338
rect 23884 4274 23940 4286
rect 26292 4340 26348 5068
rect 28476 5058 28532 5070
rect 28140 4900 28196 4910
rect 27692 4898 28196 4900
rect 27692 4846 28142 4898
rect 28194 4846 28196 4898
rect 27692 4844 28196 4846
rect 26292 4274 26348 4284
rect 26908 4340 26964 4350
rect 26908 4246 26964 4284
rect 27692 4338 27748 4844
rect 28140 4834 28196 4844
rect 29484 4452 29540 5854
rect 29596 5906 29652 6300
rect 30772 6132 30828 6142
rect 30772 6038 30828 6076
rect 30940 6020 30996 6638
rect 31220 6690 31276 6860
rect 31220 6638 31222 6690
rect 31274 6638 31276 6690
rect 31220 6626 31276 6638
rect 31388 6692 31444 6702
rect 31500 6692 31556 6702
rect 31724 6692 31780 6702
rect 32004 6692 32060 6702
rect 32172 6692 32228 8988
rect 32284 8874 32340 9604
rect 32396 9156 32452 9166
rect 32396 9042 32452 9100
rect 33124 9154 33180 9772
rect 33124 9102 33126 9154
rect 33178 9102 33180 9154
rect 33124 9090 33180 9102
rect 33516 9714 33572 9726
rect 33516 9662 33518 9714
rect 33570 9662 33572 9714
rect 33516 9156 33572 9662
rect 32396 8990 32398 9042
rect 32450 8990 32452 9042
rect 32396 8978 32452 8990
rect 33404 9044 33460 9054
rect 33404 8950 33460 8988
rect 33516 9042 33572 9100
rect 33516 8990 33518 9042
rect 33570 8990 33572 9042
rect 33516 8978 33572 8990
rect 33740 9042 33796 9884
rect 35420 9826 35476 9838
rect 35420 9774 35422 9826
rect 35474 9774 35476 9826
rect 34076 9268 34132 9278
rect 34076 9174 34132 9212
rect 35420 9268 35476 9774
rect 35420 9202 35476 9212
rect 36204 9828 36260 9838
rect 33740 8990 33742 9042
rect 33794 8990 33796 9042
rect 33740 8978 33796 8990
rect 32284 8822 32286 8874
rect 32338 8822 32340 8874
rect 32284 8810 32340 8822
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 31444 6690 31556 6692
rect 31444 6638 31502 6690
rect 31554 6638 31556 6690
rect 31444 6636 31556 6638
rect 30940 5954 30996 5964
rect 31052 6132 31108 6142
rect 29596 5854 29598 5906
rect 29650 5854 29652 5906
rect 29596 5842 29652 5854
rect 31052 5906 31108 6076
rect 31052 5854 31054 5906
rect 31106 5854 31108 5906
rect 31052 5842 31108 5854
rect 29876 5796 29932 5806
rect 29876 5702 29932 5740
rect 31276 5124 31332 5134
rect 31388 5124 31444 6636
rect 31500 6626 31556 6636
rect 31612 6690 31780 6692
rect 31612 6638 31726 6690
rect 31778 6638 31780 6690
rect 31612 6636 31780 6638
rect 31500 5945 31556 5957
rect 31500 5893 31502 5945
rect 31554 5893 31556 5945
rect 31500 5236 31556 5893
rect 31612 5796 31668 6636
rect 31724 6626 31780 6636
rect 31836 6690 32228 6692
rect 31836 6638 32006 6690
rect 32058 6638 32228 6690
rect 31836 6636 32228 6638
rect 31836 6468 31892 6636
rect 32004 6598 32060 6636
rect 31724 6412 31892 6468
rect 31724 5906 31780 6412
rect 31724 5854 31726 5906
rect 31778 5854 31780 5906
rect 31724 5842 31780 5854
rect 31836 6074 31892 6086
rect 31836 6022 31838 6074
rect 31890 6022 31892 6074
rect 31836 5908 31892 6022
rect 31836 5842 31892 5852
rect 32956 5908 33012 5918
rect 32956 5814 33012 5852
rect 31612 5460 31668 5740
rect 33292 5684 33348 5694
rect 33292 5590 33348 5628
rect 34076 5684 34132 5694
rect 31612 5404 31780 5460
rect 31612 5236 31668 5246
rect 31500 5234 31668 5236
rect 31500 5182 31614 5234
rect 31666 5182 31668 5234
rect 31500 5180 31668 5182
rect 31612 5170 31668 5180
rect 31332 5068 31444 5124
rect 31556 5092 31612 5104
rect 31276 5030 31332 5068
rect 31556 5040 31558 5092
rect 31610 5040 31612 5092
rect 31556 5012 31612 5040
rect 31724 5012 31780 5404
rect 34076 5234 34132 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34076 5182 34078 5234
rect 34130 5182 34132 5234
rect 34076 5170 34132 5182
rect 34860 5236 34916 5246
rect 32172 5124 32228 5134
rect 32172 5030 32228 5068
rect 34860 5122 34916 5180
rect 35252 5236 35308 5246
rect 35252 5142 35308 5180
rect 36204 5236 36260 9772
rect 36876 9828 36932 9996
rect 37156 9938 37212 9996
rect 37156 9886 37158 9938
rect 37210 9886 37212 9938
rect 37156 9874 37212 9886
rect 36876 9762 36932 9772
rect 36204 5170 36260 5180
rect 34860 5070 34862 5122
rect 34914 5070 34916 5122
rect 34860 5058 34916 5070
rect 31556 4956 31780 5012
rect 29596 4452 29652 4462
rect 29484 4450 29652 4452
rect 29484 4398 29598 4450
rect 29650 4398 29652 4450
rect 29484 4396 29652 4398
rect 29596 4386 29652 4396
rect 27692 4286 27694 4338
rect 27746 4286 27748 4338
rect 27692 4274 27748 4286
rect 30212 4340 30268 4350
rect 30212 4246 30268 4284
rect 18396 4162 18452 4172
rect 19964 4228 20020 4238
rect 19964 4134 20020 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
<< via2 >>
rect 13244 41804 13300 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 2156 40402 2212 40404
rect 2156 40350 2158 40402
rect 2158 40350 2210 40402
rect 2210 40350 2212 40402
rect 2156 40348 2212 40350
rect 5460 40402 5516 40404
rect 5460 40350 5462 40402
rect 5462 40350 5514 40402
rect 5514 40350 5516 40402
rect 5460 40348 5516 40350
rect 5740 40402 5796 40404
rect 5740 40350 5742 40402
rect 5742 40350 5794 40402
rect 5794 40350 5796 40402
rect 5740 40348 5796 40350
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 3052 39564 3108 39620
rect 2660 38834 2716 38836
rect 2660 38782 2662 38834
rect 2662 38782 2714 38834
rect 2714 38782 2716 38834
rect 2660 38780 2716 38782
rect 4060 39564 4116 39620
rect 3948 38668 4004 38724
rect 3276 38556 3332 38612
rect 3836 38556 3892 38612
rect 4620 39618 4676 39620
rect 4620 39566 4622 39618
rect 4622 39566 4674 39618
rect 4674 39566 4676 39618
rect 4620 39564 4676 39566
rect 5068 40236 5124 40292
rect 4844 39564 4900 39620
rect 4284 38892 4340 38948
rect 4508 38834 4564 38836
rect 4508 38782 4510 38834
rect 4510 38782 4562 38834
rect 4562 38782 4564 38834
rect 4508 38780 4564 38782
rect 4172 38556 4228 38612
rect 3948 37266 4004 37268
rect 3948 37214 3950 37266
rect 3950 37214 4002 37266
rect 4002 37214 4004 37266
rect 3948 37212 4004 37214
rect 5292 38892 5348 38948
rect 5068 38668 5124 38724
rect 4676 38556 4732 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4342 37772 4398 37828
rect 4060 37100 4116 37156
rect 5124 37826 5180 37828
rect 5124 37774 5126 37826
rect 5126 37774 5178 37826
rect 5178 37774 5180 37826
rect 5124 37772 5180 37774
rect 4688 37100 4744 37156
rect 4844 37212 4900 37268
rect 3276 33852 3332 33908
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4172 33852 4228 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4284 32562 4340 32564
rect 4284 32510 4286 32562
rect 4286 32510 4338 32562
rect 4338 32510 4340 32562
rect 4284 32508 4340 32510
rect 4508 32508 4564 32564
rect 5124 37266 5180 37268
rect 5124 37214 5126 37266
rect 5126 37214 5178 37266
rect 5178 37214 5180 37266
rect 5124 37212 5180 37214
rect 4956 34130 5012 34132
rect 4956 34078 4958 34130
rect 4958 34078 5010 34130
rect 5010 34078 5012 34130
rect 4956 34076 5012 34078
rect 5628 34130 5684 34132
rect 5628 34078 5630 34130
rect 5630 34078 5682 34130
rect 5682 34078 5684 34130
rect 5628 34076 5684 34078
rect 5124 33458 5180 33460
rect 5124 33406 5126 33458
rect 5126 33406 5178 33458
rect 5178 33406 5180 33458
rect 5124 33404 5180 33406
rect 4620 32396 4676 32452
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 3724 29389 3726 29428
rect 3726 29389 3778 29428
rect 3778 29389 3780 29428
rect 3724 29372 3780 29389
rect 2604 29260 2660 29316
rect 3612 29314 3668 29316
rect 3612 29262 3614 29314
rect 3614 29262 3666 29314
rect 3666 29262 3668 29314
rect 3612 29260 3668 29262
rect 1820 28642 1876 28644
rect 1820 28590 1822 28642
rect 1822 28590 1874 28642
rect 1874 28590 1876 28642
rect 1820 28588 1876 28590
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4060 27916 4116 27972
rect 4508 28364 4564 28420
rect 4956 31164 5012 31220
rect 5404 33404 5460 33460
rect 5516 33740 5572 33796
rect 5292 32732 5348 32788
rect 5404 33180 5460 33236
rect 5124 28642 5180 28644
rect 5124 28590 5126 28642
rect 5126 28590 5178 28642
rect 5178 28590 5180 28642
rect 5124 28588 5180 28590
rect 4844 28028 4900 28084
rect 1932 24556 1988 24612
rect 4172 23996 4228 24052
rect 1708 23212 1764 23268
rect 3948 22428 4004 22484
rect 5068 28364 5124 28420
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4620 24722 4676 24724
rect 4620 24670 4622 24722
rect 4622 24670 4674 24722
rect 4674 24670 4676 24722
rect 4620 24668 4676 24670
rect 6636 40348 6692 40404
rect 6524 40290 6580 40292
rect 6524 40238 6526 40290
rect 6526 40238 6578 40290
rect 6578 40238 6580 40290
rect 6524 40236 6580 40238
rect 6412 37772 6468 37828
rect 6412 34914 6468 34916
rect 6412 34862 6414 34914
rect 6414 34862 6466 34914
rect 6466 34862 6468 34914
rect 6412 34860 6468 34862
rect 6188 33964 6244 34020
rect 5628 33068 5684 33124
rect 5852 33292 5908 33348
rect 6412 33740 6468 33796
rect 7756 38946 7812 38948
rect 7756 38894 7758 38946
rect 7758 38894 7810 38946
rect 7810 38894 7812 38946
rect 7756 38892 7812 38894
rect 8092 38834 8148 38836
rect 8092 38782 8094 38834
rect 8094 38782 8146 38834
rect 8146 38782 8148 38834
rect 8092 38780 8148 38782
rect 8764 39506 8820 39508
rect 8764 39454 8766 39506
rect 8766 39454 8818 39506
rect 8818 39454 8820 39506
rect 8764 39452 8820 39454
rect 8428 38780 8484 38836
rect 6860 37100 6916 37156
rect 6636 35922 6692 35924
rect 6636 35870 6638 35922
rect 6638 35870 6690 35922
rect 6690 35870 6692 35922
rect 6636 35868 6692 35870
rect 7308 35868 7364 35924
rect 7028 34914 7084 34916
rect 7028 34862 7030 34914
rect 7030 34862 7082 34914
rect 7082 34862 7084 34914
rect 7028 34860 7084 34862
rect 6524 33516 6580 33572
rect 6804 33852 6860 33908
rect 6412 33404 6468 33460
rect 8764 33346 8820 33348
rect 8764 33294 8766 33346
rect 8766 33294 8818 33346
rect 8818 33294 8820 33346
rect 8764 33292 8820 33294
rect 6524 33068 6580 33124
rect 5516 30828 5572 30884
rect 5236 24610 5292 24612
rect 5236 24558 5238 24610
rect 5238 24558 5290 24610
rect 5290 24558 5292 24610
rect 5236 24556 5292 24558
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4620 23996 4676 24052
rect 4900 24050 4956 24052
rect 4900 23998 4902 24050
rect 4902 23998 4954 24050
rect 4954 23998 4956 24050
rect 4900 23996 4956 23998
rect 5068 23548 5124 23604
rect 4284 22652 4340 22708
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4620 22482 4676 22484
rect 4620 22430 4622 22482
rect 4622 22430 4674 22482
rect 4674 22430 4676 22482
rect 4620 22428 4676 22430
rect 5628 31218 5684 31220
rect 5628 31166 5630 31218
rect 5630 31166 5682 31218
rect 5682 31166 5684 31218
rect 5628 31164 5684 31166
rect 5852 32732 5908 32788
rect 6300 32549 6302 32564
rect 6302 32549 6354 32564
rect 6354 32549 6356 32564
rect 6300 32508 6356 32549
rect 5852 29372 5908 29428
rect 5684 27970 5740 27972
rect 5684 27918 5686 27970
rect 5686 27918 5738 27970
rect 5738 27918 5740 27970
rect 5684 27916 5740 27918
rect 5516 23996 5572 24052
rect 5740 24892 5796 24948
rect 6524 29372 6580 29428
rect 8428 33122 8484 33124
rect 8428 33070 8430 33122
rect 8430 33070 8482 33122
rect 8482 33070 8484 33122
rect 8428 33068 8484 33070
rect 6860 32508 6916 32564
rect 7252 32450 7308 32452
rect 7252 32398 7254 32450
rect 7254 32398 7306 32450
rect 7306 32398 7308 32450
rect 7252 32396 7308 32398
rect 7756 30940 7812 30996
rect 11788 40572 11844 40628
rect 14476 41858 14532 41860
rect 14476 41806 14478 41858
rect 14478 41806 14530 41858
rect 14530 41806 14532 41858
rect 14476 41804 14532 41806
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 17052 41804 17108 41860
rect 13468 40572 13524 40628
rect 15820 40460 15876 40516
rect 9044 40402 9100 40404
rect 9044 40350 9046 40402
rect 9046 40350 9098 40402
rect 9098 40350 9100 40402
rect 9044 40348 9100 40350
rect 13468 40348 13524 40404
rect 14476 40402 14532 40404
rect 14476 40350 14478 40402
rect 14478 40350 14530 40402
rect 14530 40350 14532 40402
rect 14476 40348 14532 40350
rect 9007 39618 9063 39620
rect 9007 39566 9009 39618
rect 9009 39566 9061 39618
rect 9061 39566 9063 39618
rect 9007 39564 9063 39566
rect 9884 38780 9940 38836
rect 10332 38780 10388 38836
rect 10892 39452 10948 39508
rect 10108 36370 10164 36372
rect 10108 36318 10110 36370
rect 10110 36318 10162 36370
rect 10162 36318 10164 36370
rect 10108 36316 10164 36318
rect 10780 36316 10836 36372
rect 10780 35698 10836 35700
rect 10780 35646 10782 35698
rect 10782 35646 10834 35698
rect 10834 35646 10836 35698
rect 10780 35644 10836 35646
rect 12236 39004 12292 39060
rect 18284 41858 18340 41860
rect 18284 41806 18286 41858
rect 18286 41806 18338 41858
rect 18338 41806 18340 41858
rect 18284 41804 18340 41806
rect 20860 41804 20916 41860
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 17276 40460 17332 40516
rect 22092 41858 22148 41860
rect 22092 41806 22094 41858
rect 22094 41806 22146 41858
rect 22146 41806 22148 41858
rect 22092 41804 22148 41806
rect 24668 41804 24724 41860
rect 25900 41858 25956 41860
rect 25900 41806 25902 41858
rect 25902 41806 25954 41858
rect 25954 41806 25956 41858
rect 25900 41804 25956 41806
rect 28476 41804 28532 41860
rect 29708 41858 29764 41860
rect 29708 41806 29710 41858
rect 29710 41806 29762 41858
rect 29762 41806 29764 41858
rect 29708 41804 29764 41806
rect 32284 41804 32340 41860
rect 33516 41858 33572 41860
rect 33516 41806 33518 41858
rect 33518 41806 33570 41858
rect 33570 41806 33572 41858
rect 33516 41804 33572 41806
rect 36092 41804 36148 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 37324 41858 37380 41860
rect 37324 41806 37326 41858
rect 37326 41806 37378 41858
rect 37378 41806 37380 41858
rect 37324 41804 37380 41806
rect 39900 41804 39956 41860
rect 18396 40402 18452 40404
rect 18396 40350 18398 40402
rect 18398 40350 18450 40402
rect 18450 40350 18452 40402
rect 18396 40348 18452 40350
rect 17724 39730 17780 39732
rect 17724 39678 17726 39730
rect 17726 39678 17778 39730
rect 17778 39678 17780 39730
rect 17724 39676 17780 39678
rect 14252 39618 14308 39620
rect 14252 39566 14254 39618
rect 14254 39566 14306 39618
rect 14306 39566 14308 39618
rect 14252 39564 14308 39566
rect 21868 40402 21924 40404
rect 21868 40350 21870 40402
rect 21870 40350 21922 40402
rect 21922 40350 21924 40402
rect 21868 40348 21924 40350
rect 19180 39788 19236 39844
rect 20188 39842 20244 39844
rect 20188 39790 20190 39842
rect 20190 39790 20242 39842
rect 20242 39790 20244 39842
rect 20188 39788 20244 39790
rect 20524 39452 20580 39508
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 16044 39058 16100 39060
rect 16044 39006 16046 39058
rect 16046 39006 16098 39058
rect 16098 39006 16100 39058
rect 16044 39004 16100 39006
rect 13468 38834 13524 38836
rect 13468 38782 13470 38834
rect 13470 38782 13522 38834
rect 13522 38782 13524 38834
rect 13468 38780 13524 38782
rect 9212 33292 9268 33348
rect 8764 30940 8820 30996
rect 8316 30210 8372 30212
rect 8316 30158 8318 30210
rect 8318 30158 8370 30210
rect 8370 30158 8372 30210
rect 8316 30156 8372 30158
rect 6972 29426 7028 29428
rect 6972 29374 6974 29426
rect 6974 29374 7026 29426
rect 7026 29374 7028 29426
rect 6972 29372 7028 29374
rect 6636 28812 6692 28868
rect 6300 28700 6356 28756
rect 6132 28082 6188 28084
rect 6132 28030 6134 28082
rect 6134 28030 6186 28082
rect 6186 28030 6188 28082
rect 6132 28028 6188 28030
rect 7420 27074 7476 27076
rect 7420 27022 7422 27074
rect 7422 27022 7474 27074
rect 7474 27022 7476 27074
rect 7420 27020 7476 27022
rect 5740 23548 5796 23604
rect 5068 22428 5124 22484
rect 4844 22316 4900 22372
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 4620 20860 4676 20916
rect 6748 24946 6804 24948
rect 6748 24894 6750 24946
rect 6750 24894 6802 24946
rect 6802 24894 6804 24946
rect 6748 24892 6804 24894
rect 5684 22594 5740 22596
rect 5684 22542 5686 22594
rect 5686 22542 5738 22594
rect 5738 22542 5740 22594
rect 5684 22540 5740 22542
rect 5404 21756 5460 21812
rect 5628 20914 5684 20916
rect 5628 20862 5630 20914
rect 5630 20862 5682 20914
rect 5682 20862 5684 20914
rect 5628 20860 5684 20862
rect 6076 22428 6132 22484
rect 5964 22370 6020 22372
rect 5964 22318 5966 22370
rect 5966 22318 6018 22370
rect 6018 22318 6020 22370
rect 5964 22316 6020 22318
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 5572 20018 5628 20020
rect 5572 19966 5574 20018
rect 5574 19966 5626 20018
rect 5626 19966 5628 20018
rect 5572 19964 5628 19966
rect 4844 19404 4900 19460
rect 4508 19346 4564 19348
rect 4508 19294 4510 19346
rect 4510 19294 4562 19346
rect 4562 19294 4564 19346
rect 4508 19292 4564 19294
rect 1820 19234 1876 19236
rect 1820 19182 1822 19234
rect 1822 19182 1874 19234
rect 1874 19182 1876 19234
rect 1820 19180 1876 19182
rect 5124 19234 5180 19236
rect 5124 19182 5126 19234
rect 5126 19182 5178 19234
rect 5178 19182 5180 19234
rect 5124 19180 5180 19182
rect 6076 20076 6132 20132
rect 7084 24722 7140 24724
rect 7084 24670 7086 24722
rect 7086 24670 7138 24722
rect 7138 24670 7140 24722
rect 7084 24668 7140 24670
rect 6412 22204 6468 22260
rect 6188 20018 6244 20020
rect 6188 19966 6190 20018
rect 6190 19966 6242 20018
rect 6242 19966 6244 20018
rect 6188 19964 6244 19966
rect 6300 20076 6356 20132
rect 5908 19458 5964 19460
rect 5908 19406 5910 19458
rect 5910 19406 5962 19458
rect 5962 19406 5964 19458
rect 5908 19404 5964 19406
rect 5740 19180 5796 19236
rect 6300 19292 6356 19348
rect 7196 19964 7252 20020
rect 7196 19404 7252 19460
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4508 15314 4564 15316
rect 4508 15262 4510 15314
rect 4510 15262 4562 15314
rect 4562 15262 4564 15314
rect 4508 15260 4564 15262
rect 6692 19234 6748 19236
rect 6692 19182 6694 19234
rect 6694 19182 6746 19234
rect 6746 19182 6748 19234
rect 6692 19180 6748 19182
rect 6412 18956 6468 19012
rect 6972 18956 7028 19012
rect 7756 28700 7812 28756
rect 7980 28588 8036 28644
rect 8092 28812 8148 28868
rect 8204 28252 8260 28308
rect 7980 24556 8036 24612
rect 9436 30210 9492 30212
rect 9436 30158 9438 30210
rect 9438 30158 9490 30210
rect 9490 30158 9492 30210
rect 9436 30156 9492 30158
rect 12012 34188 12068 34244
rect 16380 37100 16436 37156
rect 13916 35698 13972 35700
rect 13916 35646 13918 35698
rect 13918 35646 13970 35698
rect 13970 35646 13972 35698
rect 13916 35644 13972 35646
rect 14364 35698 14420 35700
rect 14364 35646 14366 35698
rect 14366 35646 14418 35698
rect 14418 35646 14420 35698
rect 14364 35644 14420 35646
rect 16380 35644 16436 35700
rect 13468 35532 13524 35588
rect 16044 35532 16100 35588
rect 14700 35308 14756 35364
rect 13860 34242 13916 34244
rect 13860 34190 13862 34242
rect 13862 34190 13914 34242
rect 13914 34190 13916 34242
rect 13860 34188 13916 34190
rect 14383 34412 14439 34468
rect 15260 34914 15316 34916
rect 15260 34862 15262 34914
rect 15262 34862 15314 34914
rect 15314 34862 15316 34914
rect 15260 34860 15316 34862
rect 14700 34524 14756 34580
rect 10108 30940 10164 30996
rect 9992 30716 10048 30772
rect 10668 30994 10724 30996
rect 10668 30942 10670 30994
rect 10670 30942 10722 30994
rect 10722 30942 10724 30994
rect 10668 30940 10724 30942
rect 10780 29426 10836 29428
rect 10780 29374 10782 29426
rect 10782 29374 10834 29426
rect 10834 29374 10836 29426
rect 10780 29372 10836 29374
rect 9324 28028 9380 28084
rect 10332 28252 10388 28308
rect 9996 26236 10052 26292
rect 9324 24892 9380 24948
rect 10892 28028 10948 28084
rect 11676 31164 11732 31220
rect 11676 30994 11732 30996
rect 11676 30942 11678 30994
rect 11678 30942 11730 30994
rect 11730 30942 11732 30994
rect 11676 30940 11732 30942
rect 12572 31778 12628 31780
rect 12572 31726 12574 31778
rect 12574 31726 12626 31778
rect 12626 31726 12628 31778
rect 12572 31724 12628 31726
rect 13804 31612 13860 31668
rect 12236 30716 12292 30772
rect 11676 30182 11732 30212
rect 11676 30156 11678 30182
rect 11678 30156 11730 30182
rect 11730 30156 11732 30182
rect 11564 29426 11620 29428
rect 11564 29374 11566 29426
rect 11566 29374 11618 29426
rect 11618 29374 11620 29426
rect 11564 29372 11620 29374
rect 12460 30044 12516 30100
rect 12852 30210 12908 30212
rect 12852 30158 12854 30210
rect 12854 30158 12906 30210
rect 12906 30158 12908 30210
rect 12852 30156 12908 30158
rect 13804 30156 13860 30212
rect 16268 34860 16324 34916
rect 16604 35532 16660 35588
rect 18060 37154 18116 37156
rect 18060 37102 18062 37154
rect 18062 37102 18114 37154
rect 18114 37102 18116 37154
rect 18060 37100 18116 37102
rect 17388 35532 17444 35588
rect 16940 34748 16996 34804
rect 14140 29820 14196 29876
rect 12572 28588 12628 28644
rect 13468 28924 13524 28980
rect 10668 25730 10724 25732
rect 10668 25678 10670 25730
rect 10670 25678 10722 25730
rect 10722 25678 10724 25730
rect 10668 25676 10724 25678
rect 10000 25468 10056 25508
rect 10000 25452 10002 25468
rect 10002 25452 10054 25468
rect 10054 25452 10056 25468
rect 9548 24668 9604 24724
rect 8988 23996 9044 24052
rect 10108 23938 10164 23940
rect 10108 23886 10110 23938
rect 10110 23886 10162 23938
rect 10162 23886 10164 23938
rect 10108 23884 10164 23886
rect 10332 25506 10388 25508
rect 10332 25454 10334 25506
rect 10334 25454 10386 25506
rect 10386 25454 10388 25506
rect 10332 25452 10388 25454
rect 11900 25116 11956 25172
rect 14140 28924 14196 28980
rect 15036 32396 15092 32452
rect 13692 28588 13748 28644
rect 13916 27746 13972 27748
rect 13916 27694 13918 27746
rect 13918 27694 13970 27746
rect 13970 27694 13972 27746
rect 13916 27692 13972 27694
rect 13916 26253 13918 26292
rect 13918 26253 13970 26292
rect 13970 26253 13972 26292
rect 13916 26236 13972 26253
rect 14812 31724 14868 31780
rect 14924 29260 14980 29316
rect 14364 27074 14420 27076
rect 14364 27022 14366 27074
rect 14366 27022 14418 27074
rect 14418 27022 14420 27074
rect 14364 27020 14420 27022
rect 14700 26908 14756 26964
rect 14924 25788 14980 25844
rect 14680 25506 14736 25508
rect 14680 25454 14682 25506
rect 14682 25454 14734 25506
rect 14734 25454 14736 25506
rect 14680 25452 14736 25454
rect 14476 25228 14532 25284
rect 13804 25116 13860 25172
rect 15484 31724 15540 31780
rect 15148 30044 15204 30100
rect 15372 30044 15428 30100
rect 16772 34130 16828 34132
rect 16772 34078 16774 34130
rect 16774 34078 16826 34130
rect 16826 34078 16828 34130
rect 16772 34076 16828 34078
rect 17276 34914 17332 34916
rect 17276 34862 17278 34914
rect 17278 34862 17330 34914
rect 17330 34862 17332 34914
rect 17276 34860 17332 34862
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 25396 40402 25452 40404
rect 25396 40350 25398 40402
rect 25398 40350 25450 40402
rect 25450 40350 25452 40402
rect 25396 40348 25452 40350
rect 26012 40402 26068 40404
rect 26012 40350 26014 40402
rect 26014 40350 26066 40402
rect 26066 40350 26068 40402
rect 26012 40348 26068 40350
rect 28588 40348 28644 40404
rect 22652 39788 22708 39844
rect 24444 39842 24500 39844
rect 24444 39790 24446 39842
rect 24446 39790 24498 39842
rect 24498 39790 24500 39842
rect 24444 39788 24500 39790
rect 23660 39676 23716 39732
rect 23436 39564 23492 39620
rect 23548 38780 23604 38836
rect 24332 38834 24388 38836
rect 24332 38782 24334 38834
rect 24334 38782 24386 38834
rect 24386 38782 24388 38834
rect 24332 38780 24388 38782
rect 24444 38220 24500 38276
rect 23660 37884 23716 37940
rect 23996 37884 24052 37940
rect 23830 37772 23886 37828
rect 17612 34412 17668 34468
rect 18004 34636 18060 34692
rect 17836 34130 17892 34132
rect 17836 34078 17838 34130
rect 17838 34078 17890 34130
rect 17890 34078 17892 34130
rect 17836 34076 17892 34078
rect 20524 36988 20580 37044
rect 19516 36876 19572 36932
rect 18396 35698 18452 35700
rect 18396 35646 18398 35698
rect 18398 35646 18450 35698
rect 18450 35646 18452 35698
rect 18396 35644 18452 35646
rect 18284 34300 18340 34356
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 18396 34860 18452 34916
rect 18172 33740 18228 33796
rect 16156 31500 16212 31556
rect 16380 31778 16436 31780
rect 16380 31726 16382 31778
rect 16382 31726 16434 31778
rect 16434 31726 16436 31778
rect 16380 31724 16436 31726
rect 16660 31724 16716 31780
rect 17164 31778 17220 31780
rect 17164 31726 17166 31778
rect 17166 31726 17218 31778
rect 17218 31726 17220 31778
rect 17164 31724 17220 31726
rect 16268 31612 16324 31668
rect 16716 31500 16772 31556
rect 16044 30940 16100 30996
rect 16268 30994 16324 30996
rect 16268 30942 16270 30994
rect 16270 30942 16322 30994
rect 16322 30942 16324 30994
rect 16268 30940 16324 30942
rect 16156 30828 16212 30884
rect 16604 30716 16660 30772
rect 16380 30268 16436 30324
rect 17500 31554 17556 31556
rect 17500 31502 17502 31554
rect 17502 31502 17554 31554
rect 17554 31502 17556 31554
rect 17500 31500 17556 31502
rect 18060 33404 18116 33460
rect 18396 34130 18452 34132
rect 18396 34078 18398 34130
rect 18398 34078 18450 34130
rect 18450 34078 18452 34130
rect 18396 34076 18452 34078
rect 18396 33740 18452 33796
rect 18676 34636 18732 34692
rect 18620 34412 18676 34468
rect 23660 34860 23716 34916
rect 18956 34524 19012 34580
rect 19292 34524 19348 34580
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 18620 33740 18676 33796
rect 19628 34130 19684 34132
rect 19628 34078 19630 34130
rect 19630 34078 19682 34130
rect 19682 34078 19684 34130
rect 19628 34076 19684 34078
rect 19404 33740 19460 33796
rect 21252 34018 21308 34020
rect 21252 33966 21254 34018
rect 21254 33966 21306 34018
rect 21306 33966 21308 34018
rect 21252 33964 21308 33966
rect 21980 33964 22036 34020
rect 22316 33964 22372 34020
rect 23044 34018 23100 34020
rect 23044 33966 23046 34018
rect 23046 33966 23098 34018
rect 23098 33966 23100 34018
rect 23044 33964 23100 33966
rect 20244 33404 20300 33460
rect 18060 31500 18116 31556
rect 17948 30994 18004 30996
rect 17948 30942 17950 30994
rect 17950 30942 18002 30994
rect 18002 30942 18004 30994
rect 17948 30940 18004 30942
rect 15260 29426 15316 29428
rect 15260 29374 15262 29426
rect 15262 29374 15314 29426
rect 15314 29374 15316 29426
rect 15260 29372 15316 29374
rect 15260 26908 15316 26964
rect 15148 25452 15204 25508
rect 14588 24780 14644 24836
rect 14476 24698 14478 24724
rect 14478 24698 14530 24724
rect 14530 24698 14532 24724
rect 14476 24668 14532 24698
rect 14700 24668 14756 24724
rect 14588 24556 14644 24612
rect 10220 22540 10276 22596
rect 13748 23884 13804 23940
rect 13580 22540 13636 22596
rect 7980 22370 8036 22372
rect 7980 22318 7982 22370
rect 7982 22318 8034 22370
rect 8034 22318 8036 22370
rect 7980 22316 8036 22318
rect 10015 21756 10071 21812
rect 12012 22428 12068 22484
rect 11284 22370 11340 22372
rect 11284 22318 11286 22370
rect 11286 22318 11338 22370
rect 11338 22318 11340 22370
rect 11284 22316 11340 22318
rect 13692 22428 13748 22484
rect 11900 21572 11902 21588
rect 11902 21572 11954 21588
rect 11954 21572 11956 21588
rect 13916 21980 13972 22036
rect 12516 21586 12572 21588
rect 11900 21532 11956 21572
rect 12516 21534 12518 21586
rect 12518 21534 12570 21586
rect 12570 21534 12572 21586
rect 12516 21532 12572 21534
rect 9772 20748 9828 20804
rect 9772 20524 9828 20580
rect 9436 19234 9492 19236
rect 9436 19182 9438 19234
rect 9438 19182 9490 19234
rect 9490 19182 9492 19234
rect 9436 19180 9492 19182
rect 11004 20412 11060 20468
rect 11564 20802 11620 20804
rect 11564 20750 11566 20802
rect 11566 20750 11618 20802
rect 11618 20750 11620 20802
rect 11564 20748 11620 20750
rect 11340 20524 11396 20580
rect 12012 20748 12068 20804
rect 13468 20802 13524 20804
rect 13468 20750 13470 20802
rect 13470 20750 13522 20802
rect 13522 20750 13524 20802
rect 13468 20748 13524 20750
rect 11900 20412 11956 20468
rect 12124 20076 12180 20132
rect 11004 19458 11060 19460
rect 11004 19406 11006 19458
rect 11006 19406 11058 19458
rect 11058 19406 11060 19458
rect 11004 19404 11060 19406
rect 12628 20130 12684 20132
rect 12628 20078 12630 20130
rect 12630 20078 12682 20130
rect 12682 20078 12684 20130
rect 12628 20076 12684 20078
rect 10108 18508 10164 18564
rect 10388 18562 10444 18564
rect 10388 18510 10390 18562
rect 10390 18510 10442 18562
rect 10442 18510 10444 18562
rect 10388 18508 10444 18510
rect 7644 18284 7700 18340
rect 5068 15260 5124 15316
rect 5516 15260 5572 15316
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5292 14588 5348 14644
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4956 12684 5012 12740
rect 7812 15314 7868 15316
rect 7812 15262 7814 15314
rect 7814 15262 7866 15314
rect 7866 15262 7868 15314
rect 7812 15260 7868 15262
rect 9436 15314 9492 15316
rect 9436 15262 9438 15314
rect 9438 15262 9490 15314
rect 9490 15262 9492 15314
rect 9436 15260 9492 15262
rect 5852 14642 5908 14644
rect 5852 14590 5854 14642
rect 5854 14590 5906 14642
rect 5906 14590 5908 14642
rect 5852 14588 5908 14590
rect 5964 14515 6020 14532
rect 5964 14476 5966 14515
rect 5966 14476 6018 14515
rect 6018 14476 6020 14515
rect 2268 12178 2324 12180
rect 2268 12126 2270 12178
rect 2270 12126 2322 12178
rect 2322 12126 2324 12178
rect 2268 12124 2324 12126
rect 5516 12124 5572 12180
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 3052 11564 3108 11620
rect 3724 11618 3780 11620
rect 3724 11566 3726 11618
rect 3726 11566 3778 11618
rect 3778 11566 3780 11618
rect 3724 11564 3780 11566
rect 4060 11394 4116 11396
rect 4060 11342 4062 11394
rect 4062 11342 4114 11394
rect 4114 11342 4116 11394
rect 4060 11340 4116 11342
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4956 9938 5012 9940
rect 4956 9886 4958 9938
rect 4958 9886 5010 9938
rect 5010 9886 5012 9938
rect 4956 9884 5012 9886
rect 6748 14530 6804 14532
rect 6748 14478 6750 14530
rect 6750 14478 6802 14530
rect 6802 14478 6804 14530
rect 6748 14476 6804 14478
rect 10332 15148 10388 15204
rect 10444 15260 10500 15316
rect 11004 15260 11060 15316
rect 12964 15202 13020 15204
rect 12964 15150 12966 15202
rect 12966 15150 13018 15202
rect 13018 15150 13020 15202
rect 12964 15148 13020 15150
rect 12460 14530 12516 14532
rect 6972 13132 7028 13188
rect 7644 13132 7700 13188
rect 7420 12962 7476 12964
rect 7420 12910 7422 12962
rect 7422 12910 7474 12962
rect 7474 12910 7476 12962
rect 7420 12908 7476 12910
rect 12460 14478 12462 14530
rect 12462 14478 12514 14530
rect 12514 14478 12516 14530
rect 12460 14476 12516 14478
rect 12908 14476 12964 14532
rect 12124 13916 12180 13972
rect 8652 13020 8708 13076
rect 7868 12908 7924 12964
rect 7028 12684 7084 12740
rect 6860 11340 6916 11396
rect 8540 12962 8596 12964
rect 8540 12910 8542 12962
rect 8542 12910 8594 12962
rect 8594 12910 8596 12962
rect 8540 12908 8596 12910
rect 8204 12796 8260 12852
rect 9324 12947 9380 12964
rect 9324 12908 9326 12947
rect 9326 12908 9378 12947
rect 9378 12908 9380 12947
rect 8988 12796 9044 12852
rect 7644 12684 7700 12740
rect 11340 13468 11396 13524
rect 12236 13020 12292 13076
rect 11564 12684 11620 12740
rect 12572 13804 12628 13860
rect 12796 13356 12852 13412
rect 12348 12684 12404 12740
rect 9436 12124 9492 12180
rect 12236 11452 12292 11508
rect 6748 10332 6804 10388
rect 3052 9212 3108 9268
rect 4172 9266 4228 9268
rect 4172 9214 4174 9266
rect 4174 9214 4226 9266
rect 4226 9214 4228 9266
rect 4172 9212 4228 9214
rect 4508 9042 4564 9044
rect 4508 8990 4510 9042
rect 4510 8990 4562 9042
rect 4562 8990 4564 9042
rect 4508 8988 4564 8990
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 9660 10386 9716 10388
rect 9660 10334 9662 10386
rect 9662 10334 9714 10386
rect 9714 10334 9716 10386
rect 9660 10332 9716 10334
rect 10444 10108 10500 10164
rect 7420 9996 7476 10052
rect 7980 9996 8036 10052
rect 7084 9884 7140 9940
rect 7420 9826 7476 9828
rect 7420 9774 7422 9826
rect 7422 9774 7474 9826
rect 7474 9774 7476 9826
rect 7420 9772 7476 9774
rect 7308 8988 7364 9044
rect 8988 9996 9044 10052
rect 8204 9826 8260 9828
rect 8204 9774 8206 9826
rect 8206 9774 8258 9826
rect 8258 9774 8260 9826
rect 8204 9772 8260 9774
rect 7868 9660 7924 9716
rect 8708 9714 8764 9716
rect 8708 9662 8710 9714
rect 8710 9662 8762 9714
rect 8762 9662 8764 9714
rect 8708 9660 8764 9662
rect 9100 9826 9156 9828
rect 9100 9774 9102 9826
rect 9102 9774 9154 9826
rect 9154 9774 9156 9826
rect 9100 9772 9156 9774
rect 8988 9324 9044 9380
rect 9772 9660 9828 9716
rect 10108 9042 10164 9044
rect 10108 8990 10110 9042
rect 10110 8990 10162 9042
rect 10162 8990 10164 9042
rect 10108 8988 10164 8990
rect 11508 10108 11564 10164
rect 10780 9772 10836 9828
rect 10612 9042 10668 9044
rect 10612 8990 10614 9042
rect 10614 8990 10666 9042
rect 10666 8990 10668 9042
rect 10612 8988 10668 8990
rect 10780 8988 10836 9044
rect 10892 9324 10948 9380
rect 11788 9212 11844 9268
rect 12124 9042 12180 9044
rect 12124 8990 12126 9042
rect 12126 8990 12178 9042
rect 12178 8990 12180 9042
rect 12124 8988 12180 8990
rect 7644 7532 7700 7588
rect 13132 13746 13188 13748
rect 13132 13694 13134 13746
rect 13134 13694 13186 13746
rect 13186 13694 13188 13746
rect 13132 13692 13188 13694
rect 15036 24668 15092 24724
rect 16492 29932 16548 29988
rect 16716 29372 16772 29428
rect 16828 30716 16884 30772
rect 16212 29314 16268 29316
rect 16212 29262 16214 29314
rect 16214 29262 16266 29314
rect 16266 29262 16268 29314
rect 16212 29260 16268 29262
rect 16716 27692 16772 27748
rect 15260 24668 15316 24724
rect 16604 25116 16660 25172
rect 15092 24050 15148 24052
rect 15092 23998 15094 24050
rect 15094 23998 15146 24050
rect 15146 23998 15148 24050
rect 15092 23996 15148 23998
rect 15260 23548 15316 23604
rect 14588 18508 14644 18564
rect 15596 23714 15652 23716
rect 15596 23662 15598 23714
rect 15598 23662 15650 23714
rect 15650 23662 15652 23714
rect 15596 23660 15652 23662
rect 15876 23548 15932 23604
rect 15036 22428 15092 22484
rect 14924 22370 14980 22372
rect 14924 22318 14926 22370
rect 14926 22318 14978 22370
rect 14978 22318 14980 22370
rect 14924 22316 14980 22318
rect 14812 22204 14868 22260
rect 14700 18450 14756 18452
rect 14700 18398 14702 18450
rect 14702 18398 14754 18450
rect 14754 18398 14756 18450
rect 14700 18396 14756 18398
rect 15316 22316 15372 22372
rect 15202 22092 15258 22148
rect 16716 22428 16772 22484
rect 16100 22258 16156 22260
rect 16100 22206 16102 22258
rect 16102 22206 16154 22258
rect 16154 22206 16156 22258
rect 16100 22204 16156 22206
rect 16604 22092 16660 22148
rect 15484 21644 15540 21700
rect 15932 21868 15988 21924
rect 16156 21644 16212 21700
rect 17556 30716 17612 30772
rect 17108 30268 17164 30324
rect 16940 30098 16996 30100
rect 16940 30046 16942 30098
rect 16942 30046 16994 30098
rect 16994 30046 16996 30098
rect 16940 30044 16996 30046
rect 17556 30098 17612 30100
rect 17556 30046 17558 30098
rect 17558 30046 17610 30098
rect 17610 30046 17612 30098
rect 17556 30044 17612 30046
rect 17388 28476 17444 28532
rect 17500 27916 17556 27972
rect 17836 28028 17892 28084
rect 17388 23660 17444 23716
rect 17836 26236 17892 26292
rect 16716 21868 16772 21924
rect 16828 21586 16884 21588
rect 16828 21534 16830 21586
rect 16830 21534 16882 21586
rect 16882 21534 16884 21586
rect 16828 21532 16884 21534
rect 15204 18450 15260 18452
rect 15204 18398 15206 18450
rect 15206 18398 15258 18450
rect 15258 18398 15260 18450
rect 15204 18396 15260 18398
rect 14084 18338 14140 18340
rect 14084 18286 14086 18338
rect 14086 18286 14138 18338
rect 14138 18286 14140 18338
rect 14084 18284 14140 18286
rect 15036 18284 15092 18340
rect 14196 17612 14252 17668
rect 14476 17724 14532 17780
rect 14140 14812 14196 14868
rect 13468 13356 13524 13412
rect 13580 14476 13636 14532
rect 13692 13804 13748 13860
rect 14700 17666 14756 17668
rect 14700 17614 14702 17666
rect 14702 17614 14754 17666
rect 14754 17614 14756 17666
rect 14700 17612 14756 17614
rect 16324 18956 16380 19012
rect 15596 18396 15652 18452
rect 15764 18284 15820 18340
rect 15372 17778 15428 17780
rect 15372 17726 15374 17778
rect 15374 17726 15426 17778
rect 15426 17726 15428 17778
rect 15372 17724 15428 17726
rect 15260 17612 15316 17668
rect 16604 18450 16660 18452
rect 16604 18398 16606 18450
rect 16606 18398 16658 18450
rect 16658 18398 16660 18450
rect 16604 18396 16660 18398
rect 16716 18284 16772 18340
rect 17724 22370 17780 22372
rect 17724 22318 17726 22370
rect 17726 22318 17778 22370
rect 17778 22318 17780 22370
rect 17724 22316 17780 22318
rect 17556 22258 17612 22260
rect 17556 22206 17558 22258
rect 17558 22206 17610 22258
rect 17610 22206 17612 22258
rect 17556 22204 17612 22206
rect 18060 27858 18116 27860
rect 18060 27806 18062 27858
rect 18062 27806 18114 27858
rect 18114 27806 18116 27858
rect 18060 27804 18116 27806
rect 18450 33346 18506 33348
rect 18450 33294 18452 33346
rect 18452 33294 18504 33346
rect 18504 33294 18506 33346
rect 18450 33292 18506 33294
rect 19292 33292 19348 33348
rect 18284 30940 18340 30996
rect 18396 33068 18452 33124
rect 18844 31500 18900 31556
rect 19180 30994 19236 30996
rect 19180 30942 19182 30994
rect 19182 30942 19234 30994
rect 19234 30942 19236 30994
rect 19180 30940 19236 30942
rect 18732 30268 18788 30324
rect 18284 30044 18340 30100
rect 18284 28700 18340 28756
rect 19068 28476 19124 28532
rect 18788 28082 18844 28084
rect 18788 28030 18790 28082
rect 18790 28030 18842 28082
rect 18842 28030 18844 28082
rect 18788 28028 18844 28030
rect 19460 33346 19516 33348
rect 19460 33294 19462 33346
rect 19462 33294 19514 33346
rect 19514 33294 19516 33346
rect 19460 33292 19516 33294
rect 22484 33906 22540 33908
rect 22484 33854 22486 33906
rect 22486 33854 22538 33906
rect 22538 33854 22540 33906
rect 22484 33852 22540 33854
rect 23324 33852 23380 33908
rect 21644 33516 21700 33572
rect 22596 33516 22652 33572
rect 23660 33516 23716 33572
rect 25004 37772 25060 37828
rect 26348 37324 26404 37380
rect 25900 37250 25902 37268
rect 25902 37250 25954 37268
rect 25954 37250 25956 37268
rect 28028 37996 28084 38052
rect 27804 37324 27860 37380
rect 25900 37212 25956 37250
rect 25564 37100 25620 37156
rect 21532 33068 21588 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 21196 32060 21252 32116
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20076 30940 20132 30996
rect 19964 30044 20020 30100
rect 20412 30044 20468 30100
rect 21084 30044 21140 30100
rect 20188 29932 20244 29988
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19516 29372 19572 29428
rect 20860 29426 20916 29428
rect 20860 29374 20862 29426
rect 20862 29374 20914 29426
rect 20914 29374 20916 29426
rect 20860 29372 20916 29374
rect 20188 28812 20244 28868
rect 20636 28866 20692 28868
rect 20636 28814 20638 28866
rect 20638 28814 20690 28866
rect 20690 28814 20692 28866
rect 20636 28812 20692 28814
rect 19292 28028 19348 28084
rect 20412 28588 20468 28644
rect 18620 27804 18676 27860
rect 18508 26908 18564 26964
rect 18228 26402 18284 26404
rect 18228 26350 18230 26402
rect 18230 26350 18282 26402
rect 18282 26350 18284 26402
rect 18228 26348 18284 26350
rect 18508 26290 18564 26292
rect 18508 26238 18510 26290
rect 18510 26238 18562 26290
rect 18562 26238 18564 26290
rect 18508 26236 18564 26238
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19404 27692 19460 27748
rect 18900 27580 18956 27636
rect 18900 26962 18956 26964
rect 18900 26910 18902 26962
rect 18902 26910 18954 26962
rect 18954 26910 18956 26962
rect 18900 26908 18956 26910
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19124 26348 19180 26404
rect 18172 25676 18228 25732
rect 17948 25116 18004 25172
rect 18396 25116 18452 25172
rect 19068 26124 19124 26180
rect 18844 26012 18900 26068
rect 18060 22540 18116 22596
rect 17948 22428 18004 22484
rect 18228 22258 18284 22260
rect 18228 22206 18230 22258
rect 18230 22206 18282 22258
rect 18282 22206 18284 22258
rect 18228 22204 18284 22206
rect 18620 22540 18676 22596
rect 18396 21980 18452 22036
rect 17780 19234 17836 19236
rect 17780 19182 17782 19234
rect 17782 19182 17834 19234
rect 17834 19182 17836 19234
rect 17780 19180 17836 19182
rect 17388 18284 17444 18340
rect 16940 16044 16996 16100
rect 18956 22482 19012 22484
rect 18956 22430 18958 22482
rect 18958 22430 19010 22482
rect 19010 22430 19012 22482
rect 18956 22428 19012 22430
rect 18956 21980 19012 22036
rect 19180 25676 19236 25732
rect 19292 25452 19348 25508
rect 19180 25228 19236 25284
rect 19684 26066 19740 26068
rect 19684 26014 19686 26066
rect 19686 26014 19738 26066
rect 19738 26014 19740 26066
rect 19684 26012 19740 26014
rect 19628 25340 19684 25396
rect 20300 25340 20356 25396
rect 19628 25116 19684 25172
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20188 24892 20244 24948
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20076 22540 20132 22596
rect 19460 22204 19516 22260
rect 19628 22204 19684 22260
rect 20412 22428 20468 22484
rect 20076 22204 20132 22260
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19292 21532 19348 21588
rect 20972 21644 21028 21700
rect 20300 21586 20356 21588
rect 20300 21534 20302 21586
rect 20302 21534 20354 21586
rect 20354 21534 20356 21586
rect 20300 21532 20356 21534
rect 19068 21420 19124 21476
rect 19796 21474 19852 21476
rect 19796 21422 19798 21474
rect 19798 21422 19850 21474
rect 19850 21422 19852 21474
rect 19796 21420 19852 21422
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19964 18284 20020 18340
rect 20188 18172 20244 18228
rect 17836 17836 17892 17892
rect 20860 19234 20916 19236
rect 20860 19182 20862 19234
rect 20862 19182 20914 19234
rect 20914 19182 20916 19234
rect 20860 19180 20916 19182
rect 20748 17836 20804 17892
rect 20860 18732 20916 18788
rect 20748 17612 20804 17668
rect 17724 17442 17780 17444
rect 17724 17390 17726 17442
rect 17726 17390 17778 17442
rect 17778 17390 17780 17442
rect 17724 17388 17780 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 21084 18732 21140 18788
rect 20972 18226 21028 18228
rect 20972 18174 20974 18226
rect 20974 18174 21026 18226
rect 21026 18174 21028 18226
rect 20972 18172 21028 18174
rect 20860 17388 20916 17444
rect 20748 16882 20804 16884
rect 20748 16830 20750 16882
rect 20750 16830 20802 16882
rect 20802 16830 20804 16882
rect 20748 16828 20804 16830
rect 21868 31836 21924 31892
rect 21980 31948 22036 32004
rect 21532 30716 21588 30772
rect 21476 30098 21532 30100
rect 21476 30046 21478 30098
rect 21478 30046 21530 30098
rect 21530 30046 21532 30098
rect 21476 30044 21532 30046
rect 23660 33346 23716 33348
rect 23660 33294 23662 33346
rect 23662 33294 23714 33346
rect 23714 33294 23716 33346
rect 23660 33292 23716 33294
rect 23268 33122 23324 33124
rect 23268 33070 23270 33122
rect 23270 33070 23322 33122
rect 23322 33070 23324 33122
rect 23268 33068 23324 33070
rect 22652 32620 22708 32676
rect 24836 34914 24892 34916
rect 24836 34862 24838 34914
rect 24838 34862 24890 34914
rect 24890 34862 24892 34914
rect 24836 34860 24892 34862
rect 25620 34914 25676 34916
rect 25620 34862 25622 34914
rect 25622 34862 25674 34914
rect 25674 34862 25676 34914
rect 25620 34860 25676 34862
rect 25788 34636 25844 34692
rect 27580 37266 27636 37268
rect 27580 37214 27582 37266
rect 27582 37214 27634 37266
rect 27634 37214 27636 37266
rect 27580 37212 27636 37214
rect 26504 37100 26560 37156
rect 25900 34914 25956 34916
rect 25900 34862 25902 34914
rect 25902 34862 25954 34914
rect 25954 34862 25956 34914
rect 25900 34860 25956 34862
rect 24668 33292 24724 33348
rect 24556 32620 24612 32676
rect 22428 32060 22484 32116
rect 23324 32060 23380 32116
rect 26852 35196 26908 35252
rect 27356 34914 27412 34916
rect 27356 34862 27358 34914
rect 27358 34862 27410 34914
rect 27410 34862 27412 34914
rect 27356 34860 27412 34862
rect 28364 37996 28420 38052
rect 28364 35308 28420 35364
rect 28028 34860 28084 34916
rect 27804 34636 27860 34692
rect 28252 34300 28308 34356
rect 28476 34748 28532 34804
rect 27300 33516 27356 33572
rect 24556 31724 24612 31780
rect 24668 31836 24724 31892
rect 21980 30044 22036 30100
rect 22428 30156 22484 30212
rect 21420 29202 21476 29204
rect 21420 29150 21422 29202
rect 21422 29150 21474 29202
rect 21474 29150 21476 29202
rect 21420 29148 21476 29150
rect 21756 27074 21812 27076
rect 21756 27022 21758 27074
rect 21758 27022 21810 27074
rect 21810 27022 21812 27074
rect 21756 27020 21812 27022
rect 21420 26236 21476 26292
rect 21420 25340 21476 25396
rect 21868 24668 21924 24724
rect 21364 23266 21420 23268
rect 21364 23214 21366 23266
rect 21366 23214 21418 23266
rect 21418 23214 21420 23266
rect 21364 23212 21420 23214
rect 21644 23212 21700 23268
rect 24108 29932 24164 29988
rect 22652 27916 22708 27972
rect 22764 28700 22820 28756
rect 22540 26290 22596 26292
rect 22540 26238 22542 26290
rect 22542 26238 22594 26290
rect 22594 26238 22596 26290
rect 22540 26236 22596 26238
rect 22540 25452 22596 25508
rect 22988 25506 23044 25508
rect 22988 25454 22990 25506
rect 22990 25454 23042 25506
rect 23042 25454 23044 25506
rect 22988 25452 23044 25454
rect 27132 33292 27188 33348
rect 25340 31836 25396 31892
rect 25228 27804 25284 27860
rect 24724 27746 24780 27748
rect 24724 27694 24726 27746
rect 24726 27694 24778 27746
rect 24778 27694 24780 27746
rect 24724 27692 24780 27694
rect 25004 27692 25060 27748
rect 25564 27858 25620 27860
rect 25564 27806 25566 27858
rect 25566 27806 25618 27858
rect 25618 27806 25620 27858
rect 25564 27804 25620 27806
rect 25788 31778 25844 31780
rect 25788 31726 25790 31778
rect 25790 31726 25842 31778
rect 25842 31726 25844 31778
rect 25788 31724 25844 31726
rect 27748 31890 27804 31892
rect 27748 31838 27750 31890
rect 27750 31838 27802 31890
rect 27802 31838 27804 31890
rect 27748 31836 27804 31838
rect 28476 33516 28532 33572
rect 28476 31948 28532 32004
rect 29316 40402 29372 40404
rect 29316 40350 29318 40402
rect 29318 40350 29370 40402
rect 29370 40350 29372 40402
rect 29316 40348 29372 40350
rect 29708 40402 29764 40404
rect 29708 40350 29710 40402
rect 29710 40350 29762 40402
rect 29762 40350 29764 40402
rect 29708 40348 29764 40350
rect 36092 40460 36148 40516
rect 32788 40348 32844 40404
rect 33292 40402 33348 40404
rect 33292 40350 33294 40402
rect 33294 40350 33346 40402
rect 33346 40350 33348 40402
rect 33292 40348 33348 40350
rect 32844 39842 32900 39844
rect 32844 39790 32846 39842
rect 32846 39790 32898 39842
rect 32898 39790 32900 39842
rect 32844 39788 32900 39790
rect 39676 40626 39732 40628
rect 39676 40574 39678 40626
rect 39678 40574 39730 40626
rect 39730 40574 39732 40626
rect 39676 40572 39732 40574
rect 41132 41858 41188 41860
rect 41132 41806 41134 41858
rect 41134 41806 41186 41858
rect 41186 41806 41188 41858
rect 41132 41804 41188 41806
rect 40124 40572 40180 40628
rect 39004 40514 39060 40516
rect 39004 40462 39006 40514
rect 39006 40462 39058 40514
rect 39058 40462 39060 40514
rect 39004 40460 39060 40462
rect 39340 40460 39396 40516
rect 36372 40402 36428 40404
rect 36372 40350 36374 40402
rect 36374 40350 36426 40402
rect 36426 40350 36428 40402
rect 36372 40348 36428 40350
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34076 39788 34132 39844
rect 29148 39452 29204 39508
rect 28924 38780 28980 38836
rect 28700 37772 28756 37828
rect 28700 37100 28756 37156
rect 29036 38050 29092 38052
rect 29036 37998 29038 38050
rect 29038 37998 29090 38050
rect 29090 37998 29092 38050
rect 29036 37996 29092 37998
rect 29260 38780 29316 38836
rect 29540 37938 29596 37940
rect 29540 37886 29542 37938
rect 29542 37886 29594 37938
rect 29594 37886 29596 37938
rect 29540 37884 29596 37886
rect 28958 35308 29014 35364
rect 28812 35196 28868 35252
rect 29372 37324 29428 37380
rect 29596 35196 29652 35252
rect 28700 34860 28756 34916
rect 29148 34914 29204 34916
rect 29148 34862 29150 34914
rect 29150 34862 29202 34914
rect 29202 34862 29204 34914
rect 29148 34860 29204 34862
rect 29372 34636 29428 34692
rect 29260 34300 29316 34356
rect 28364 31836 28420 31892
rect 28588 31836 28644 31892
rect 28700 33292 28756 33348
rect 28196 31554 28252 31556
rect 28196 31502 28198 31554
rect 28198 31502 28250 31554
rect 28250 31502 28252 31554
rect 28196 31500 28252 31502
rect 27132 30380 27188 30436
rect 26908 30044 26964 30100
rect 27580 30994 27636 30996
rect 27580 30942 27582 30994
rect 27582 30942 27634 30994
rect 27634 30942 27636 30994
rect 27580 30940 27636 30942
rect 26684 29932 26740 29988
rect 25900 27692 25956 27748
rect 28700 30940 28756 30996
rect 29148 31500 29204 31556
rect 28476 30380 28532 30436
rect 29148 30268 29204 30324
rect 28140 30044 28196 30100
rect 27020 28642 27076 28644
rect 27020 28590 27022 28642
rect 27022 28590 27074 28642
rect 27074 28590 27076 28642
rect 27020 28588 27076 28590
rect 26572 27858 26628 27860
rect 26572 27806 26574 27858
rect 26574 27806 26626 27858
rect 26626 27806 26628 27858
rect 26572 27804 26628 27806
rect 29484 33346 29540 33348
rect 29484 33294 29486 33346
rect 29486 33294 29538 33346
rect 29538 33294 29540 33346
rect 29484 33292 29540 33294
rect 30156 37826 30212 37828
rect 30156 37774 30158 37826
rect 30158 37774 30210 37826
rect 30210 37774 30212 37826
rect 30156 37772 30212 37774
rect 35812 38722 35868 38724
rect 35812 38670 35814 38722
rect 35814 38670 35866 38722
rect 35866 38670 35868 38722
rect 35812 38668 35868 38670
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 32508 37324 32564 37380
rect 32956 37772 33012 37828
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 29820 34300 29876 34356
rect 30156 34748 30212 34804
rect 33740 36204 33796 36260
rect 34132 36258 34188 36260
rect 34132 36206 34134 36258
rect 34134 36206 34186 36258
rect 34186 36206 34188 36258
rect 34132 36204 34188 36206
rect 29988 33852 30044 33908
rect 30604 33404 30660 33460
rect 32508 33852 32564 33908
rect 29820 33346 29876 33348
rect 29820 33294 29822 33346
rect 29822 33294 29874 33346
rect 29874 33294 29876 33346
rect 29820 33292 29876 33294
rect 31276 33292 31332 33348
rect 32844 31948 32900 32004
rect 30156 31836 30212 31892
rect 31836 31836 31892 31892
rect 33460 31890 33516 31892
rect 33460 31838 33462 31890
rect 33462 31838 33514 31890
rect 33514 31838 33516 31890
rect 33460 31836 33516 31838
rect 32564 31500 32620 31556
rect 33068 31500 33124 31556
rect 36390 38668 36446 38724
rect 39340 39564 39396 39620
rect 41804 39788 41860 39844
rect 42588 39842 42644 39844
rect 42588 39790 42590 39842
rect 42590 39790 42642 39842
rect 42642 39790 42644 39842
rect 42588 39788 42644 39790
rect 36540 36204 36596 36260
rect 37156 36258 37212 36260
rect 37156 36206 37158 36258
rect 37158 36206 37210 36258
rect 37210 36206 37212 36258
rect 37156 36204 37212 36206
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36428 35644 36484 35700
rect 34748 34188 34804 34244
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 34636 31948 34692 32004
rect 34412 31052 34468 31108
rect 31388 28812 31444 28868
rect 28252 27074 28308 27076
rect 28252 27022 28254 27074
rect 28254 27022 28306 27074
rect 28306 27022 28308 27074
rect 28252 27020 28308 27022
rect 29036 27804 29092 27860
rect 26236 26908 26292 26964
rect 28364 26908 28420 26964
rect 24108 25788 24164 25844
rect 28252 26684 28308 26740
rect 25340 25340 25396 25396
rect 25844 25394 25900 25396
rect 25844 25342 25846 25394
rect 25846 25342 25898 25394
rect 25898 25342 25900 25394
rect 25844 25340 25900 25342
rect 24108 25116 24164 25172
rect 23436 24946 23492 24948
rect 23436 24894 23438 24946
rect 23438 24894 23490 24946
rect 23490 24894 23492 24946
rect 23436 24892 23492 24894
rect 23772 24892 23828 24948
rect 22932 24722 22988 24724
rect 22932 24670 22934 24722
rect 22934 24670 22986 24722
rect 22986 24670 22988 24722
rect 22932 24668 22988 24670
rect 22932 23884 22988 23940
rect 23548 23938 23604 23940
rect 23548 23886 23550 23938
rect 23550 23886 23602 23938
rect 23602 23886 23604 23938
rect 23548 23884 23604 23886
rect 25284 24444 25340 24500
rect 23268 23212 23324 23268
rect 23772 23212 23828 23268
rect 21868 20076 21924 20132
rect 21588 18338 21644 18340
rect 21588 18286 21590 18338
rect 21590 18286 21642 18338
rect 21642 18286 21644 18338
rect 21588 18284 21644 18286
rect 21364 17890 21420 17892
rect 21364 17838 21366 17890
rect 21366 17838 21418 17890
rect 21418 17838 21420 17890
rect 21364 17836 21420 17838
rect 21196 17052 21252 17108
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 15708 15484 15764 15540
rect 14700 15148 14756 15204
rect 14700 14588 14756 14644
rect 15036 15148 15092 15204
rect 14476 13804 14532 13860
rect 13860 13580 13916 13636
rect 14028 13692 14084 13748
rect 14700 13746 14756 13748
rect 14700 13694 14702 13746
rect 14702 13694 14754 13746
rect 14754 13694 14756 13746
rect 14700 13692 14756 13694
rect 14364 13580 14420 13636
rect 14252 13522 14308 13524
rect 14252 13470 14254 13522
rect 14254 13470 14306 13522
rect 14306 13470 14308 13522
rect 14252 13468 14308 13470
rect 13244 12178 13300 12180
rect 13244 12126 13246 12178
rect 13246 12126 13298 12178
rect 13298 12126 13300 12178
rect 13244 12124 13300 12126
rect 13580 12178 13636 12180
rect 13580 12126 13582 12178
rect 13582 12126 13634 12178
rect 13634 12126 13636 12178
rect 13580 12124 13636 12126
rect 12908 11452 12964 11508
rect 12348 9324 12404 9380
rect 13132 9884 13188 9940
rect 13468 9884 13524 9940
rect 12460 9212 12516 9268
rect 12348 9100 12404 9156
rect 13300 9100 13356 9156
rect 13580 9212 13636 9268
rect 9660 8204 9716 8260
rect 10668 8258 10724 8260
rect 10668 8206 10670 8258
rect 10670 8206 10722 8258
rect 10722 8206 10724 8258
rect 10668 8204 10724 8206
rect 7756 5906 7812 5908
rect 7756 5854 7758 5906
rect 7758 5854 7810 5906
rect 7810 5854 7812 5906
rect 7756 5852 7812 5854
rect 9604 5852 9660 5908
rect 9212 5740 9268 5796
rect 8428 5628 8484 5684
rect 5852 5068 5908 5124
rect 6524 5122 6580 5124
rect 6524 5070 6526 5122
rect 6526 5070 6578 5122
rect 6578 5070 6580 5122
rect 6524 5068 6580 5070
rect 8932 5682 8988 5684
rect 8932 5630 8934 5682
rect 8934 5630 8986 5682
rect 8986 5630 8988 5682
rect 8932 5628 8988 5630
rect 9772 5906 9828 5908
rect 9772 5854 9774 5906
rect 9774 5854 9826 5906
rect 9826 5854 9828 5906
rect 9772 5852 9828 5854
rect 9828 5234 9884 5236
rect 9828 5182 9830 5234
rect 9830 5182 9882 5234
rect 9882 5182 9884 5234
rect 9828 5180 9884 5182
rect 10108 5180 10164 5236
rect 12572 7532 12628 7588
rect 12012 5906 12068 5908
rect 12012 5854 12014 5906
rect 12014 5854 12066 5906
rect 12066 5854 12068 5906
rect 12012 5852 12068 5854
rect 12460 5893 12462 5908
rect 12462 5893 12514 5908
rect 12514 5893 12516 5908
rect 12460 5852 12516 5893
rect 16716 15202 16772 15204
rect 16716 15150 16718 15202
rect 16718 15150 16770 15202
rect 16770 15150 16772 15202
rect 16716 15148 16772 15150
rect 15372 14812 15428 14868
rect 17500 14812 17556 14868
rect 17332 14642 17388 14644
rect 17332 14590 17334 14642
rect 17334 14590 17386 14642
rect 17386 14590 17388 14642
rect 17332 14588 17388 14590
rect 15652 13970 15708 13972
rect 15652 13918 15654 13970
rect 15654 13918 15706 13970
rect 15706 13918 15708 13970
rect 15652 13916 15708 13918
rect 15652 13468 15708 13524
rect 19628 14252 19684 14308
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21868 17666 21924 17668
rect 21868 17614 21870 17666
rect 21870 17614 21922 17666
rect 21922 17614 21924 17666
rect 21868 17612 21924 17614
rect 22260 17666 22316 17668
rect 22260 17614 22262 17666
rect 22262 17614 22314 17666
rect 22314 17614 22316 17666
rect 22260 17612 22316 17614
rect 21700 17106 21756 17108
rect 21700 17054 21702 17106
rect 21702 17054 21754 17106
rect 21754 17054 21756 17106
rect 21700 17052 21756 17054
rect 22204 17106 22260 17108
rect 22204 17054 22206 17106
rect 22206 17054 22258 17106
rect 22258 17054 22260 17106
rect 22204 17052 22260 17054
rect 21756 16828 21812 16884
rect 21532 16268 21588 16324
rect 20356 14306 20412 14308
rect 20356 14254 20358 14306
rect 20358 14254 20410 14306
rect 20410 14254 20412 14306
rect 20356 14252 20412 14254
rect 20188 13916 20244 13972
rect 20300 13804 20356 13860
rect 20076 13746 20132 13748
rect 20076 13694 20078 13746
rect 20078 13694 20130 13746
rect 20130 13694 20132 13746
rect 20076 13692 20132 13694
rect 21084 13804 21140 13860
rect 20524 13746 20580 13748
rect 20524 13694 20526 13746
rect 20526 13694 20578 13746
rect 20578 13694 20580 13746
rect 20524 13692 20580 13694
rect 21308 13746 21364 13748
rect 21308 13694 21310 13746
rect 21310 13694 21362 13746
rect 21362 13694 21364 13746
rect 21308 13692 21364 13694
rect 21644 13692 21700 13748
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 14812 12124 14868 12180
rect 28588 26012 28644 26068
rect 28924 26290 28980 26292
rect 28924 26238 28926 26290
rect 28926 26238 28978 26290
rect 28978 26238 28980 26290
rect 28924 26236 28980 26238
rect 28924 25676 28980 25732
rect 29932 26908 29988 26964
rect 29708 26796 29764 26852
rect 30268 26684 30324 26740
rect 30492 26908 30548 26964
rect 29596 26236 29652 26292
rect 30360 26124 30416 26180
rect 30156 26012 30212 26068
rect 30604 26796 30660 26852
rect 31220 26178 31276 26180
rect 31220 26126 31222 26178
rect 31222 26126 31274 26178
rect 31274 26126 31276 26178
rect 31220 26124 31276 26126
rect 30716 26012 30772 26068
rect 24556 20802 24612 20804
rect 24556 20750 24558 20802
rect 24558 20750 24610 20802
rect 24610 20750 24612 20802
rect 24556 20748 24612 20750
rect 27356 22204 27412 22260
rect 28364 22204 28420 22260
rect 28232 21756 28288 21812
rect 24948 20748 25004 20804
rect 24444 18284 24500 18340
rect 24444 17724 24500 17780
rect 22652 16156 22708 16212
rect 23884 16268 23940 16324
rect 23044 16098 23100 16100
rect 23044 16046 23046 16098
rect 23046 16046 23098 16098
rect 23098 16046 23100 16098
rect 23044 16044 23100 16046
rect 23548 15314 23604 15316
rect 23548 15262 23550 15314
rect 23550 15262 23602 15314
rect 23602 15262 23604 15314
rect 23548 15260 23604 15262
rect 22652 14588 22708 14644
rect 27804 20130 27860 20132
rect 27804 20078 27806 20130
rect 27806 20078 27858 20130
rect 27858 20078 27860 20130
rect 27804 20076 27860 20078
rect 25116 20018 25172 20020
rect 25116 19966 25118 20018
rect 25118 19966 25170 20018
rect 25170 19966 25172 20018
rect 25116 19964 25172 19966
rect 30584 25506 30640 25508
rect 30584 25454 30586 25506
rect 30586 25454 30638 25506
rect 30638 25454 30640 25506
rect 30584 25452 30640 25454
rect 30136 23154 30192 23156
rect 30136 23102 30138 23154
rect 30138 23102 30190 23154
rect 30190 23102 30192 23154
rect 30136 23100 30192 23102
rect 30828 25730 30884 25732
rect 30828 25678 30830 25730
rect 30830 25678 30882 25730
rect 30882 25678 30884 25730
rect 30828 25676 30884 25678
rect 29036 21756 29092 21812
rect 28812 21644 28868 21700
rect 30248 22370 30304 22372
rect 30248 22318 30250 22370
rect 30250 22318 30302 22370
rect 30302 22318 30304 22370
rect 30248 22316 30304 22318
rect 31276 22204 31332 22260
rect 29036 20972 29092 21028
rect 29260 20802 29316 20804
rect 29260 20750 29262 20802
rect 29262 20750 29314 20802
rect 29314 20750 29316 20802
rect 29260 20748 29316 20750
rect 29540 21026 29596 21028
rect 29540 20974 29542 21026
rect 29542 20974 29594 21026
rect 29594 20974 29596 21026
rect 29540 20972 29596 20974
rect 28700 20076 28756 20132
rect 29092 20018 29148 20020
rect 29092 19966 29094 20018
rect 29094 19966 29146 20018
rect 29146 19966 29148 20018
rect 29092 19964 29148 19966
rect 28140 18620 28196 18676
rect 26908 18508 26964 18564
rect 27692 18508 27748 18564
rect 26180 18338 26236 18340
rect 26180 18286 26182 18338
rect 26182 18286 26234 18338
rect 26234 18286 26236 18338
rect 26180 18284 26236 18286
rect 26460 18284 26516 18340
rect 27132 18284 27188 18340
rect 27804 18413 27806 18452
rect 27806 18413 27858 18452
rect 27858 18413 27860 18452
rect 27804 18396 27860 18413
rect 27412 17442 27468 17444
rect 27412 17390 27414 17442
rect 27414 17390 27466 17442
rect 27466 17390 27468 17442
rect 27412 17388 27468 17390
rect 28364 18620 28420 18676
rect 28924 18620 28980 18676
rect 28756 18450 28812 18452
rect 28756 18398 28758 18450
rect 28758 18398 28810 18450
rect 28810 18398 28812 18450
rect 28756 18396 28812 18398
rect 28756 18060 28812 18116
rect 27804 17388 27860 17444
rect 28028 17164 28084 17220
rect 28476 16940 28532 16996
rect 27468 16716 27524 16772
rect 24444 14476 24500 14532
rect 25900 14588 25956 14644
rect 27020 14642 27076 14644
rect 27020 14590 27022 14642
rect 27022 14590 27074 14642
rect 27074 14590 27076 14642
rect 27020 14588 27076 14590
rect 27860 16210 27916 16212
rect 27860 16158 27862 16210
rect 27862 16158 27914 16210
rect 27914 16158 27916 16210
rect 27860 16156 27916 16158
rect 28364 16882 28420 16884
rect 28364 16830 28366 16882
rect 28366 16830 28418 16882
rect 28418 16830 28420 16882
rect 28364 16828 28420 16830
rect 28868 16716 28924 16772
rect 29148 18508 29204 18564
rect 29260 18396 29316 18452
rect 29148 18172 29204 18228
rect 29148 16940 29204 16996
rect 29428 18338 29484 18340
rect 29428 18286 29430 18338
rect 29430 18286 29482 18338
rect 29482 18286 29484 18338
rect 29428 18284 29484 18286
rect 31052 19740 31108 19796
rect 30156 18450 30212 18452
rect 30156 18398 30158 18450
rect 30158 18398 30210 18450
rect 30210 18398 30212 18450
rect 34300 26796 34356 26852
rect 33964 26290 34020 26292
rect 33964 26238 33966 26290
rect 33966 26238 34018 26290
rect 34018 26238 34020 26290
rect 33964 26236 34020 26238
rect 34076 26124 34132 26180
rect 32060 25452 32116 25508
rect 31948 23100 32004 23156
rect 31388 21644 31444 21700
rect 32396 25340 32452 25396
rect 32191 22204 32247 22260
rect 32060 20748 32116 20804
rect 32060 20188 32116 20244
rect 32228 19628 32284 19684
rect 30156 18396 30212 18398
rect 29596 17164 29652 17220
rect 31836 17612 31892 17668
rect 30156 16940 30212 16996
rect 29260 16882 29316 16884
rect 29260 16830 29262 16882
rect 29262 16830 29314 16882
rect 29314 16830 29316 16882
rect 29260 16828 29316 16830
rect 30044 16828 30100 16884
rect 29036 16268 29092 16324
rect 28588 15314 28644 15316
rect 28588 15262 28590 15314
rect 28590 15262 28642 15314
rect 28642 15262 28644 15314
rect 28588 15260 28644 15262
rect 28140 15148 28196 15204
rect 24892 14306 24948 14308
rect 24892 14254 24894 14306
rect 24894 14254 24946 14306
rect 24946 14254 24948 14306
rect 24892 14252 24948 14254
rect 27244 14252 27300 14308
rect 21532 13244 21588 13300
rect 14364 10108 14420 10164
rect 19852 11788 19908 11844
rect 18172 11452 18228 11508
rect 19740 11506 19796 11508
rect 19740 11454 19742 11506
rect 19742 11454 19794 11506
rect 19794 11454 19796 11506
rect 19740 11452 19796 11454
rect 20524 11788 20580 11844
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 21756 10668 21812 10724
rect 20972 9212 21028 9268
rect 13468 8258 13524 8260
rect 13468 8206 13470 8258
rect 13470 8206 13522 8258
rect 13522 8206 13524 8258
rect 13468 8204 13524 8206
rect 13132 5852 13188 5908
rect 13804 8204 13860 8260
rect 19180 8988 19236 9044
rect 19740 9042 19796 9044
rect 19740 8990 19742 9042
rect 19742 8990 19794 9042
rect 19794 8990 19796 9042
rect 19740 8988 19796 8990
rect 20188 8988 20244 9044
rect 19964 8428 20020 8484
rect 14140 7532 14196 7588
rect 14028 5852 14084 5908
rect 13580 5180 13636 5236
rect 13804 5180 13860 5236
rect 15932 5234 15988 5236
rect 15932 5182 15934 5234
rect 15934 5182 15986 5234
rect 15986 5182 15988 5234
rect 15932 5180 15988 5182
rect 19740 8316 19796 8372
rect 18396 7980 18452 8036
rect 19740 7980 19796 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20804 8540 20860 8596
rect 20804 8316 20860 8372
rect 20300 7980 20356 8036
rect 20356 6466 20412 6468
rect 20356 6414 20358 6466
rect 20358 6414 20410 6466
rect 20410 6414 20412 6466
rect 20356 6412 20412 6414
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19740 6076 19796 6132
rect 20356 6076 20412 6132
rect 21868 8988 21924 9044
rect 21644 8370 21700 8372
rect 21644 8318 21646 8370
rect 21646 8318 21698 8370
rect 21698 8318 21700 8370
rect 21644 8316 21700 8318
rect 22484 10722 22540 10724
rect 22484 10670 22486 10722
rect 22486 10670 22538 10722
rect 22538 10670 22540 10722
rect 22484 10668 22540 10670
rect 22204 10610 22260 10612
rect 22204 10558 22206 10610
rect 22206 10558 22258 10610
rect 22258 10558 22260 10610
rect 22204 10556 22260 10558
rect 23772 10556 23828 10612
rect 24444 10610 24500 10612
rect 24444 10558 24446 10610
rect 24446 10558 24498 10610
rect 24498 10558 24500 10610
rect 24444 10556 24500 10558
rect 24612 10556 24668 10612
rect 25754 10780 25810 10836
rect 26516 10834 26572 10836
rect 26516 10782 26518 10834
rect 26518 10782 26570 10834
rect 26570 10782 26572 10834
rect 26516 10780 26572 10782
rect 24444 9660 24500 9716
rect 24220 8316 24276 8372
rect 22316 8258 22372 8260
rect 22316 8206 22318 8258
rect 22318 8206 22370 8258
rect 22370 8206 22372 8258
rect 22316 8204 22372 8206
rect 26012 10610 26068 10612
rect 26012 10558 26014 10610
rect 26014 10558 26066 10610
rect 26066 10558 26068 10610
rect 26012 10556 26068 10558
rect 26684 10556 26740 10612
rect 26572 9884 26628 9940
rect 25900 9772 25956 9828
rect 25676 9042 25732 9044
rect 25676 8990 25678 9042
rect 25678 8990 25730 9042
rect 25730 8990 25732 9042
rect 25676 8988 25732 8990
rect 25900 8428 25956 8484
rect 27020 9811 27076 9828
rect 27020 9772 27022 9811
rect 27022 9772 27074 9811
rect 27074 9772 27076 9811
rect 27132 8988 27188 9044
rect 20972 6412 21028 6468
rect 19964 5906 20020 5908
rect 19964 5854 19966 5906
rect 19966 5854 20018 5906
rect 20018 5854 20020 5906
rect 19964 5852 20020 5854
rect 20468 5906 20524 5908
rect 20468 5854 20470 5906
rect 20470 5854 20522 5906
rect 20522 5854 20524 5906
rect 20468 5852 20524 5854
rect 16716 5180 16772 5236
rect 17444 5234 17500 5236
rect 17444 5182 17446 5234
rect 17446 5182 17498 5234
rect 17498 5182 17500 5234
rect 17444 5180 17500 5182
rect 20412 5628 20468 5684
rect 20300 5234 20356 5236
rect 20300 5182 20302 5234
rect 20302 5182 20354 5234
rect 20354 5182 20356 5234
rect 20300 5180 20356 5182
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21588 5682 21644 5684
rect 21588 5630 21590 5682
rect 21590 5630 21642 5682
rect 21642 5630 21644 5682
rect 21588 5628 21644 5630
rect 20860 5180 20916 5236
rect 22820 5906 22876 5908
rect 22820 5854 22822 5906
rect 22822 5854 22874 5906
rect 22874 5854 22876 5906
rect 22820 5852 22876 5854
rect 23548 5906 23604 5908
rect 23548 5854 23550 5906
rect 23550 5854 23602 5906
rect 23602 5854 23604 5906
rect 23548 5852 23604 5854
rect 22540 5628 22596 5684
rect 27132 6300 27188 6356
rect 27468 9884 27524 9940
rect 27804 10332 27860 10388
rect 29148 16156 29204 16212
rect 29148 15820 29204 15876
rect 29708 15484 29764 15540
rect 29036 15148 29092 15204
rect 29540 15148 29596 15204
rect 29876 15372 29932 15428
rect 31164 16716 31220 16772
rect 30940 16604 30996 16660
rect 30156 16322 30212 16324
rect 30156 16270 30158 16322
rect 30158 16270 30210 16322
rect 30210 16270 30212 16322
rect 30156 16268 30212 16270
rect 30940 15372 30996 15428
rect 30436 15314 30492 15316
rect 30436 15262 30438 15314
rect 30438 15262 30490 15314
rect 30490 15262 30492 15314
rect 30436 15260 30492 15262
rect 29708 10780 29764 10836
rect 31480 10610 31536 10612
rect 31480 10558 31482 10610
rect 31482 10558 31534 10610
rect 31534 10558 31536 10610
rect 31480 10556 31536 10558
rect 31724 10386 31780 10388
rect 31724 10334 31726 10386
rect 31726 10334 31778 10386
rect 31778 10334 31780 10386
rect 31724 10332 31780 10334
rect 30156 10108 30212 10164
rect 34300 25340 34356 25396
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34972 30156 35028 30212
rect 34806 28642 34862 28644
rect 34806 28590 34808 28642
rect 34808 28590 34860 28642
rect 34860 28590 34862 28642
rect 34806 28588 34862 28590
rect 36092 34242 36148 34244
rect 36092 34190 36094 34242
rect 36094 34190 36146 34242
rect 36146 34190 36148 34242
rect 36092 34188 36148 34190
rect 35980 31106 36036 31108
rect 35980 31054 35982 31106
rect 35982 31054 36034 31106
rect 36034 31054 36036 31106
rect 35980 31052 36036 31054
rect 35644 30156 35700 30212
rect 35532 30044 35588 30100
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 28812 35140 28868
rect 35868 28700 35924 28756
rect 35644 27692 35700 27748
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35532 27244 35588 27300
rect 34916 26850 34972 26852
rect 34916 26798 34918 26850
rect 34918 26798 34970 26850
rect 34970 26798 34972 26850
rect 34916 26796 34972 26798
rect 35196 26796 35252 26852
rect 34636 26236 34692 26292
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35532 25452 35588 25508
rect 35868 27468 35924 27524
rect 36316 31778 36372 31780
rect 36316 31726 36318 31778
rect 36318 31726 36370 31778
rect 36370 31726 36372 31778
rect 36316 31724 36372 31726
rect 36204 31500 36260 31556
rect 36428 30156 36484 30212
rect 37100 35756 37156 35812
rect 38892 35756 38948 35812
rect 36652 35698 36708 35700
rect 36652 35646 36654 35698
rect 36654 35646 36706 35698
rect 36706 35646 36708 35698
rect 36652 35644 36708 35646
rect 37976 35698 38032 35700
rect 37976 35646 37978 35698
rect 37978 35646 38030 35698
rect 38030 35646 38032 35698
rect 37976 35644 38032 35646
rect 39676 36204 39732 36260
rect 39228 35644 39284 35700
rect 40124 36316 40180 36372
rect 38220 34860 38276 34916
rect 38892 34914 38948 34916
rect 36764 32674 36820 32676
rect 36764 32622 36766 32674
rect 36766 32622 36818 32674
rect 36818 32622 36820 32674
rect 36764 32620 36820 32622
rect 37100 32562 37156 32564
rect 36652 32396 36708 32452
rect 37100 32510 37102 32562
rect 37102 32510 37154 32562
rect 37154 32510 37156 32562
rect 37100 32508 37156 32510
rect 37660 32562 37716 32564
rect 37660 32510 37662 32562
rect 37662 32510 37714 32562
rect 37714 32510 37716 32562
rect 37660 32508 37716 32510
rect 38892 34862 38894 34914
rect 38894 34862 38946 34914
rect 38946 34862 38948 34914
rect 38892 34860 38948 34862
rect 38612 34636 38668 34692
rect 38780 34802 38836 34804
rect 38780 34750 38782 34802
rect 38782 34750 38834 34802
rect 38834 34750 38836 34802
rect 38780 34748 38836 34750
rect 38444 32508 38500 32564
rect 37324 31948 37380 32004
rect 36876 31778 36932 31780
rect 36876 31726 36878 31778
rect 36878 31726 36930 31778
rect 36930 31726 36932 31778
rect 36876 31724 36932 31726
rect 37044 31554 37100 31556
rect 37044 31502 37046 31554
rect 37046 31502 37098 31554
rect 37098 31502 37100 31554
rect 37044 31500 37100 31502
rect 36540 29148 36596 29204
rect 36148 28530 36204 28532
rect 36148 28478 36150 28530
rect 36150 28478 36202 28530
rect 36202 28478 36204 28530
rect 36148 28476 36204 28478
rect 34412 24498 34468 24500
rect 34412 24446 34414 24498
rect 34414 24446 34466 24498
rect 34466 24446 34468 24498
rect 34412 24444 34468 24446
rect 35644 24444 35700 24500
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35476 23436 35532 23492
rect 34860 22876 34916 22932
rect 34524 22482 34580 22484
rect 34524 22430 34526 22482
rect 34526 22430 34578 22482
rect 34578 22430 34580 22482
rect 34524 22428 34580 22430
rect 34280 22370 34336 22372
rect 34280 22318 34282 22370
rect 34282 22318 34334 22370
rect 34334 22318 34336 22370
rect 34280 22316 34336 22318
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34860 22204 34916 22260
rect 33292 21644 33348 21700
rect 33124 20076 33180 20132
rect 35028 22316 35084 22372
rect 33404 21532 33460 21588
rect 34524 21586 34580 21588
rect 34524 21534 34526 21586
rect 34526 21534 34578 21586
rect 34578 21534 34580 21586
rect 34524 21532 34580 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 37100 28588 37156 28644
rect 39340 34972 39396 35028
rect 40572 34972 40628 35028
rect 40404 34914 40460 34916
rect 40404 34862 40406 34914
rect 40406 34862 40458 34914
rect 40458 34862 40460 34914
rect 40404 34860 40460 34862
rect 39676 32508 39732 32564
rect 40012 34802 40068 34804
rect 40012 34750 40014 34802
rect 40014 34750 40066 34802
rect 40066 34750 40068 34802
rect 40012 34748 40068 34750
rect 39788 34636 39844 34692
rect 39004 30044 39060 30100
rect 39340 30210 39396 30212
rect 39340 30158 39342 30210
rect 39342 30158 39394 30210
rect 39394 30158 39396 30210
rect 42924 39618 42980 39620
rect 42924 39566 42926 39618
rect 42926 39566 42978 39618
rect 42978 39566 42980 39618
rect 42924 39564 42980 39566
rect 43316 39618 43372 39620
rect 43316 39566 43318 39618
rect 43318 39566 43370 39618
rect 43370 39566 43372 39618
rect 43316 39564 43372 39566
rect 41132 36876 41188 36932
rect 42364 36876 42420 36932
rect 41132 36316 41188 36372
rect 41300 36258 41356 36260
rect 41300 36206 41302 36258
rect 41302 36206 41354 36258
rect 41354 36206 41356 36258
rect 41300 36204 41356 36206
rect 40964 34914 41020 34916
rect 40964 34862 40966 34914
rect 40966 34862 41018 34914
rect 41018 34862 41020 34914
rect 40964 34860 41020 34862
rect 42812 35308 42868 35364
rect 41580 34972 41636 35028
rect 41356 34636 41412 34692
rect 43820 35308 43876 35364
rect 40908 32562 40964 32564
rect 40908 32510 40910 32562
rect 40910 32510 40962 32562
rect 40962 32510 40964 32562
rect 41244 32674 41300 32676
rect 41244 32622 41246 32674
rect 41246 32622 41298 32674
rect 41298 32622 41300 32674
rect 41244 32620 41300 32622
rect 40908 32508 40964 32510
rect 41244 31500 41300 31556
rect 42644 34690 42700 34692
rect 42644 34638 42646 34690
rect 42646 34638 42698 34690
rect 42698 34638 42700 34690
rect 42644 34636 42700 34638
rect 41356 32396 41412 32452
rect 39340 30156 39396 30158
rect 38780 28588 38836 28644
rect 39004 28588 39060 28644
rect 37940 27970 37996 27972
rect 37940 27918 37942 27970
rect 37942 27918 37994 27970
rect 37994 27918 37996 27970
rect 37940 27916 37996 27918
rect 38444 27858 38500 27860
rect 38444 27806 38446 27858
rect 38446 27806 38498 27858
rect 38498 27806 38500 27858
rect 38444 27804 38500 27806
rect 37884 27692 37940 27748
rect 36484 26962 36540 26964
rect 36484 26910 36486 26962
rect 36486 26910 36538 26962
rect 36538 26910 36540 26962
rect 36484 26908 36540 26910
rect 36652 27468 36708 27524
rect 37212 27298 37268 27300
rect 37212 27246 37214 27298
rect 37214 27246 37266 27298
rect 37266 27246 37268 27298
rect 37212 27244 37268 27246
rect 39452 27356 39508 27412
rect 36652 27020 36708 27076
rect 37324 26908 37380 26964
rect 35980 22876 36036 22932
rect 36316 23938 36372 23940
rect 36316 23886 36318 23938
rect 36318 23886 36370 23938
rect 36370 23886 36372 23938
rect 36316 23884 36372 23886
rect 37100 26290 37156 26292
rect 37100 26238 37102 26290
rect 37102 26238 37154 26290
rect 37154 26238 37156 26290
rect 37100 26236 37156 26238
rect 36092 23436 36148 23492
rect 36708 23042 36764 23044
rect 36708 22990 36710 23042
rect 36710 22990 36762 23042
rect 36762 22990 36764 23042
rect 36708 22988 36764 22990
rect 36092 22540 36148 22596
rect 35980 22370 36036 22372
rect 33404 20188 33460 20244
rect 35980 22318 35982 22370
rect 35982 22318 36034 22370
rect 36034 22318 36036 22370
rect 35980 22316 36036 22318
rect 36372 22370 36428 22372
rect 36372 22318 36374 22370
rect 36374 22318 36426 22370
rect 36426 22318 36428 22370
rect 36372 22316 36428 22318
rect 33124 19740 33180 19796
rect 35364 19964 35420 20020
rect 34972 19628 35028 19684
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 36092 20300 36148 20356
rect 35980 20188 36036 20244
rect 35812 20076 35868 20132
rect 35644 20018 35700 20020
rect 35644 19966 35646 20018
rect 35646 19966 35698 20018
rect 35698 19966 35700 20018
rect 35644 19964 35700 19966
rect 35532 19404 35588 19460
rect 35644 18396 35700 18452
rect 34076 18060 34132 18116
rect 32956 16604 33012 16660
rect 33684 17612 33740 17668
rect 33404 15820 33460 15876
rect 32508 15484 32564 15540
rect 31948 15277 31950 15316
rect 31950 15277 32002 15316
rect 32002 15277 32004 15316
rect 31948 15260 32004 15277
rect 32732 15148 32788 15204
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36092 18450 36148 18452
rect 36092 18398 36094 18450
rect 36094 18398 36146 18450
rect 36146 18398 36148 18450
rect 36092 18396 36148 18398
rect 36484 18450 36540 18452
rect 36484 18398 36486 18450
rect 36486 18398 36538 18450
rect 36538 18398 36540 18450
rect 36484 18396 36540 18398
rect 37100 23884 37156 23940
rect 37436 26066 37492 26068
rect 37436 26014 37438 26066
rect 37438 26014 37490 26066
rect 37490 26014 37492 26066
rect 37436 26012 37492 26014
rect 34188 17106 34244 17108
rect 34188 17054 34190 17106
rect 34190 17054 34242 17106
rect 34242 17054 34244 17106
rect 34188 17052 34244 17054
rect 36988 17052 37044 17108
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 37996 23714 38052 23716
rect 37996 23662 37998 23714
rect 37998 23662 38050 23714
rect 38050 23662 38052 23714
rect 37996 23660 38052 23662
rect 37100 22988 37156 23044
rect 37548 20076 37604 20132
rect 37548 18396 37604 18452
rect 38668 20188 38724 20244
rect 37324 18284 37380 18340
rect 38668 18172 38724 18228
rect 37100 16940 37156 16996
rect 37492 16994 37548 16996
rect 37492 16942 37494 16994
rect 37494 16942 37546 16994
rect 37546 16942 37548 16994
rect 37492 16940 37548 16942
rect 38332 16716 38388 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 37996 15596 38052 15652
rect 34972 15314 35028 15316
rect 34972 15262 34974 15314
rect 34974 15262 35026 15314
rect 35026 15262 35028 15314
rect 34972 15260 35028 15262
rect 36316 15260 36372 15316
rect 33796 14530 33852 14532
rect 33796 14478 33798 14530
rect 33798 14478 33850 14530
rect 33850 14478 33852 14530
rect 33796 14476 33852 14478
rect 34076 14530 34132 14532
rect 34076 14478 34078 14530
rect 34078 14478 34130 14530
rect 34130 14478 34132 14530
rect 34076 14476 34132 14478
rect 33628 13746 33684 13748
rect 33628 13694 33630 13746
rect 33630 13694 33682 13746
rect 33682 13694 33684 13746
rect 33628 13692 33684 13694
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34188 13020 34244 13076
rect 38332 15426 38388 15428
rect 38332 15374 38334 15426
rect 38334 15374 38386 15426
rect 38386 15374 38388 15426
rect 38332 15372 38388 15374
rect 38164 15314 38220 15316
rect 38164 15262 38166 15314
rect 38166 15262 38218 15314
rect 38218 15262 38220 15314
rect 38164 15260 38220 15262
rect 38668 16716 38724 16772
rect 39452 27074 39508 27076
rect 39452 27022 39454 27074
rect 39454 27022 39506 27074
rect 39506 27022 39508 27074
rect 39452 27020 39508 27022
rect 40236 30044 40292 30100
rect 41224 30210 41280 30212
rect 41224 30158 41226 30210
rect 41226 30158 41278 30210
rect 41278 30158 41280 30210
rect 41224 30156 41280 30158
rect 41692 31500 41748 31556
rect 39900 27468 39956 27524
rect 39676 27020 39732 27076
rect 39788 26908 39844 26964
rect 39116 26012 39172 26068
rect 40012 26908 40068 26964
rect 39228 24668 39284 24724
rect 41076 28364 41132 28420
rect 40908 27858 40964 27860
rect 40908 27806 40910 27858
rect 40910 27806 40962 27858
rect 40962 27806 40964 27858
rect 40908 27804 40964 27806
rect 41244 27692 41300 27748
rect 41076 27244 41132 27300
rect 40908 27132 40964 27188
rect 42140 30828 42196 30884
rect 43820 30882 43876 30884
rect 43820 30830 43822 30882
rect 43822 30830 43874 30882
rect 43874 30830 43876 30882
rect 43820 30828 43876 30830
rect 42140 30210 42196 30212
rect 42140 30158 42142 30210
rect 42142 30158 42194 30210
rect 42194 30158 42196 30210
rect 42140 30156 42196 30158
rect 41692 28364 41748 28420
rect 40236 26124 40292 26180
rect 40124 24668 40180 24724
rect 41244 25228 41300 25284
rect 39228 23660 39284 23716
rect 39060 22370 39116 22372
rect 39060 22318 39062 22370
rect 39062 22318 39114 22370
rect 39114 22318 39116 22370
rect 39060 22316 39116 22318
rect 39116 20300 39172 20356
rect 39452 21756 39508 21812
rect 39340 21644 39396 21700
rect 42812 25506 42868 25508
rect 42812 25454 42814 25506
rect 42814 25454 42866 25506
rect 42866 25454 42868 25506
rect 42812 25452 42868 25454
rect 43820 25452 43876 25508
rect 41580 25228 41636 25284
rect 42644 25282 42700 25284
rect 42644 25230 42646 25282
rect 42646 25230 42698 25282
rect 42698 25230 42700 25282
rect 42644 25228 42700 25230
rect 39564 21586 39620 21588
rect 39564 21534 39566 21586
rect 39566 21534 39618 21586
rect 39618 21534 39620 21586
rect 39900 21756 39956 21812
rect 39564 21532 39620 21534
rect 39732 21308 39788 21364
rect 40012 21644 40068 21700
rect 40012 20300 40068 20356
rect 39900 20188 39956 20244
rect 40908 21586 40964 21588
rect 40908 21534 40910 21586
rect 40910 21534 40962 21586
rect 40962 21534 40964 21586
rect 41244 21756 41300 21812
rect 41356 21644 41412 21700
rect 40908 21532 40964 21534
rect 41244 21308 41300 21364
rect 42644 21362 42700 21364
rect 42644 21310 42646 21362
rect 42646 21310 42698 21362
rect 42698 21310 42700 21362
rect 42644 21308 42700 21310
rect 40236 19628 40292 19684
rect 40572 20076 40628 20132
rect 39564 19458 39620 19460
rect 39564 19406 39566 19458
rect 39566 19406 39618 19458
rect 39618 19406 39620 19458
rect 39564 19404 39620 19406
rect 39004 18284 39060 18340
rect 39340 18172 39396 18228
rect 39340 16716 39396 16772
rect 40740 19628 40796 19684
rect 40908 19404 40964 19460
rect 41356 19404 41412 19460
rect 41020 18450 41076 18452
rect 41020 18398 41022 18450
rect 41022 18398 41074 18450
rect 41074 18398 41076 18450
rect 41020 18396 41076 18398
rect 43596 18396 43652 18452
rect 39004 15596 39060 15652
rect 39340 15596 39396 15652
rect 38780 15484 38836 15540
rect 39004 15372 39060 15428
rect 38724 15314 38780 15316
rect 38724 15262 38726 15314
rect 38726 15262 38778 15314
rect 38778 15262 38780 15314
rect 38724 15260 38780 15262
rect 38444 15148 38500 15204
rect 38892 15148 38948 15204
rect 39564 15484 39620 15540
rect 36932 14364 36988 14420
rect 36932 13692 36988 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 38220 13074 38276 13076
rect 38220 13022 38222 13074
rect 38222 13022 38274 13074
rect 38274 13022 38276 13074
rect 38220 13020 38276 13022
rect 38332 12124 38388 12180
rect 39822 15299 39824 15316
rect 39824 15299 39876 15316
rect 39876 15299 39878 15316
rect 39822 15260 39878 15299
rect 39228 12908 39284 12964
rect 39900 12962 39956 12964
rect 39900 12910 39902 12962
rect 39902 12910 39954 12962
rect 39954 12910 39956 12962
rect 39900 12908 39956 12910
rect 39340 12178 39396 12180
rect 39340 12126 39342 12178
rect 39342 12126 39394 12178
rect 39394 12126 39396 12178
rect 39340 12124 39396 12126
rect 40236 15090 40292 15092
rect 40236 15038 40238 15090
rect 40238 15038 40290 15090
rect 40290 15038 40292 15090
rect 40236 15036 40292 15038
rect 43820 15484 43876 15540
rect 40348 14476 40404 14532
rect 40460 15036 40516 15092
rect 41132 14530 41188 14532
rect 41132 14478 41134 14530
rect 41134 14478 41186 14530
rect 41186 14478 41188 14530
rect 41132 14476 41188 14478
rect 30940 10108 30996 10164
rect 30548 9938 30604 9940
rect 30548 9886 30550 9938
rect 30550 9886 30602 9938
rect 30602 9886 30604 9938
rect 30548 9884 30604 9886
rect 32172 10556 32228 10612
rect 28588 9660 28644 9716
rect 27412 9266 27468 9268
rect 27412 9214 27414 9266
rect 27414 9214 27466 9266
rect 27466 9214 27468 9266
rect 27412 9212 27468 9214
rect 31388 8988 31444 9044
rect 27244 8540 27300 8596
rect 32060 9660 32116 9716
rect 32956 10610 33012 10612
rect 32956 10558 32958 10610
rect 32958 10558 33010 10610
rect 33010 10558 33012 10610
rect 32956 10556 33012 10558
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 40012 12124 40068 12180
rect 40572 12124 40628 12180
rect 43708 12908 43764 12964
rect 41132 12178 41188 12180
rect 41132 12126 41134 12178
rect 41134 12126 41186 12178
rect 41186 12126 41188 12178
rect 41132 12124 41188 12126
rect 32172 9042 32228 9044
rect 32172 8990 32174 9042
rect 32174 8990 32226 9042
rect 32226 8990 32228 9042
rect 32172 8988 32228 8990
rect 30828 6690 30884 6692
rect 30828 6638 30830 6690
rect 30830 6638 30882 6690
rect 30882 6638 30884 6690
rect 30828 6636 30884 6638
rect 27244 6076 27300 6132
rect 27580 6300 27636 6356
rect 29596 6300 29652 6356
rect 28252 6076 28308 6132
rect 27916 5964 27972 6020
rect 27468 5794 27524 5796
rect 27468 5742 27470 5794
rect 27470 5742 27522 5794
rect 27522 5742 27524 5794
rect 27468 5740 27524 5742
rect 29484 5964 29540 6020
rect 28588 5740 28644 5796
rect 28924 5740 28980 5796
rect 26292 4284 26348 4340
rect 26908 4338 26964 4340
rect 26908 4286 26910 4338
rect 26910 4286 26962 4338
rect 26962 4286 26964 4338
rect 26908 4284 26964 4286
rect 30772 6130 30828 6132
rect 30772 6078 30774 6130
rect 30774 6078 30826 6130
rect 30826 6078 30828 6130
rect 30772 6076 30828 6078
rect 32396 9100 32452 9156
rect 33516 9100 33572 9156
rect 33404 9042 33460 9044
rect 33404 8990 33406 9042
rect 33406 8990 33458 9042
rect 33458 8990 33460 9042
rect 33404 8988 33460 8990
rect 34076 9266 34132 9268
rect 34076 9214 34078 9266
rect 34078 9214 34130 9266
rect 34130 9214 34132 9266
rect 34076 9212 34132 9214
rect 35420 9212 35476 9268
rect 36204 9826 36260 9828
rect 36204 9774 36206 9826
rect 36206 9774 36258 9826
rect 36258 9774 36260 9826
rect 36204 9772 36260 9774
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 31388 6636 31444 6692
rect 30940 5964 30996 6020
rect 31052 6076 31108 6132
rect 29876 5794 29932 5796
rect 29876 5742 29878 5794
rect 29878 5742 29930 5794
rect 29930 5742 29932 5794
rect 29876 5740 29932 5742
rect 31836 5852 31892 5908
rect 32956 5906 33012 5908
rect 32956 5854 32958 5906
rect 32958 5854 33010 5906
rect 33010 5854 33012 5906
rect 32956 5852 33012 5854
rect 31612 5740 31668 5796
rect 33292 5682 33348 5684
rect 33292 5630 33294 5682
rect 33294 5630 33346 5682
rect 33346 5630 33348 5682
rect 33292 5628 33348 5630
rect 34076 5628 34132 5684
rect 31276 5122 31332 5124
rect 31276 5070 31278 5122
rect 31278 5070 31330 5122
rect 31330 5070 31332 5122
rect 31276 5068 31332 5070
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34860 5180 34916 5236
rect 32172 5122 32228 5124
rect 32172 5070 32174 5122
rect 32174 5070 32226 5122
rect 32226 5070 32228 5122
rect 32172 5068 32228 5070
rect 35252 5234 35308 5236
rect 35252 5182 35254 5234
rect 35254 5182 35306 5234
rect 35306 5182 35308 5234
rect 35252 5180 35308 5182
rect 36876 9772 36932 9828
rect 36204 5180 36260 5236
rect 30212 4338 30268 4340
rect 30212 4286 30214 4338
rect 30214 4286 30266 4338
rect 30266 4286 30268 4338
rect 30212 4284 30268 4286
rect 18396 4172 18452 4228
rect 19964 4226 20020 4228
rect 19964 4174 19966 4226
rect 19966 4174 20018 4226
rect 20018 4174 20020 4226
rect 19964 4172 20020 4174
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 13234 41804 13244 41860
rect 13300 41804 14476 41860
rect 14532 41804 14542 41860
rect 17042 41804 17052 41860
rect 17108 41804 18284 41860
rect 18340 41804 18350 41860
rect 20850 41804 20860 41860
rect 20916 41804 22092 41860
rect 22148 41804 22158 41860
rect 24658 41804 24668 41860
rect 24724 41804 25900 41860
rect 25956 41804 25966 41860
rect 28466 41804 28476 41860
rect 28532 41804 29708 41860
rect 29764 41804 29774 41860
rect 32274 41804 32284 41860
rect 32340 41804 33516 41860
rect 33572 41804 33582 41860
rect 36082 41804 36092 41860
rect 36148 41804 37324 41860
rect 37380 41804 37390 41860
rect 39890 41804 39900 41860
rect 39956 41804 41132 41860
rect 41188 41804 41198 41860
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 11778 40572 11788 40628
rect 11844 40572 13468 40628
rect 13524 40572 13534 40628
rect 39666 40572 39676 40628
rect 39732 40572 40124 40628
rect 40180 40572 40190 40628
rect 15810 40460 15820 40516
rect 15876 40460 17276 40516
rect 17332 40460 17342 40516
rect 36082 40460 36092 40516
rect 36148 40460 39004 40516
rect 39060 40460 39340 40516
rect 39396 40460 39406 40516
rect 2146 40348 2156 40404
rect 2212 40348 5460 40404
rect 5516 40348 5740 40404
rect 5796 40348 6636 40404
rect 6692 40348 9044 40404
rect 9100 40348 9110 40404
rect 13458 40348 13468 40404
rect 13524 40348 14476 40404
rect 14532 40348 18396 40404
rect 18452 40348 18462 40404
rect 21858 40348 21868 40404
rect 21924 40348 25396 40404
rect 25452 40348 26012 40404
rect 26068 40348 28588 40404
rect 28644 40348 29316 40404
rect 29372 40348 29708 40404
rect 29764 40348 32788 40404
rect 32844 40348 32854 40404
rect 33282 40348 33292 40404
rect 33348 40348 36372 40404
rect 36428 40348 36438 40404
rect 5058 40236 5068 40292
rect 5124 40236 6524 40292
rect 6580 40236 6590 40292
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 19170 39788 19180 39844
rect 19236 39788 20188 39844
rect 20244 39788 20254 39844
rect 22642 39788 22652 39844
rect 22708 39788 24444 39844
rect 24500 39788 24510 39844
rect 32834 39788 32844 39844
rect 32900 39788 34076 39844
rect 34132 39788 34142 39844
rect 41794 39788 41804 39844
rect 41860 39788 42588 39844
rect 42644 39788 42654 39844
rect 17714 39676 17724 39732
rect 17780 39676 23660 39732
rect 23716 39676 23726 39732
rect 3042 39564 3052 39620
rect 3108 39564 4060 39620
rect 4116 39564 4620 39620
rect 4676 39564 4686 39620
rect 4834 39564 4844 39620
rect 4900 39564 9007 39620
rect 9063 39564 9073 39620
rect 14242 39564 14252 39620
rect 14308 39564 23436 39620
rect 23492 39564 23502 39620
rect 39330 39564 39340 39620
rect 39396 39564 42924 39620
rect 42980 39564 43316 39620
rect 43372 39564 43382 39620
rect 8754 39452 8764 39508
rect 8820 39452 10892 39508
rect 10948 39452 10958 39508
rect 20514 39452 20524 39508
rect 20580 39452 29148 39508
rect 29204 39452 29214 39508
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 12226 39004 12236 39060
rect 12292 39004 16044 39060
rect 16100 39004 16110 39060
rect 4274 38892 4284 38948
rect 4340 38892 5292 38948
rect 5348 38892 7756 38948
rect 7812 38892 7822 38948
rect 2650 38780 2660 38836
rect 2716 38780 4508 38836
rect 4564 38780 4574 38836
rect 8082 38780 8092 38836
rect 8148 38780 8428 38836
rect 8484 38780 9884 38836
rect 9940 38780 9950 38836
rect 10322 38780 10332 38836
rect 10388 38780 13468 38836
rect 13524 38780 13534 38836
rect 23538 38780 23548 38836
rect 23604 38780 24332 38836
rect 24388 38780 28924 38836
rect 28980 38780 29260 38836
rect 29316 38780 29326 38836
rect 3938 38668 3948 38724
rect 4004 38668 5068 38724
rect 5124 38668 5134 38724
rect 35802 38668 35812 38724
rect 35868 38668 36390 38724
rect 36446 38668 36456 38724
rect 3266 38556 3276 38612
rect 3332 38556 3836 38612
rect 3892 38556 3902 38612
rect 4162 38556 4172 38612
rect 4228 38556 4676 38612
rect 4732 38556 4742 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 24434 38220 24444 38276
rect 24500 38220 24510 38276
rect 24444 37940 24500 38220
rect 28018 37996 28028 38052
rect 28084 37996 28364 38052
rect 28420 37996 29036 38052
rect 29092 37996 29102 38052
rect 23650 37884 23660 37940
rect 23716 37884 23996 37940
rect 24052 37884 29540 37940
rect 29596 37884 29606 37940
rect 4332 37772 4342 37828
rect 4398 37772 5124 37828
rect 5180 37772 6412 37828
rect 6468 37772 6478 37828
rect 23820 37772 23830 37828
rect 23886 37772 25004 37828
rect 25060 37772 25070 37828
rect 28690 37772 28700 37828
rect 28756 37772 30156 37828
rect 30212 37772 32956 37828
rect 33012 37772 33022 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 26338 37324 26348 37380
rect 26404 37324 27804 37380
rect 27860 37324 27870 37380
rect 29362 37324 29372 37380
rect 29428 37324 32508 37380
rect 32564 37324 32574 37380
rect 3938 37212 3948 37268
rect 4004 37212 4844 37268
rect 4900 37212 5124 37268
rect 5180 37212 5190 37268
rect 25890 37212 25900 37268
rect 25956 37212 27580 37268
rect 27636 37212 27646 37268
rect 4050 37100 4060 37156
rect 4116 37100 4688 37156
rect 4744 37100 6860 37156
rect 6916 37100 6926 37156
rect 16370 37100 16380 37156
rect 16436 37100 18060 37156
rect 18116 37100 18126 37156
rect 25554 37100 25564 37156
rect 25620 37100 26504 37156
rect 26560 37100 28700 37156
rect 28756 37100 28766 37156
rect 19516 36988 20524 37044
rect 20580 36988 20590 37044
rect 19516 36932 19572 36988
rect 19506 36876 19516 36932
rect 19572 36876 19582 36932
rect 41122 36876 41132 36932
rect 41188 36876 42364 36932
rect 42420 36876 42430 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 10098 36316 10108 36372
rect 10164 36316 10780 36372
rect 10836 36316 10846 36372
rect 40114 36316 40124 36372
rect 40180 36316 41132 36372
rect 41188 36316 41198 36372
rect 33730 36204 33740 36260
rect 33796 36204 34132 36260
rect 34188 36204 36540 36260
rect 36596 36204 37156 36260
rect 37212 36204 39676 36260
rect 39732 36204 41300 36260
rect 41356 36204 41366 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 6626 35868 6636 35924
rect 6692 35868 7308 35924
rect 7364 35868 7374 35924
rect 37090 35756 37100 35812
rect 37156 35756 38892 35812
rect 38948 35756 38958 35812
rect 10770 35644 10780 35700
rect 10836 35644 13916 35700
rect 13972 35644 14364 35700
rect 14420 35644 14430 35700
rect 16370 35644 16380 35700
rect 16436 35644 18396 35700
rect 18452 35644 18462 35700
rect 36418 35644 36428 35700
rect 36484 35644 36652 35700
rect 36708 35644 37976 35700
rect 38032 35644 38042 35700
rect 39218 35644 39228 35700
rect 39284 35644 39294 35700
rect 13458 35532 13468 35588
rect 13524 35532 16044 35588
rect 16100 35532 16604 35588
rect 16660 35532 17388 35588
rect 17444 35532 17454 35588
rect 14690 35308 14700 35364
rect 14756 35308 14766 35364
rect 28354 35308 28364 35364
rect 28420 35308 28958 35364
rect 29014 35308 29024 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 14700 34916 14756 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 26842 35196 26852 35252
rect 26908 35196 28812 35252
rect 28868 35196 29596 35252
rect 29652 35196 29662 35252
rect 39228 35028 39284 35644
rect 42802 35308 42812 35364
rect 42868 35308 43820 35364
rect 43876 35308 43886 35364
rect 39228 34972 39340 35028
rect 39396 34972 39406 35028
rect 40562 34972 40572 35028
rect 40628 34972 41580 35028
rect 41636 34972 41646 35028
rect 6402 34860 6412 34916
rect 6468 34860 7028 34916
rect 7084 34860 7094 34916
rect 14700 34860 15260 34916
rect 15316 34860 16268 34916
rect 16324 34860 16996 34916
rect 17266 34860 17276 34916
rect 17332 34860 18396 34916
rect 18452 34860 18462 34916
rect 23650 34860 23660 34916
rect 23716 34860 24836 34916
rect 24892 34860 25620 34916
rect 25676 34860 25686 34916
rect 25890 34860 25900 34916
rect 25956 34860 27356 34916
rect 27412 34860 27422 34916
rect 28018 34860 28028 34916
rect 28084 34860 28700 34916
rect 28756 34860 29148 34916
rect 29204 34860 29214 34916
rect 38210 34860 38220 34916
rect 38276 34860 38892 34916
rect 38948 34860 38958 34916
rect 40394 34860 40404 34916
rect 40460 34860 40964 34916
rect 41020 34860 41030 34916
rect 14700 34580 14756 34860
rect 16940 34804 16996 34860
rect 16930 34748 16940 34804
rect 16996 34748 17006 34804
rect 28466 34748 28476 34804
rect 28532 34748 30156 34804
rect 30212 34748 30222 34804
rect 38770 34748 38780 34804
rect 38836 34748 40012 34804
rect 40068 34748 40078 34804
rect 17994 34636 18004 34692
rect 18060 34636 18676 34692
rect 18732 34636 18742 34692
rect 25778 34636 25788 34692
rect 25844 34636 27804 34692
rect 27860 34636 29372 34692
rect 29428 34636 29438 34692
rect 38602 34636 38612 34692
rect 38668 34636 39788 34692
rect 39844 34636 39854 34692
rect 41346 34636 41356 34692
rect 41412 34636 42644 34692
rect 42700 34636 42710 34692
rect 14690 34524 14700 34580
rect 14756 34524 14766 34580
rect 17388 34524 18956 34580
rect 19012 34524 19292 34580
rect 19348 34524 19358 34580
rect 17388 34468 17444 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 14373 34412 14383 34468
rect 14439 34412 17444 34468
rect 17602 34412 17612 34468
rect 17668 34412 18620 34468
rect 18676 34412 18686 34468
rect 18274 34300 18284 34356
rect 18340 34300 18396 34356
rect 18452 34300 18462 34356
rect 28242 34300 28252 34356
rect 28308 34300 29260 34356
rect 29316 34300 29820 34356
rect 29876 34300 29886 34356
rect 12002 34188 12012 34244
rect 12068 34188 13860 34244
rect 13916 34188 13926 34244
rect 34738 34188 34748 34244
rect 34804 34188 36092 34244
rect 36148 34188 36158 34244
rect 4946 34076 4956 34132
rect 5012 34076 5628 34132
rect 5684 34076 5694 34132
rect 16762 34076 16772 34132
rect 16828 34076 17836 34132
rect 17892 34076 17902 34132
rect 18386 34076 18396 34132
rect 18452 34076 19628 34132
rect 19684 34076 19694 34132
rect 6178 33964 6188 34020
rect 6244 33964 21252 34020
rect 21308 33964 21980 34020
rect 22036 33964 22316 34020
rect 22372 33964 23044 34020
rect 23100 33964 23110 34020
rect 3266 33852 3276 33908
rect 3332 33852 4172 33908
rect 4228 33852 6804 33908
rect 6860 33852 6870 33908
rect 22474 33852 22484 33908
rect 22540 33852 23324 33908
rect 23380 33852 29988 33908
rect 30044 33852 32508 33908
rect 32564 33852 32574 33908
rect 5506 33740 5516 33796
rect 5572 33740 6412 33796
rect 6468 33740 6478 33796
rect 18162 33740 18172 33796
rect 18228 33740 18396 33796
rect 18452 33740 18462 33796
rect 18610 33740 18620 33796
rect 18676 33740 19404 33796
rect 19460 33740 19470 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 18620 33684 18676 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 18060 33628 18676 33684
rect 5180 33516 6524 33572
rect 6580 33516 6590 33572
rect 5114 33404 5124 33460
rect 5180 33404 5236 33516
rect 18060 33460 18116 33628
rect 21634 33516 21644 33572
rect 21700 33516 22596 33572
rect 22652 33516 23660 33572
rect 23716 33516 23726 33572
rect 27290 33516 27300 33572
rect 27356 33516 28476 33572
rect 28532 33516 28542 33572
rect 5394 33404 5404 33460
rect 5460 33404 6412 33460
rect 6468 33404 6478 33460
rect 18050 33404 18060 33460
rect 18116 33404 18126 33460
rect 20132 33404 20244 33460
rect 20300 33404 20310 33460
rect 29484 33404 30604 33460
rect 30660 33404 30670 33460
rect 20132 33348 20188 33404
rect 29484 33348 29540 33404
rect 5404 33292 5852 33348
rect 5908 33292 5918 33348
rect 8754 33292 8764 33348
rect 8820 33292 9212 33348
rect 9268 33292 9278 33348
rect 18440 33292 18450 33348
rect 18506 33292 19292 33348
rect 19348 33292 19460 33348
rect 19516 33292 20188 33348
rect 23650 33292 23660 33348
rect 23716 33292 24668 33348
rect 24724 33292 27132 33348
rect 27188 33292 27198 33348
rect 28690 33292 28700 33348
rect 28756 33292 29484 33348
rect 29540 33292 29550 33348
rect 29810 33292 29820 33348
rect 29876 33292 31276 33348
rect 31332 33292 31342 33348
rect 5404 33236 5460 33292
rect 5394 33180 5404 33236
rect 5460 33180 5470 33236
rect 5618 33068 5628 33124
rect 5684 33068 6524 33124
rect 6580 33068 8428 33124
rect 8484 33068 8494 33124
rect 18358 33068 18396 33124
rect 18452 33068 18462 33124
rect 21522 33068 21532 33124
rect 21588 33068 23268 33124
rect 23324 33068 23334 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 5282 32732 5292 32788
rect 5348 32732 5852 32788
rect 5908 32732 5918 32788
rect 22642 32620 22652 32676
rect 22708 32620 24556 32676
rect 24612 32620 24622 32676
rect 36754 32620 36764 32676
rect 36820 32620 41244 32676
rect 41300 32620 41310 32676
rect 4274 32508 4284 32564
rect 4340 32508 4508 32564
rect 4564 32508 6300 32564
rect 6356 32508 6860 32564
rect 6916 32508 6926 32564
rect 37090 32508 37100 32564
rect 37156 32508 37660 32564
rect 37716 32508 38444 32564
rect 38500 32508 39676 32564
rect 39732 32508 40908 32564
rect 40964 32508 40974 32564
rect 4610 32396 4620 32452
rect 4676 32396 7252 32452
rect 7308 32396 15036 32452
rect 15092 32396 15102 32452
rect 36642 32396 36652 32452
rect 36708 32396 41356 32452
rect 41412 32396 41422 32452
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 21186 32060 21196 32116
rect 21252 32060 22428 32116
rect 22484 32060 23324 32116
rect 23380 32060 23390 32116
rect 21970 31948 21980 32004
rect 22036 31948 28476 32004
rect 28532 31948 28542 32004
rect 32834 31948 32844 32004
rect 32900 31948 34636 32004
rect 34692 31948 37324 32004
rect 37380 31948 37390 32004
rect 21858 31836 21868 31892
rect 21924 31836 24668 31892
rect 24724 31836 25340 31892
rect 25396 31836 27748 31892
rect 27804 31836 28364 31892
rect 28420 31836 28588 31892
rect 28644 31836 30156 31892
rect 30212 31836 31836 31892
rect 31892 31836 33460 31892
rect 33516 31836 33526 31892
rect 12562 31724 12572 31780
rect 12628 31724 14812 31780
rect 14868 31724 14878 31780
rect 15474 31724 15484 31780
rect 15540 31724 16380 31780
rect 16436 31724 16446 31780
rect 16650 31724 16660 31780
rect 16716 31724 17164 31780
rect 17220 31724 17230 31780
rect 24546 31724 24556 31780
rect 24612 31724 25788 31780
rect 25844 31724 25854 31780
rect 36306 31724 36316 31780
rect 36372 31724 36876 31780
rect 36932 31724 36942 31780
rect 13794 31612 13804 31668
rect 13860 31612 16268 31668
rect 16324 31612 16334 31668
rect 16146 31500 16156 31556
rect 16212 31500 16716 31556
rect 16772 31500 16782 31556
rect 17490 31500 17500 31556
rect 17556 31500 18060 31556
rect 18116 31500 18844 31556
rect 18900 31500 18910 31556
rect 28186 31500 28196 31556
rect 28252 31500 29148 31556
rect 29204 31500 32564 31556
rect 32620 31500 33068 31556
rect 33124 31500 33134 31556
rect 36194 31500 36204 31556
rect 36260 31500 37044 31556
rect 37100 31500 37110 31556
rect 41234 31500 41244 31556
rect 41300 31500 41692 31556
rect 41748 31500 41758 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4946 31164 4956 31220
rect 5012 31164 5628 31220
rect 5684 31164 5694 31220
rect 8372 31164 11676 31220
rect 11732 31164 11742 31220
rect 8372 30996 8428 31164
rect 34402 31052 34412 31108
rect 34468 31052 35980 31108
rect 36036 31052 36046 31108
rect 7746 30940 7756 30996
rect 7812 30940 8428 30996
rect 8754 30940 8764 30996
rect 8820 30940 10108 30996
rect 10164 30940 10668 30996
rect 10724 30940 10734 30996
rect 11666 30940 11676 30996
rect 11732 30940 16044 30996
rect 16100 30940 16110 30996
rect 16258 30940 16268 30996
rect 16324 30940 17948 30996
rect 18004 30940 18284 30996
rect 18340 30940 18350 30996
rect 19170 30940 19180 30996
rect 19236 30940 20076 30996
rect 20132 30940 20142 30996
rect 27570 30940 27580 30996
rect 27636 30940 28700 30996
rect 28756 30940 28766 30996
rect 5506 30828 5516 30884
rect 5572 30828 16156 30884
rect 16212 30828 16222 30884
rect 42130 30828 42140 30884
rect 42196 30828 43820 30884
rect 43876 30828 43886 30884
rect 9982 30716 9992 30772
rect 10048 30716 12236 30772
rect 12292 30716 12302 30772
rect 16594 30716 16604 30772
rect 16660 30716 16828 30772
rect 16884 30716 17556 30772
rect 17612 30716 21532 30772
rect 21588 30716 21598 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 27122 30380 27132 30436
rect 27188 30380 28476 30436
rect 28532 30380 28542 30436
rect 16370 30268 16380 30324
rect 16436 30268 16446 30324
rect 17098 30268 17108 30324
rect 17164 30268 18732 30324
rect 18788 30268 18798 30324
rect 28476 30268 29148 30324
rect 29204 30268 29214 30324
rect 16380 30212 16436 30268
rect 28476 30212 28532 30268
rect 8306 30156 8316 30212
rect 8372 30156 9436 30212
rect 9492 30156 9502 30212
rect 11666 30156 11676 30212
rect 11732 30156 12852 30212
rect 12908 30156 13804 30212
rect 13860 30156 13870 30212
rect 16380 30156 22428 30212
rect 22484 30156 28532 30212
rect 34962 30156 34972 30212
rect 35028 30156 35644 30212
rect 35700 30156 36428 30212
rect 36484 30156 39340 30212
rect 39396 30156 39406 30212
rect 41214 30156 41224 30212
rect 41280 30156 42140 30212
rect 42196 30156 42206 30212
rect 12450 30044 12460 30100
rect 12516 30044 15148 30100
rect 15204 30044 15214 30100
rect 15362 30044 15372 30100
rect 15428 30044 16940 30100
rect 16996 30044 17006 30100
rect 17164 30044 17556 30100
rect 17612 30044 18284 30100
rect 18340 30044 18350 30100
rect 18508 30044 19964 30100
rect 20020 30044 20030 30100
rect 20402 30044 20412 30100
rect 20468 30044 21084 30100
rect 21140 30044 21476 30100
rect 21532 30044 21980 30100
rect 22036 30044 22046 30100
rect 26898 30044 26908 30100
rect 26964 30044 28140 30100
rect 28196 30044 28206 30100
rect 28466 30044 28476 30100
rect 28532 30044 35532 30100
rect 35588 30044 35598 30100
rect 38994 30044 39004 30100
rect 39060 30044 40236 30100
rect 40292 30044 40302 30100
rect 17164 29988 17220 30044
rect 16482 29932 16492 29988
rect 16548 29932 17220 29988
rect 18508 29876 18564 30044
rect 20178 29932 20188 29988
rect 20244 29932 24108 29988
rect 24164 29932 26684 29988
rect 26740 29932 26750 29988
rect 14130 29820 14140 29876
rect 14196 29820 18564 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 3714 29372 3724 29428
rect 3780 29372 5852 29428
rect 5908 29372 5918 29428
rect 6514 29372 6524 29428
rect 6580 29372 6972 29428
rect 7028 29372 7038 29428
rect 10770 29372 10780 29428
rect 10836 29372 11564 29428
rect 11620 29372 15260 29428
rect 15316 29372 16716 29428
rect 16772 29372 16782 29428
rect 19506 29372 19516 29428
rect 19572 29372 20860 29428
rect 20916 29372 20926 29428
rect 2594 29260 2604 29316
rect 2660 29260 3612 29316
rect 3668 29260 3678 29316
rect 14914 29260 14924 29316
rect 14980 29260 16212 29316
rect 16268 29260 16278 29316
rect 21410 29148 21420 29204
rect 21476 29148 36540 29204
rect 36596 29148 36606 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 13458 28924 13468 28980
rect 13524 28924 14140 28980
rect 14196 28924 14206 28980
rect 6626 28812 6636 28868
rect 6692 28812 8092 28868
rect 8148 28812 8158 28868
rect 20178 28812 20188 28868
rect 20244 28812 20636 28868
rect 20692 28812 20702 28868
rect 31378 28812 31388 28868
rect 31444 28812 35084 28868
rect 35140 28812 35150 28868
rect 6290 28700 6300 28756
rect 6356 28700 7756 28756
rect 7812 28700 7822 28756
rect 18274 28700 18284 28756
rect 18340 28700 22764 28756
rect 22820 28700 22830 28756
rect 35858 28700 35868 28756
rect 35924 28700 37156 28756
rect 37100 28644 37156 28700
rect 1810 28588 1820 28644
rect 1876 28588 5124 28644
rect 5180 28588 7980 28644
rect 8036 28588 8046 28644
rect 12562 28588 12572 28644
rect 12628 28588 13692 28644
rect 13748 28588 13758 28644
rect 20402 28588 20412 28644
rect 20468 28588 27020 28644
rect 27076 28588 27086 28644
rect 34796 28588 34806 28644
rect 34862 28588 36148 28644
rect 37090 28588 37100 28644
rect 37156 28588 38780 28644
rect 38836 28588 39004 28644
rect 39060 28588 39070 28644
rect 17378 28476 17388 28532
rect 17444 28476 19068 28532
rect 19124 28476 19134 28532
rect 36092 28476 36148 28588
rect 36204 28476 36214 28532
rect 4498 28364 4508 28420
rect 4564 28364 5068 28420
rect 5124 28364 5134 28420
rect 41066 28364 41076 28420
rect 41132 28364 41692 28420
rect 41748 28364 41758 28420
rect 8194 28252 8204 28308
rect 8260 28252 10332 28308
rect 10388 28252 10398 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4834 28028 4844 28084
rect 4900 28028 6132 28084
rect 6188 28028 6198 28084
rect 9314 28028 9324 28084
rect 9380 28028 10892 28084
rect 10948 28028 10958 28084
rect 17826 28028 17836 28084
rect 17892 28028 18788 28084
rect 18844 28028 19292 28084
rect 19348 28028 20188 28084
rect 20132 27972 20188 28028
rect 4050 27916 4060 27972
rect 4116 27916 5684 27972
rect 5740 27916 17500 27972
rect 17556 27916 17566 27972
rect 20132 27916 22652 27972
rect 22708 27916 37940 27972
rect 37996 27916 38006 27972
rect 18050 27804 18060 27860
rect 18116 27804 18620 27860
rect 18676 27804 25228 27860
rect 25284 27804 25564 27860
rect 25620 27804 25630 27860
rect 26562 27804 26572 27860
rect 26628 27804 29036 27860
rect 29092 27804 29102 27860
rect 38434 27804 38444 27860
rect 38500 27804 40908 27860
rect 40964 27804 40974 27860
rect 13906 27692 13916 27748
rect 13972 27692 16716 27748
rect 16772 27692 19404 27748
rect 19460 27692 19470 27748
rect 20132 27692 24724 27748
rect 24780 27692 25004 27748
rect 25060 27692 25900 27748
rect 25956 27692 25966 27748
rect 35634 27692 35644 27748
rect 35700 27692 37884 27748
rect 37940 27692 41244 27748
rect 41300 27692 41310 27748
rect 20132 27636 20188 27692
rect 18890 27580 18900 27636
rect 18956 27580 20188 27636
rect 35858 27468 35868 27524
rect 35924 27468 36652 27524
rect 36708 27468 36718 27524
rect 39452 27468 39900 27524
rect 39956 27468 39966 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 39452 27412 39508 27468
rect 39442 27356 39452 27412
rect 39508 27356 39518 27412
rect 35522 27244 35532 27300
rect 35588 27244 37212 27300
rect 37268 27244 41076 27300
rect 41132 27244 41142 27300
rect 39778 27132 39788 27188
rect 39844 27132 40908 27188
rect 40964 27132 40974 27188
rect 7410 27020 7420 27076
rect 7476 27020 14364 27076
rect 14420 27020 21756 27076
rect 21812 27020 21822 27076
rect 28242 27020 28252 27076
rect 28308 27020 29988 27076
rect 36642 27020 36652 27076
rect 36708 27020 39452 27076
rect 39508 27020 39518 27076
rect 39666 27020 39676 27076
rect 39732 27020 40068 27076
rect 29932 26964 29988 27020
rect 40012 26964 40068 27020
rect 14690 26908 14700 26964
rect 14756 26908 15260 26964
rect 15316 26908 15326 26964
rect 18498 26908 18508 26964
rect 18564 26908 18900 26964
rect 18956 26908 18966 26964
rect 26226 26908 26236 26964
rect 26292 26908 28364 26964
rect 28420 26908 28430 26964
rect 29922 26908 29932 26964
rect 29988 26908 30492 26964
rect 30548 26908 30558 26964
rect 36474 26908 36484 26964
rect 36540 26908 37324 26964
rect 37380 26908 37390 26964
rect 39750 26908 39788 26964
rect 39844 26908 39854 26964
rect 40002 26908 40012 26964
rect 40068 26908 40078 26964
rect 29698 26796 29708 26852
rect 29764 26796 30604 26852
rect 30660 26796 30670 26852
rect 34290 26796 34300 26852
rect 34356 26796 34916 26852
rect 34972 26796 35196 26852
rect 35252 26796 35262 26852
rect 28242 26684 28252 26740
rect 28308 26684 30268 26740
rect 30324 26684 30334 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 18218 26348 18228 26404
rect 18284 26348 19124 26404
rect 19180 26348 19190 26404
rect 9986 26236 9996 26292
rect 10052 26236 13916 26292
rect 13972 26236 17836 26292
rect 17892 26236 17902 26292
rect 18498 26236 18508 26292
rect 18564 26236 19124 26292
rect 21410 26236 21420 26292
rect 21476 26236 22540 26292
rect 22596 26236 22606 26292
rect 28914 26236 28924 26292
rect 28980 26236 29596 26292
rect 29652 26236 29662 26292
rect 33954 26236 33964 26292
rect 34020 26236 34636 26292
rect 34692 26236 37100 26292
rect 37156 26236 37166 26292
rect 19068 26180 19124 26236
rect 19058 26124 19068 26180
rect 19124 26124 19134 26180
rect 30350 26124 30360 26180
rect 30416 26124 31220 26180
rect 31276 26124 34076 26180
rect 34132 26124 40236 26180
rect 40292 26124 40302 26180
rect 18834 26012 18844 26068
rect 18900 26012 19684 26068
rect 19740 26012 19750 26068
rect 28578 26012 28588 26068
rect 28644 26012 30156 26068
rect 30212 26012 30716 26068
rect 30772 26012 30782 26068
rect 37426 26012 37436 26068
rect 37492 26012 39116 26068
rect 39172 26012 39182 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14886 25788 14924 25844
rect 14980 25788 14990 25844
rect 24098 25788 24108 25844
rect 24164 25788 24174 25844
rect 10658 25676 10668 25732
rect 10724 25676 18172 25732
rect 18228 25676 19180 25732
rect 19236 25676 19246 25732
rect 9990 25452 10000 25508
rect 10056 25452 10332 25508
rect 10388 25452 10398 25508
rect 14670 25452 14680 25508
rect 14736 25452 15148 25508
rect 15204 25452 19292 25508
rect 19348 25452 19358 25508
rect 22530 25452 22540 25508
rect 22596 25452 22988 25508
rect 23044 25452 23054 25508
rect 19618 25340 19628 25396
rect 19684 25340 20300 25396
rect 20356 25340 21420 25396
rect 21476 25340 21486 25396
rect 14466 25228 14476 25284
rect 14532 25228 14542 25284
rect 19170 25228 19180 25284
rect 19236 25228 19684 25284
rect 14476 25172 14532 25228
rect 19628 25172 19684 25228
rect 24108 25172 24164 25788
rect 28914 25676 28924 25732
rect 28980 25676 30828 25732
rect 30884 25676 30894 25732
rect 30574 25452 30584 25508
rect 30640 25452 32060 25508
rect 32116 25452 35532 25508
rect 35588 25452 35598 25508
rect 42802 25452 42812 25508
rect 42868 25452 43820 25508
rect 43876 25452 43886 25508
rect 25330 25340 25340 25396
rect 25396 25340 25844 25396
rect 25900 25340 32396 25396
rect 32452 25340 34300 25396
rect 34356 25340 34366 25396
rect 41234 25228 41244 25284
rect 41300 25228 41580 25284
rect 41636 25228 42644 25284
rect 42700 25228 42710 25284
rect 11890 25116 11900 25172
rect 11956 25116 13804 25172
rect 13860 25116 14532 25172
rect 16594 25116 16604 25172
rect 16660 25116 17948 25172
rect 18004 25116 18396 25172
rect 18452 25116 18462 25172
rect 19618 25116 19628 25172
rect 19684 25116 19694 25172
rect 24098 25116 24108 25172
rect 24164 25116 24174 25172
rect 5730 24892 5740 24948
rect 5796 24892 6748 24948
rect 6804 24892 9324 24948
rect 9380 24892 9390 24948
rect 14476 24836 14532 25116
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 20178 24892 20188 24948
rect 20244 24892 23436 24948
rect 23492 24892 23772 24948
rect 23828 24892 23838 24948
rect 14476 24780 14588 24836
rect 14644 24780 14654 24836
rect 4610 24668 4620 24724
rect 4676 24668 7084 24724
rect 7140 24668 9548 24724
rect 9604 24668 9614 24724
rect 14466 24668 14476 24724
rect 14532 24668 14700 24724
rect 14756 24668 15036 24724
rect 15092 24668 15102 24724
rect 15250 24668 15260 24724
rect 15316 24668 21868 24724
rect 21924 24668 22932 24724
rect 22988 24668 22998 24724
rect 39218 24668 39228 24724
rect 39284 24668 40124 24724
rect 40180 24668 40190 24724
rect 1922 24556 1932 24612
rect 1988 24556 5236 24612
rect 5292 24556 7980 24612
rect 8036 24556 8046 24612
rect 14578 24556 14588 24612
rect 14644 24556 14924 24612
rect 14980 24556 14990 24612
rect 25274 24444 25284 24500
rect 25340 24444 34412 24500
rect 34468 24444 35644 24500
rect 35700 24444 35710 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 4162 23996 4172 24052
rect 4228 23996 4620 24052
rect 4676 23996 4900 24052
rect 4956 23996 5516 24052
rect 5572 23996 5582 24052
rect 8978 23996 8988 24052
rect 9044 23996 15092 24052
rect 15148 23996 15158 24052
rect 10098 23884 10108 23940
rect 10164 23884 13748 23940
rect 13804 23884 13814 23940
rect 22922 23884 22932 23940
rect 22988 23884 23548 23940
rect 23604 23884 23614 23940
rect 36306 23884 36316 23940
rect 36372 23884 37100 23940
rect 37156 23884 37660 23940
rect 37716 23884 37726 23940
rect 15586 23660 15596 23716
rect 15652 23660 17388 23716
rect 17444 23660 17454 23716
rect 37986 23660 37996 23716
rect 38052 23660 39228 23716
rect 39284 23660 39294 23716
rect 5058 23548 5068 23604
rect 5124 23548 5740 23604
rect 5796 23548 5806 23604
rect 15250 23548 15260 23604
rect 15316 23548 15876 23604
rect 15932 23548 15942 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 35466 23436 35476 23492
rect 35532 23436 36092 23492
rect 36148 23436 36158 23492
rect 1698 23212 1708 23268
rect 1764 23212 21364 23268
rect 21420 23212 21644 23268
rect 21700 23212 21710 23268
rect 23258 23212 23268 23268
rect 23324 23212 23772 23268
rect 23828 23212 23838 23268
rect 30126 23100 30136 23156
rect 30192 23100 31948 23156
rect 32004 23100 32014 23156
rect 36698 22988 36708 23044
rect 36764 22988 37100 23044
rect 37156 22988 37166 23044
rect 34850 22876 34860 22932
rect 34916 22876 35980 22932
rect 36036 22876 36046 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 4274 22652 4284 22708
rect 4340 22652 4350 22708
rect 4284 22596 4340 22652
rect 4284 22540 5684 22596
rect 5740 22540 5750 22596
rect 10210 22540 10220 22596
rect 10276 22540 13580 22596
rect 13636 22540 18060 22596
rect 18116 22540 18620 22596
rect 18676 22540 18686 22596
rect 20066 22540 20076 22596
rect 20132 22540 36092 22596
rect 36148 22540 36158 22596
rect 3938 22428 3948 22484
rect 4004 22428 4620 22484
rect 4676 22428 4686 22484
rect 5058 22428 5068 22484
rect 5124 22428 6076 22484
rect 6132 22428 6142 22484
rect 12002 22428 12012 22484
rect 12068 22428 13692 22484
rect 13748 22428 15036 22484
rect 15092 22428 15102 22484
rect 16706 22428 16716 22484
rect 16772 22428 17948 22484
rect 18004 22428 18014 22484
rect 18946 22428 18956 22484
rect 19012 22428 20412 22484
rect 20468 22428 20478 22484
rect 31892 22428 34524 22484
rect 34580 22428 34590 22484
rect 31892 22372 31948 22428
rect 4834 22316 4844 22372
rect 4900 22316 5964 22372
rect 6020 22316 6030 22372
rect 7970 22316 7980 22372
rect 8036 22316 11284 22372
rect 11340 22316 11350 22372
rect 14914 22316 14924 22372
rect 14980 22316 15316 22372
rect 15372 22316 17724 22372
rect 17780 22316 17790 22372
rect 30238 22316 30248 22372
rect 30304 22316 31948 22372
rect 34270 22316 34280 22372
rect 34336 22316 35028 22372
rect 35084 22316 35980 22372
rect 36036 22316 36046 22372
rect 36362 22316 36372 22372
rect 36428 22316 39060 22372
rect 39116 22316 39126 22372
rect 6402 22204 6412 22260
rect 6468 22204 8428 22260
rect 14802 22204 14812 22260
rect 14868 22204 16100 22260
rect 16156 22204 16166 22260
rect 17546 22204 17556 22260
rect 17612 22204 18228 22260
rect 18284 22204 19460 22260
rect 19516 22204 19628 22260
rect 19684 22204 20076 22260
rect 20132 22204 20142 22260
rect 27346 22204 27356 22260
rect 27412 22204 28364 22260
rect 28420 22204 31276 22260
rect 31332 22204 31342 22260
rect 32181 22204 32191 22260
rect 32247 22204 34860 22260
rect 34916 22204 34926 22260
rect 8372 22148 8428 22204
rect 8372 22092 15202 22148
rect 15258 22092 16604 22148
rect 16660 22092 16670 22148
rect 13906 21980 13916 22036
rect 13972 21980 18396 22036
rect 18452 21980 18956 22036
rect 19012 21980 19022 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 15922 21868 15932 21924
rect 15988 21868 16716 21924
rect 16772 21868 16782 21924
rect 5394 21756 5404 21812
rect 5460 21756 10015 21812
rect 10071 21756 10081 21812
rect 28222 21756 28232 21812
rect 28288 21756 29036 21812
rect 29092 21756 29102 21812
rect 39442 21756 39452 21812
rect 39508 21756 39900 21812
rect 39956 21756 41244 21812
rect 41300 21756 41310 21812
rect 15474 21644 15484 21700
rect 15540 21644 16156 21700
rect 16212 21644 20972 21700
rect 21028 21644 21038 21700
rect 28802 21644 28812 21700
rect 28868 21644 31388 21700
rect 31444 21644 33292 21700
rect 33348 21644 33358 21700
rect 39330 21644 39340 21700
rect 39396 21644 40012 21700
rect 40068 21644 41356 21700
rect 41412 21644 41422 21700
rect 11890 21532 11900 21588
rect 11956 21532 12516 21588
rect 12572 21532 16660 21588
rect 16818 21532 16828 21588
rect 16884 21532 19292 21588
rect 19348 21532 20300 21588
rect 20356 21532 20366 21588
rect 33394 21532 33404 21588
rect 33460 21532 34524 21588
rect 34580 21532 34590 21588
rect 39554 21532 39564 21588
rect 39620 21532 40908 21588
rect 40964 21532 40974 21588
rect 16604 21476 16660 21532
rect 16604 21420 19068 21476
rect 19124 21420 19796 21476
rect 19852 21420 19862 21476
rect 39722 21308 39732 21364
rect 39788 21308 41244 21364
rect 41300 21308 42644 21364
rect 42700 21308 42710 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 29026 20972 29036 21028
rect 29092 20972 29540 21028
rect 29596 20972 29606 21028
rect 4610 20860 4620 20916
rect 4676 20860 5628 20916
rect 5684 20860 5694 20916
rect 9762 20748 9772 20804
rect 9828 20748 11564 20804
rect 11620 20748 11630 20804
rect 12002 20748 12012 20804
rect 12068 20748 13468 20804
rect 13524 20748 13534 20804
rect 24546 20748 24556 20804
rect 24612 20748 24948 20804
rect 25004 20748 25014 20804
rect 29250 20748 29260 20804
rect 29316 20748 32060 20804
rect 32116 20748 32126 20804
rect 9762 20524 9772 20580
rect 9828 20524 11340 20580
rect 11396 20524 11406 20580
rect 10994 20412 11004 20468
rect 11060 20412 11900 20468
rect 11956 20412 11966 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 36082 20300 36092 20356
rect 36148 20300 39116 20356
rect 39172 20300 40012 20356
rect 40068 20300 40078 20356
rect 32050 20188 32060 20244
rect 32116 20188 33404 20244
rect 33460 20188 33470 20244
rect 35970 20188 35980 20244
rect 36036 20188 38668 20244
rect 38724 20188 39900 20244
rect 39956 20188 39966 20244
rect 6066 20076 6076 20132
rect 6132 20076 6300 20132
rect 6356 20076 6366 20132
rect 12114 20076 12124 20132
rect 12180 20076 12628 20132
rect 12684 20076 21868 20132
rect 21924 20076 21934 20132
rect 27794 20076 27804 20132
rect 27860 20076 28700 20132
rect 28756 20076 28766 20132
rect 33114 20076 33124 20132
rect 33180 20076 35812 20132
rect 35868 20076 35878 20132
rect 37538 20076 37548 20132
rect 37604 20076 40572 20132
rect 40628 20076 40638 20132
rect 4274 19964 4284 20020
rect 4340 19964 5572 20020
rect 5628 19964 5638 20020
rect 6178 19964 6188 20020
rect 6244 19964 7196 20020
rect 7252 19964 7262 20020
rect 25106 19964 25116 20020
rect 25172 19964 29092 20020
rect 29148 19964 29158 20020
rect 35354 19964 35364 20020
rect 35420 19964 35644 20020
rect 35700 19964 35710 20020
rect 31042 19740 31052 19796
rect 31108 19740 33124 19796
rect 33180 19740 33190 19796
rect 32218 19628 32228 19684
rect 32284 19628 34972 19684
rect 35028 19628 35038 19684
rect 40226 19628 40236 19684
rect 40292 19628 40740 19684
rect 40796 19628 40806 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4834 19404 4844 19460
rect 4900 19404 5908 19460
rect 5964 19404 5974 19460
rect 7186 19404 7196 19460
rect 7252 19404 11004 19460
rect 11060 19404 11070 19460
rect 35522 19404 35532 19460
rect 35588 19404 39564 19460
rect 39620 19404 40908 19460
rect 40964 19404 41356 19460
rect 41412 19404 41422 19460
rect 4498 19292 4508 19348
rect 4564 19292 6300 19348
rect 6356 19292 6366 19348
rect 1810 19180 1820 19236
rect 1876 19180 5124 19236
rect 5180 19180 5190 19236
rect 5730 19180 5740 19236
rect 5796 19180 6692 19236
rect 6748 19180 9436 19236
rect 9492 19180 9502 19236
rect 17770 19180 17780 19236
rect 17836 19180 20860 19236
rect 20916 19180 20926 19236
rect 6402 18956 6412 19012
rect 6468 18956 6972 19012
rect 7028 18956 16324 19012
rect 16380 18956 16390 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 20850 18732 20860 18788
rect 20916 18732 21084 18788
rect 21140 18732 21150 18788
rect 28130 18620 28140 18676
rect 28196 18620 28364 18676
rect 28420 18620 28924 18676
rect 28980 18620 28990 18676
rect 10098 18508 10108 18564
rect 10164 18508 10388 18564
rect 10444 18508 14588 18564
rect 14644 18508 14654 18564
rect 26898 18508 26908 18564
rect 26964 18508 27692 18564
rect 27748 18508 27758 18564
rect 29036 18508 29148 18564
rect 29204 18508 29214 18564
rect 7634 18284 7644 18340
rect 7700 18284 14084 18340
rect 14140 18284 14150 18340
rect 14476 18228 14532 18508
rect 29036 18452 29092 18508
rect 14690 18396 14700 18452
rect 14756 18396 15204 18452
rect 15260 18396 15270 18452
rect 15586 18396 15596 18452
rect 15652 18396 16604 18452
rect 16660 18396 16670 18452
rect 27794 18396 27804 18452
rect 27860 18396 28756 18452
rect 28812 18396 29092 18452
rect 29250 18396 29260 18452
rect 29316 18396 30156 18452
rect 30212 18396 30222 18452
rect 35634 18396 35644 18452
rect 35700 18396 36092 18452
rect 36148 18396 36484 18452
rect 36540 18396 37548 18452
rect 37604 18396 37614 18452
rect 39340 18396 41020 18452
rect 41076 18396 43596 18452
rect 43652 18396 43662 18452
rect 15596 18340 15652 18396
rect 15026 18284 15036 18340
rect 15092 18284 15652 18340
rect 15754 18284 15764 18340
rect 15820 18284 16716 18340
rect 16772 18284 17388 18340
rect 17444 18284 17454 18340
rect 19954 18284 19964 18340
rect 20020 18284 21588 18340
rect 21644 18284 21654 18340
rect 24434 18284 24444 18340
rect 24500 18284 26180 18340
rect 26236 18284 26460 18340
rect 26516 18284 26526 18340
rect 27122 18284 27132 18340
rect 27188 18284 29428 18340
rect 29484 18284 29494 18340
rect 37314 18284 37324 18340
rect 37380 18284 39004 18340
rect 39060 18284 39070 18340
rect 29148 18228 29204 18284
rect 38668 18228 38724 18284
rect 39340 18228 39396 18396
rect 14476 18172 15652 18228
rect 20178 18172 20188 18228
rect 20244 18172 20972 18228
rect 21028 18172 21038 18228
rect 29138 18172 29148 18228
rect 29204 18172 29214 18228
rect 38658 18172 38668 18228
rect 38724 18172 38734 18228
rect 39330 18172 39340 18228
rect 39396 18172 39406 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 15596 17780 15652 18172
rect 28746 18060 28756 18116
rect 28812 18060 34076 18116
rect 34132 18060 34142 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 17826 17836 17836 17892
rect 17892 17836 20748 17892
rect 20804 17836 21364 17892
rect 21420 17836 21430 17892
rect 14466 17724 14476 17780
rect 14532 17724 15372 17780
rect 15428 17724 15438 17780
rect 15596 17724 24444 17780
rect 24500 17724 24510 17780
rect 14186 17612 14196 17668
rect 14252 17612 14700 17668
rect 14756 17612 15260 17668
rect 15316 17612 15326 17668
rect 20738 17612 20748 17668
rect 20804 17612 21868 17668
rect 21924 17612 22260 17668
rect 22316 17612 31836 17668
rect 31892 17612 33684 17668
rect 33740 17612 33750 17668
rect 17714 17388 17724 17444
rect 17780 17388 20860 17444
rect 20916 17388 27412 17444
rect 27468 17388 27804 17444
rect 27860 17388 27870 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 28018 17164 28028 17220
rect 28084 17164 29596 17220
rect 29652 17164 29662 17220
rect 21186 17052 21196 17108
rect 21252 17052 21700 17108
rect 21756 17052 21766 17108
rect 22194 17052 22204 17108
rect 22260 17052 31948 17108
rect 34178 17052 34188 17108
rect 34244 17052 36988 17108
rect 37044 17052 37054 17108
rect 31892 16996 31948 17052
rect 28466 16940 28476 16996
rect 28532 16940 29148 16996
rect 29204 16940 30156 16996
rect 30212 16940 30222 16996
rect 31892 16940 37100 16996
rect 37156 16940 37492 16996
rect 37548 16940 37558 16996
rect 20738 16828 20748 16884
rect 20804 16828 21756 16884
rect 21812 16828 21822 16884
rect 28354 16828 28364 16884
rect 28420 16828 29260 16884
rect 29316 16828 30044 16884
rect 30100 16828 30110 16884
rect 27458 16716 27468 16772
rect 27524 16716 28868 16772
rect 28924 16716 31164 16772
rect 31220 16716 31230 16772
rect 38322 16716 38332 16772
rect 38388 16716 38668 16772
rect 38724 16716 39340 16772
rect 39396 16716 39406 16772
rect 30930 16604 30940 16660
rect 30996 16604 32956 16660
rect 33012 16604 33022 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 21522 16268 21532 16324
rect 21588 16268 23884 16324
rect 23940 16268 23950 16324
rect 29026 16268 29036 16324
rect 29092 16268 30156 16324
rect 30212 16268 30222 16324
rect 22642 16156 22652 16212
rect 22708 16156 27860 16212
rect 27916 16156 29148 16212
rect 29204 16156 29214 16212
rect 16930 16044 16940 16100
rect 16996 16044 23044 16100
rect 23100 16044 23110 16100
rect 29138 15820 29148 15876
rect 29204 15820 33404 15876
rect 33460 15820 33470 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 37986 15596 37996 15652
rect 38052 15596 39004 15652
rect 39060 15596 39340 15652
rect 39396 15596 39406 15652
rect 15698 15484 15708 15540
rect 15764 15484 15774 15540
rect 29698 15484 29708 15540
rect 29764 15484 32508 15540
rect 32564 15484 32574 15540
rect 38770 15484 38780 15540
rect 38836 15484 39564 15540
rect 39620 15484 43820 15540
rect 43876 15484 43886 15540
rect 4498 15260 4508 15316
rect 4564 15260 5068 15316
rect 5124 15260 5516 15316
rect 5572 15260 7812 15316
rect 7868 15260 9436 15316
rect 9492 15260 10444 15316
rect 10500 15260 11004 15316
rect 11060 15260 11070 15316
rect 15708 15204 15764 15484
rect 29866 15372 29876 15428
rect 29932 15372 30940 15428
rect 30996 15372 31006 15428
rect 38322 15372 38332 15428
rect 38388 15372 39004 15428
rect 39060 15372 39070 15428
rect 23538 15260 23548 15316
rect 23604 15260 28588 15316
rect 28644 15260 28654 15316
rect 30426 15260 30436 15316
rect 30492 15260 31948 15316
rect 32004 15260 32014 15316
rect 34962 15260 34972 15316
rect 35028 15260 36316 15316
rect 36372 15260 38164 15316
rect 38220 15260 38230 15316
rect 38714 15260 38724 15316
rect 38780 15260 39822 15316
rect 39878 15260 39888 15316
rect 10322 15148 10332 15204
rect 10388 15148 12964 15204
rect 13020 15148 14700 15204
rect 14756 15148 14766 15204
rect 15026 15148 15036 15204
rect 15092 15148 16716 15204
rect 16772 15148 16782 15204
rect 28130 15148 28140 15204
rect 28196 15148 29036 15204
rect 29092 15148 29540 15204
rect 29596 15148 32732 15204
rect 32788 15148 32798 15204
rect 38434 15148 38444 15204
rect 38500 15148 38892 15204
rect 38948 15148 38958 15204
rect 40226 15036 40236 15092
rect 40292 15036 40460 15092
rect 40516 15036 40526 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 14130 14812 14140 14868
rect 14196 14812 15372 14868
rect 15428 14812 17500 14868
rect 17556 14812 17566 14868
rect 5282 14588 5292 14644
rect 5348 14588 5852 14644
rect 5908 14588 5918 14644
rect 14690 14588 14700 14644
rect 14756 14588 17332 14644
rect 17388 14588 22652 14644
rect 22708 14588 22718 14644
rect 25890 14588 25900 14644
rect 25956 14588 27020 14644
rect 27076 14588 27086 14644
rect 5954 14476 5964 14532
rect 6020 14476 6748 14532
rect 6804 14476 6814 14532
rect 12450 14476 12460 14532
rect 12516 14476 12908 14532
rect 12964 14476 13580 14532
rect 13636 14476 13646 14532
rect 24434 14476 24444 14532
rect 24500 14476 33796 14532
rect 33852 14476 34076 14532
rect 34132 14476 34142 14532
rect 40338 14476 40348 14532
rect 40404 14476 41132 14532
rect 41188 14476 41198 14532
rect 40348 14420 40404 14476
rect 36922 14364 36932 14420
rect 36988 14364 40404 14420
rect 19618 14252 19628 14308
rect 19684 14252 20356 14308
rect 20412 14252 24892 14308
rect 24948 14252 27244 14308
rect 27300 14252 27310 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 12114 13916 12124 13972
rect 12180 13916 12190 13972
rect 15642 13916 15652 13972
rect 15708 13916 20188 13972
rect 20244 13916 20254 13972
rect 12124 13860 12180 13916
rect 12124 13804 12572 13860
rect 12628 13804 13692 13860
rect 13748 13804 14476 13860
rect 14532 13804 14542 13860
rect 20290 13804 20300 13860
rect 20356 13804 21084 13860
rect 21140 13804 21150 13860
rect 13122 13692 13132 13748
rect 13188 13692 14028 13748
rect 14084 13692 14700 13748
rect 14756 13692 14766 13748
rect 20066 13692 20076 13748
rect 20132 13692 20524 13748
rect 20580 13692 21308 13748
rect 21364 13692 21374 13748
rect 21532 13692 21644 13748
rect 21700 13692 21710 13748
rect 33618 13692 33628 13748
rect 33684 13692 36932 13748
rect 36988 13692 36998 13748
rect 13850 13580 13860 13636
rect 13916 13580 14364 13636
rect 14420 13580 14532 13636
rect 14476 13524 14532 13580
rect 11330 13468 11340 13524
rect 11396 13468 14252 13524
rect 14308 13468 14318 13524
rect 14476 13468 15652 13524
rect 15708 13468 15718 13524
rect 12786 13356 12796 13412
rect 12852 13356 13468 13412
rect 13524 13356 13534 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 21532 13300 21588 13692
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 21522 13244 21532 13300
rect 21588 13244 21598 13300
rect 6962 13132 6972 13188
rect 7028 13132 7644 13188
rect 7700 13132 7710 13188
rect 8642 13020 8652 13076
rect 8708 13020 12236 13076
rect 12292 13020 12302 13076
rect 34178 13020 34188 13076
rect 34244 13020 38220 13076
rect 38276 13020 38286 13076
rect 7410 12908 7420 12964
rect 7476 12908 7868 12964
rect 7924 12908 8540 12964
rect 8596 12908 9324 12964
rect 9380 12908 9390 12964
rect 39218 12908 39228 12964
rect 39284 12908 39900 12964
rect 39956 12908 43708 12964
rect 43764 12908 43774 12964
rect 7420 12796 8204 12852
rect 8260 12796 8988 12852
rect 9044 12796 9054 12852
rect 7420 12740 7476 12796
rect 4946 12684 4956 12740
rect 5012 12684 7028 12740
rect 7084 12684 7476 12740
rect 7634 12684 7644 12740
rect 7700 12684 11564 12740
rect 11620 12684 12348 12740
rect 12404 12684 12414 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 2258 12124 2268 12180
rect 2324 12124 5516 12180
rect 5572 12124 5582 12180
rect 9426 12124 9436 12180
rect 9492 12124 13244 12180
rect 13300 12124 13310 12180
rect 13570 12124 13580 12180
rect 13636 12124 14812 12180
rect 14868 12124 14878 12180
rect 38322 12124 38332 12180
rect 38388 12124 39340 12180
rect 39396 12124 40012 12180
rect 40068 12124 40078 12180
rect 40562 12124 40572 12180
rect 40628 12124 41132 12180
rect 41188 12124 41198 12180
rect 19842 11788 19852 11844
rect 19908 11788 20524 11844
rect 20580 11788 20590 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 3042 11564 3052 11620
rect 3108 11564 3724 11620
rect 3780 11564 3790 11620
rect 12226 11452 12236 11508
rect 12292 11452 12908 11508
rect 12964 11452 12974 11508
rect 18162 11452 18172 11508
rect 18228 11452 19740 11508
rect 19796 11452 19806 11508
rect 4050 11340 4060 11396
rect 4116 11340 6860 11396
rect 6916 11340 6926 11396
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 25744 10780 25754 10836
rect 25810 10780 26516 10836
rect 26572 10780 29708 10836
rect 29764 10780 29774 10836
rect 21746 10668 21756 10724
rect 21812 10668 22484 10724
rect 22540 10668 22550 10724
rect 22194 10556 22204 10612
rect 22260 10556 23772 10612
rect 23828 10556 24444 10612
rect 24500 10556 24510 10612
rect 24602 10556 24612 10612
rect 24668 10556 26012 10612
rect 26068 10556 26684 10612
rect 26740 10556 26750 10612
rect 31470 10556 31480 10612
rect 31536 10556 32172 10612
rect 32228 10556 32956 10612
rect 33012 10556 33022 10612
rect 6738 10332 6748 10388
rect 6804 10332 9660 10388
rect 9716 10332 9726 10388
rect 27794 10332 27804 10388
rect 27860 10332 31724 10388
rect 31780 10332 31790 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 10434 10108 10444 10164
rect 10500 10108 11508 10164
rect 11564 10108 14364 10164
rect 14420 10108 14430 10164
rect 30146 10108 30156 10164
rect 30212 10108 30940 10164
rect 30996 10108 31006 10164
rect 7410 9996 7420 10052
rect 7476 9996 7980 10052
rect 8036 9996 8988 10052
rect 9044 9996 9054 10052
rect 4946 9884 4956 9940
rect 5012 9884 7084 9940
rect 7140 9884 13132 9940
rect 13188 9884 13468 9940
rect 13524 9884 13534 9940
rect 26562 9884 26572 9940
rect 26628 9884 27468 9940
rect 27524 9884 30548 9940
rect 30604 9884 30614 9940
rect 7410 9772 7420 9828
rect 7476 9772 8204 9828
rect 8260 9772 9100 9828
rect 9156 9772 10780 9828
rect 10836 9772 10846 9828
rect 25890 9772 25900 9828
rect 25956 9772 27020 9828
rect 27076 9772 27086 9828
rect 36194 9772 36204 9828
rect 36260 9772 36876 9828
rect 36932 9772 36942 9828
rect 7858 9660 7868 9716
rect 7924 9660 8708 9716
rect 8764 9660 9772 9716
rect 9828 9660 9838 9716
rect 24434 9660 24444 9716
rect 24500 9660 28588 9716
rect 28644 9660 32060 9716
rect 32116 9660 32126 9716
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 8978 9324 8988 9380
rect 9044 9324 10892 9380
rect 10948 9324 12348 9380
rect 12404 9324 12414 9380
rect 3042 9212 3052 9268
rect 3108 9212 4172 9268
rect 4228 9212 4238 9268
rect 11778 9212 11788 9268
rect 11844 9212 12460 9268
rect 12516 9212 13580 9268
rect 13636 9212 13646 9268
rect 20962 9212 20972 9268
rect 21028 9212 27412 9268
rect 27468 9212 27478 9268
rect 34066 9212 34076 9268
rect 34132 9212 35420 9268
rect 35476 9212 35486 9268
rect 10556 9100 12348 9156
rect 12404 9100 13300 9156
rect 13356 9100 13366 9156
rect 31892 9100 32396 9156
rect 32452 9100 33516 9156
rect 33572 9100 33582 9156
rect 10556 9044 10612 9100
rect 31892 9044 31948 9100
rect 4498 8988 4508 9044
rect 4564 8988 7308 9044
rect 7364 8988 7374 9044
rect 10098 8988 10108 9044
rect 10164 8988 10612 9044
rect 10668 8988 10678 9044
rect 10770 8988 10780 9044
rect 10836 8988 12124 9044
rect 12180 8988 12190 9044
rect 19170 8988 19180 9044
rect 19236 8988 19740 9044
rect 19796 8988 20188 9044
rect 20244 8988 21868 9044
rect 21924 8988 21934 9044
rect 25666 8988 25676 9044
rect 25732 8988 27132 9044
rect 27188 8988 27198 9044
rect 31378 8988 31388 9044
rect 31444 8988 31948 9044
rect 32162 8988 32172 9044
rect 32228 8988 33404 9044
rect 33460 8988 33470 9044
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 20794 8540 20804 8596
rect 20860 8540 27244 8596
rect 27300 8540 27310 8596
rect 19954 8428 19964 8484
rect 20020 8428 21028 8484
rect 19730 8316 19740 8372
rect 19796 8316 20804 8372
rect 20860 8316 20870 8372
rect 20972 8260 21028 8428
rect 24220 8428 25900 8484
rect 25956 8428 25966 8484
rect 24220 8372 24276 8428
rect 21634 8316 21644 8372
rect 21700 8316 24220 8372
rect 24276 8316 24286 8372
rect 9650 8204 9660 8260
rect 9716 8204 10668 8260
rect 10724 8204 10734 8260
rect 13458 8204 13468 8260
rect 13524 8204 13804 8260
rect 13860 8204 13870 8260
rect 20300 8204 22316 8260
rect 22372 8204 22382 8260
rect 20300 8036 20356 8204
rect 18386 7980 18396 8036
rect 18452 7980 19740 8036
rect 19796 7980 19806 8036
rect 20290 7980 20300 8036
rect 20356 7980 20366 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 7634 7532 7644 7588
rect 7700 7532 12572 7588
rect 12628 7532 14140 7588
rect 14196 7532 14206 7588
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 30818 6636 30828 6692
rect 30884 6636 31388 6692
rect 31444 6636 31454 6692
rect 20346 6412 20356 6468
rect 20412 6412 20972 6468
rect 21028 6412 21038 6468
rect 27122 6300 27132 6356
rect 27188 6300 27580 6356
rect 27636 6300 29596 6356
rect 29652 6300 29662 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 19730 6076 19740 6132
rect 19796 6076 20356 6132
rect 20412 6076 20422 6132
rect 27234 6076 27244 6132
rect 27300 6076 28252 6132
rect 28308 6076 30772 6132
rect 30828 6076 31052 6132
rect 31108 6076 31118 6132
rect 27906 5964 27916 6020
rect 27972 5964 29484 6020
rect 29540 5964 30940 6020
rect 30996 5964 31006 6020
rect 7746 5852 7756 5908
rect 7812 5852 9604 5908
rect 9660 5852 9670 5908
rect 9762 5852 9772 5908
rect 9828 5852 12012 5908
rect 12068 5852 12078 5908
rect 12450 5852 12460 5908
rect 12516 5852 13132 5908
rect 13188 5852 14028 5908
rect 14084 5852 14094 5908
rect 19954 5852 19964 5908
rect 20020 5852 20468 5908
rect 20524 5852 20534 5908
rect 22810 5852 22820 5908
rect 22876 5852 23548 5908
rect 23604 5852 23614 5908
rect 31826 5852 31836 5908
rect 31892 5852 32956 5908
rect 33012 5852 33022 5908
rect 9772 5796 9828 5852
rect 9202 5740 9212 5796
rect 9268 5740 9828 5796
rect 27458 5740 27468 5796
rect 27524 5740 28588 5796
rect 28644 5740 28654 5796
rect 28914 5740 28924 5796
rect 28980 5740 29876 5796
rect 29932 5740 31612 5796
rect 31668 5740 31678 5796
rect 8418 5628 8428 5684
rect 8484 5628 8932 5684
rect 8988 5628 8998 5684
rect 20402 5628 20412 5684
rect 20468 5628 21588 5684
rect 21644 5628 22540 5684
rect 22596 5628 22606 5684
rect 33282 5628 33292 5684
rect 33348 5628 34076 5684
rect 34132 5628 34142 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 8372 5180 9828 5236
rect 9884 5180 10108 5236
rect 10164 5180 13580 5236
rect 13636 5180 13646 5236
rect 13794 5180 13804 5236
rect 13860 5180 15932 5236
rect 15988 5180 15998 5236
rect 16706 5180 16716 5236
rect 16772 5180 17444 5236
rect 17500 5180 17510 5236
rect 20290 5180 20300 5236
rect 20356 5180 20860 5236
rect 20916 5180 20926 5236
rect 34850 5180 34860 5236
rect 34916 5180 35252 5236
rect 35308 5180 36204 5236
rect 36260 5180 36270 5236
rect 8372 5124 8428 5180
rect 5842 5068 5852 5124
rect 5908 5068 6524 5124
rect 6580 5068 8428 5124
rect 31266 5068 31276 5124
rect 31332 5068 32172 5124
rect 32228 5068 32238 5124
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 26282 4284 26292 4340
rect 26348 4284 26908 4340
rect 26964 4284 30212 4340
rect 30268 4284 30278 4340
rect 18386 4172 18396 4228
rect 18452 4172 19964 4228
rect 20020 4172 20030 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 18396 34300 18452 34356
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 18396 33068 18452 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 28476 31948 28532 32004
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 28476 30044 28532 30100
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 39788 27132 39844 27188
rect 39788 26908 39844 26964
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 14924 25788 14980 25844
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 14924 24556 14980 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 18396 34356 18452 34366
rect 18396 33124 18452 34300
rect 18396 33058 18452 33068
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 28476 32004 28532 32014
rect 28476 30100 28532 31948
rect 28476 30034 28532 30044
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 24332 4768 25844
rect 14924 25844 14980 25854
rect 14924 24612 14980 25788
rect 14924 24546 14980 24556
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 39788 27188 39844 27198
rect 39788 26964 39844 27132
rect 39788 26898 39844 26908
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_as_sc_mcu7t3v3__buff_2  _367_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform -1 0 22064 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _368_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 25760 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _369_
timestamp 1751534193
transform 1 0 10304 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _370_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform 1 0 9408 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _371_
timestamp 1751534193
transform -1 0 11984 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _372_
timestamp 1751905124
transform 1 0 9968 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _373_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform -1 0 10976 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _374_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform -1 0 10752 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _375_
timestamp 1753277515
transform -1 0 7616 0 1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _376_
timestamp 1753277515
transform -1 0 7952 0 1 31360
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _377_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform 1 0 7616 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _378_
timestamp 1751534193
transform -1 0 7168 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _379_
timestamp 1751905124
transform -1 0 10192 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _380_
timestamp 1751905124
transform 1 0 9856 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _381_
timestamp 1753277515
transform -1 0 10080 0 1 39200
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _382_
timestamp 1752345181
transform 1 0 10752 0 1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _383_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform 1 0 9856 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _384_
timestamp 1753277515
transform -1 0 11088 0 -1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _385_
timestamp 1753277515
transform -1 0 12320 0 -1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _386_
timestamp 1751531619
transform 1 0 11424 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _387_
timestamp 1751532043
transform -1 0 13216 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _388_
timestamp 1753182340
transform 1 0 11872 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _389_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform 1 0 8848 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _390_
timestamp 1751740063
transform 1 0 14560 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _391_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753172561
transform 1 0 12432 0 -1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _392_
timestamp 1751740063
transform 1 0 13328 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _393_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform 1 0 30688 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _394_
timestamp 1753182340
transform 1 0 30800 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _395_
timestamp 1751889808
transform 1 0 20272 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _396_
timestamp 1751889808
transform 1 0 21952 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _397_
timestamp 1751889808
transform 1 0 21616 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _398_
timestamp 1753182340
transform 1 0 21168 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _399_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform -1 0 21952 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _400_
timestamp 1751532043
transform -1 0 15568 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _401_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform 1 0 11536 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _402_
timestamp 1751534193
transform 1 0 11536 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _403_
timestamp 1751740063
transform 1 0 13440 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _404_
timestamp 1751534193
transform 1 0 13440 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _405_
timestamp 1752061876
transform 1 0 13216 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _406_
timestamp 1751740063
transform 1 0 14224 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _407_
timestamp 1753172561
transform 1 0 13552 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _408_
timestamp 1751889408
transform 1 0 17696 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _409_
timestamp 1753172561
transform 1 0 18480 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _410_
timestamp 1751534193
transform 1 0 26880 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _411_
timestamp 1751534193
transform 1 0 28000 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _412_
timestamp 1751532043
transform -1 0 33376 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _413_
timestamp 1753277515
transform 1 0 30016 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _414_
timestamp 1751889408
transform 1 0 29008 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _415_
timestamp 1753277515
transform 1 0 27216 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__maj3_2  _416_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753272495
transform 1 0 28448 0 -1 21952
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _417_
timestamp 1753277515
transform -1 0 33264 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _418_
timestamp 1753277515
transform 1 0 29120 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _419_
timestamp 1751531619
transform -1 0 28784 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _420_
timestamp 1751532043
transform 1 0 34832 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _421_
timestamp 1753277515
transform 1 0 33264 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _422_
timestamp 1753277515
transform 1 0 29232 0 1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _423_
timestamp 1751534193
transform -1 0 28784 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _424_
timestamp 1751532043
transform 1 0 32032 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _425_
timestamp 1753277515
transform 1 0 29568 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _426_
timestamp 1752345181
transform 1 0 28112 0 -1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _427_
timestamp 1752061876
transform 1 0 26320 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_4  _428_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753864693
transform 1 0 26320 0 -1 31360
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _429_
timestamp 1751889408
transform 1 0 23408 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _430_
timestamp 1751534193
transform 1 0 24192 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _431_
timestamp 1751889408
transform 1 0 18032 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _432_
timestamp 1751889408
transform -1 0 20384 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _433_
timestamp 1751534193
transform -1 0 34608 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _434_
timestamp 1753277515
transform 1 0 29344 0 -1 26656
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _435_
timestamp 1751531619
transform 1 0 28784 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _436_
timestamp 1753172561
transform 1 0 25424 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _437_
timestamp 1751531619
transform -1 0 30016 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _438_
timestamp 1751531619
transform 1 0 27440 0 -1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _439_
timestamp 1751531619
transform -1 0 30352 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _440_
timestamp 1752345181
transform -1 0 30464 0 1 26656
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _441_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform 1 0 29008 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _442_
timestamp 1751532043
transform 1 0 22288 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _443_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform -1 0 31024 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _444_
timestamp 1751531619
transform 1 0 29680 0 -1 36064
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _445_
timestamp 1751889808
transform 1 0 29008 0 1 37632
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _446_
timestamp 1751534193
transform 1 0 23296 0 -1 34496
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _447_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform -1 0 26096 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _448_
timestamp 1751534193
transform 1 0 29792 0 1 37632
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _449_
timestamp 1753371985
transform -1 0 25872 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _450_
timestamp 1753441877
transform -1 0 24304 0 1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _451_
timestamp 1751534193
transform -1 0 14336 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _452_
timestamp 1751534193
transform 1 0 21616 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _453_
timestamp 1751534193
transform 1 0 20272 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _454_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform 1 0 26432 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _455_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753579406
transform 1 0 27216 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _456_
timestamp 1753182340
transform -1 0 28672 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _457_
timestamp 1753441877
transform -1 0 24640 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _458_
timestamp 1751534193
transform 1 0 24080 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _459_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform 1 0 25312 0 -1 37632
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _460_
timestamp 1751740063
transform 1 0 28224 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _461_
timestamp 1751889808
transform 1 0 29008 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _462_
timestamp 1751534193
transform 1 0 29904 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _463_
timestamp 1751532043
transform 1 0 26656 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _464_
timestamp 1753441877
transform 1 0 28560 0 -1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _465_
timestamp 1751534193
transform 1 0 32480 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _466_
timestamp 1753172561
transform 1 0 29008 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _467_
timestamp 1751534193
transform -1 0 20608 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _468_
timestamp 1751531619
transform -1 0 24080 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _469_
timestamp 1751534193
transform 1 0 32480 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _470_
timestamp 1751534193
transform -1 0 34832 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _471_
timestamp 1751534193
transform -1 0 25312 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _472_
timestamp 1751740063
transform -1 0 20272 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _473_
timestamp 1751889408
transform 1 0 21056 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _474_
timestamp 1751534193
transform 1 0 23184 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _475_
timestamp 1751534193
transform 1 0 23520 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _476_
timestamp 1751531619
transform -1 0 21168 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _477_
timestamp 1751740063
transform -1 0 20384 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _478_
timestamp 1751740063
transform 1 0 19488 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _479_
timestamp 1751889408
transform 1 0 20048 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _480_
timestamp 1753182340
transform 1 0 19488 0 1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _481_
timestamp 1751534193
transform -1 0 18480 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _482_
timestamp 1751889408
transform 1 0 21056 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _483_
timestamp 1751889808
transform -1 0 21056 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _484_
timestamp 1751531619
transform 1 0 19488 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _485_
timestamp 1751740063
transform -1 0 20608 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _486_
timestamp 1751889808
transform 1 0 22288 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _487_
timestamp 1753172561
transform 1 0 21168 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _488_
timestamp 1751889408
transform -1 0 24528 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _489_
timestamp 1751889408
transform 1 0 23520 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _490_
timestamp 1751534193
transform 1 0 23856 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _491_
timestamp 1751532043
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _492_
timestamp 1751740063
transform 1 0 26544 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _493_
timestamp 1751534193
transform 1 0 33936 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _494_
timestamp 1753441877
transform -1 0 26208 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _495_
timestamp 1751740063
transform -1 0 25872 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _496_
timestamp 1751740063
transform -1 0 28112 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _497_
timestamp 1751889408
transform 1 0 29344 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _498_
timestamp 1753182340
transform 1 0 28112 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _499_
timestamp 1751534193
transform -1 0 28560 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _500_
timestamp 1751740063
transform 1 0 31024 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _501_
timestamp 1751889408
transform 1 0 31472 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _502_
timestamp 1753182340
transform 1 0 30912 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _503_
timestamp 1751534193
transform 1 0 32928 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _504_
timestamp 1751531619
transform -1 0 32704 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _505_
timestamp 1751889808
transform -1 0 33712 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _506_
timestamp 1751889408
transform 1 0 32032 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _507_
timestamp 1751889408
transform 1 0 32928 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _508_
timestamp 1751534193
transform 1 0 33712 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _509_
timestamp 1753277515
transform 1 0 30464 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _510_
timestamp 1751889408
transform 1 0 27552 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _511_
timestamp 1751534193
transform 1 0 27888 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _512_
timestamp 1751534193
transform 1 0 33824 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _513_
timestamp 1751534193
transform 1 0 21840 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _514_
timestamp 1751531619
transform 1 0 36848 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _515_
timestamp 1751534193
transform 1 0 37632 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _516_
timestamp 1751534193
transform 1 0 39200 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _517_
timestamp 1751534193
transform 1 0 36960 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _518_
timestamp 1751534193
transform -1 0 39088 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _519_
timestamp 1751534193
transform 1 0 37632 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _520_
timestamp 1751534193
transform 1 0 39088 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _521_
timestamp 1753960525
transform 1 0 35504 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _522_
timestamp 1753371985
transform 1 0 34832 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _523_
timestamp 1751534193
transform -1 0 39536 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _524_
timestamp 1751534193
transform -1 0 36960 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _525_
timestamp 1751534193
transform 1 0 36736 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _526_
timestamp 1753960525
transform 1 0 35280 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _527_
timestamp 1753441877
transform -1 0 35280 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _528_
timestamp 1751534193
transform -1 0 33712 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _529_
timestamp 1751532043
transform -1 0 40096 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _530_
timestamp 1751534193
transform 1 0 22400 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _531_
timestamp 1751534193
transform 1 0 38080 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _532_
timestamp 1753960525
transform -1 0 39984 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _533_
timestamp 1753371985
transform 1 0 35392 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _534_
timestamp 1751534193
transform 1 0 37072 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _535_
timestamp 1753960525
transform 1 0 38976 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _536_
timestamp 1753441877
transform 1 0 39088 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _537_
timestamp 1751534193
transform 1 0 40656 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _538_
timestamp 1751534193
transform -1 0 39648 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _539_
timestamp 1753960525
transform 1 0 37856 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _540_
timestamp 1753441877
transform 1 0 39424 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _541_
timestamp 1751534193
transform 1 0 40432 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _542_
timestamp 1751534193
transform -1 0 24864 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _543_
timestamp 1751740063
transform -1 0 38864 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _544_
timestamp 1751534193
transform -1 0 17920 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _545_
timestamp 1751534193
transform 1 0 17360 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _546_
timestamp 1751740063
transform -1 0 35168 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _547_
timestamp 1753182340
transform 1 0 33936 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _548_
timestamp 1751534193
transform 1 0 34272 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _549_
timestamp 1753960525
transform -1 0 39536 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _550_
timestamp 1753441877
transform -1 0 39648 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _551_
timestamp 1751534193
transform -1 0 38976 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _552_
timestamp 1753960525
transform 1 0 38864 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _553_
timestamp 1753441877
transform 1 0 39760 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _554_
timestamp 1751534193
transform 1 0 41104 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _555_
timestamp 1751532043
transform 1 0 40992 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _556_
timestamp 1751532043
transform -1 0 42896 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _557_
timestamp 1753960525
transform 1 0 39424 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _558_
timestamp 1753371985
transform -1 0 41776 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _559_
timestamp 1751532043
transform -1 0 42896 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _560_
timestamp 1753960525
transform 1 0 40768 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _561_
timestamp 1753371985
transform 1 0 40656 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _562_
timestamp 1751534193
transform 1 0 40096 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _563_
timestamp 1751534193
transform 1 0 36848 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _564_
timestamp 1751534193
transform 1 0 37520 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _565_
timestamp 1753277515
transform 1 0 40208 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _566_
timestamp 1753960525
transform 1 0 40768 0 -1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _567_
timestamp 1753371985
transform 1 0 40992 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _568_
timestamp 1751532043
transform -1 0 42224 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _569_
timestamp 1751532043
transform -1 0 42896 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _570_
timestamp 1751534193
transform 1 0 37296 0 -1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _571_
timestamp 1753960525
transform 1 0 40768 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _572_
timestamp 1753371985
transform 1 0 41104 0 1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _573_
timestamp 1753277515
transform 1 0 38976 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _574_
timestamp 1753960525
transform 1 0 39536 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _575_
timestamp 1753371985
transform -1 0 42000 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _576_
timestamp 1751532043
transform -1 0 41216 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _577_
timestamp 1753277515
transform 1 0 36960 0 -1 36064
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _578_
timestamp 1753960525
transform 1 0 38304 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _579_
timestamp 1753371985
transform -1 0 40992 0 1 36064
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _580_
timestamp 1751532043
transform -1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _581_
timestamp 1751532043
transform 1 0 36848 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _582_
timestamp 1753960525
transform -1 0 37296 0 -1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _583_
timestamp 1753371985
transform 1 0 35280 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _584_
timestamp 1753960525
transform 1 0 35056 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _585_
timestamp 1753371985
transform -1 0 36848 0 -1 31360
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _586_
timestamp 1751531619
transform 1 0 13440 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _587_
timestamp 1751534193
transform 1 0 10640 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _588_
timestamp 1753371985
transform -1 0 12208 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _589_
timestamp 1751534193
transform 1 0 15232 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _590_
timestamp 1751889808
transform -1 0 16240 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _591_
timestamp 1751889408
transform -1 0 16912 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _592_
timestamp 1751889408
transform -1 0 7280 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _593_
timestamp 1753182340
transform -1 0 10304 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _594_
timestamp 1751534193
transform -1 0 10080 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _595_
timestamp 1751531619
transform -1 0 17024 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _596_
timestamp 1753441877
transform 1 0 14784 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _597_
timestamp 1751534193
transform 1 0 16240 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _598_
timestamp 1751531619
transform -1 0 16800 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _599_
timestamp 1751740063
transform -1 0 6272 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _600_
timestamp 1751889408
transform -1 0 6496 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _601_
timestamp 1751889408
transform -1 0 6496 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _602_
timestamp 1753182340
transform 1 0 4032 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _603_
timestamp 1751534193
transform -1 0 3584 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _604_
timestamp 1751889408
transform -1 0 6272 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _605_
timestamp 1751740063
transform -1 0 5264 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _606_
timestamp 1753182340
transform -1 0 4816 0 -1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _607_
timestamp 1751534193
transform -1 0 3584 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _608_
timestamp 1751889408
transform -1 0 16688 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _609_
timestamp 1751534193
transform -1 0 15120 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _610_
timestamp 1753182340
transform 1 0 17248 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _611_
timestamp 1753579406
transform -1 0 5376 0 -1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _612_
timestamp 1753172561
transform 1 0 5152 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _613_
timestamp 1751740063
transform -1 0 6496 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _614_
timestamp 1751740063
transform -1 0 4256 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _615_
timestamp 1751534193
transform -1 0 8848 0 1 32928
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _616_
timestamp 1751740063
transform 1 0 5488 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _617_
timestamp 1751889408
transform 1 0 5488 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _618_
timestamp 1753182340
transform -1 0 6720 0 1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _619_
timestamp 1751534193
transform 1 0 6272 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _620_
timestamp 1753579406
transform 1 0 4032 0 -1 32928
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _621_
timestamp 1751889408
transform 1 0 4704 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _622_
timestamp 1751889408
transform 1 0 6272 0 1 32928
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _623_
timestamp 1751740063
transform -1 0 3808 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _624_
timestamp 1751534193
transform -1 0 8176 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _625_
timestamp 1753441877
transform -1 0 4816 0 1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _626_
timestamp 1751740063
transform -1 0 5600 0 -1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _627_
timestamp 1751740063
transform 1 0 4480 0 1 39200
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _628_
timestamp 1751905124
transform -1 0 4816 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _629_
timestamp 1753371985
transform 1 0 3696 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _630_
timestamp 1753371985
transform -1 0 3696 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _631_
timestamp 1752345181
transform 1 0 5712 0 -1 32928
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _632_
timestamp 1751740063
transform 1 0 5936 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _633_
timestamp 1751889408
transform 1 0 6720 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _634_
timestamp 1753172561
transform -1 0 15904 0 1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _635_
timestamp 1753960525
transform -1 0 16128 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _636_
timestamp 1751889408
transform -1 0 15008 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _637_
timestamp 1751889408
transform 1 0 14448 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _638_
timestamp 1751534193
transform 1 0 14896 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _639_
timestamp 1751532043
transform -1 0 13776 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _640_
timestamp 1751740063
transform -1 0 12656 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _641_
timestamp 1753960525
transform -1 0 21392 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _642_
timestamp 1753441877
transform 1 0 13440 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _643_
timestamp 1751740063
transform -1 0 11872 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _644_
timestamp 1751534193
transform -1 0 10080 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _645_
timestamp 1753277515
transform -1 0 8064 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _646_
timestamp 1751740063
transform -1 0 6496 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _647_
timestamp 1753371985
transform -1 0 8064 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _648_
timestamp 1751531619
transform 1 0 8064 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _649_
timestamp 1753182340
transform -1 0 13104 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _650_
timestamp 1751534193
transform -1 0 12768 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _651_
timestamp 1753182340
transform 1 0 6608 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _652_
timestamp 1751534193
transform -1 0 4144 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _653_
timestamp 1751534193
transform 1 0 7056 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _654_
timestamp 1751740063
transform -1 0 8512 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _655_
timestamp 1751889408
transform -1 0 9296 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _656_
timestamp 1753182340
transform 1 0 7056 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _657_
timestamp 1751534193
transform -1 0 4592 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _658_
timestamp 1751534193
transform -1 0 13104 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _659_
timestamp 1751740063
transform -1 0 10304 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _660_
timestamp 1753960525
transform 1 0 10304 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _661_
timestamp 1751740063
transform 1 0 10528 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _662_
timestamp 1753172561
transform -1 0 12992 0 -1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _663_
timestamp 1753960525
transform 1 0 12992 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _664_
timestamp 1752061876
transform 1 0 13328 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _665_
timestamp 1751889408
transform 1 0 14112 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _666_
timestamp 1751534193
transform -1 0 14224 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _667_
timestamp 1751532043
transform -1 0 9856 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _668_
timestamp 1751889808
transform 1 0 7616 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _669_
timestamp 1753371985
transform 1 0 7392 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _670_
timestamp 1751889408
transform 1 0 8400 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _671_
timestamp 1751534193
transform -1 0 7952 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _672_
timestamp 1751534193
transform 1 0 23072 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _673_
timestamp 1751532043
transform 1 0 23744 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _674_
timestamp 1751534193
transform 1 0 17920 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _675_
timestamp 1751889808
transform -1 0 23856 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _676_
timestamp 1753371985
transform 1 0 23856 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _677_
timestamp 1751889408
transform 1 0 23744 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _678_
timestamp 1751534193
transform -1 0 23856 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _679_
timestamp 1751534193
transform -1 0 21840 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _680_
timestamp 1751532043
transform 1 0 22512 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _681_
timestamp 1753277515
transform 1 0 22848 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _682_
timestamp 1753960525
transform -1 0 25536 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _683_
timestamp 1753371985
transform 1 0 22736 0 1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _684_
timestamp 1751889408
transform -1 0 18816 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _685_
timestamp 1752345181
transform 1 0 19040 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _686_
timestamp 1753441877
transform -1 0 20384 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _687_
timestamp 1751889408
transform 1 0 18144 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _688_
timestamp 1753960525
transform 1 0 18816 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _689_
timestamp 1751889408
transform 1 0 19824 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _690_
timestamp 1751534193
transform 1 0 20608 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _691_
timestamp 1753277515
transform 1 0 13664 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _692_
timestamp 1751740063
transform -1 0 20608 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _693_
timestamp 1753868718
transform -1 0 14784 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _694_
timestamp 1751534193
transform -1 0 10192 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _695_
timestamp 1752061876
transform 1 0 14448 0 -1 26656
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _696_
timestamp 1751889408
transform 1 0 16128 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _697_
timestamp 1751534193
transform 1 0 17136 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _698_
timestamp 1751740063
transform -1 0 19376 0 -1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _699_
timestamp 1753371985
transform 1 0 16128 0 1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _700_
timestamp 1751740063
transform 1 0 15120 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _701_
timestamp 1753182340
transform 1 0 14784 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _702_
timestamp 1751534193
transform -1 0 12544 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _703_
timestamp 1751534193
transform 1 0 18368 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _704_
timestamp 1751889808
transform 1 0 18368 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _705_
timestamp 1751531619
transform -1 0 19936 0 -1 34496
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _706_
timestamp 1753441877
transform 1 0 18032 0 1 32928
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _707_
timestamp 1753960525
transform 1 0 18368 0 1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _708_
timestamp 1751534193
transform 1 0 19152 0 1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _709_
timestamp 1751534193
transform 1 0 14336 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _710_
timestamp 1753277515
transform -1 0 15456 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _711_
timestamp 1753868718
transform -1 0 14896 0 -1 34496
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _712_
timestamp 1751534193
transform -1 0 12096 0 -1 36064
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _713_
timestamp 1753960525
transform 1 0 15904 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _714_
timestamp 1753172561
transform 1 0 16464 0 1 34496
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _715_
timestamp 1753960525
transform -1 0 18368 0 -1 34496
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _716_
timestamp 1753441877
transform 1 0 17248 0 -1 37632
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _717_
timestamp 1751534193
transform -1 0 16464 0 -1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _718_
timestamp 1751740063
transform -1 0 28336 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _719_
timestamp 1751889408
transform 1 0 28896 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _720_
timestamp 1753182340
transform 1 0 26320 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _721_
timestamp 1751534193
transform -1 0 26320 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _722_
timestamp 1751889408
transform -1 0 29456 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _723_
timestamp 1751889808
transform 1 0 28000 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _724_
timestamp 1751531619
transform -1 0 28896 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _725_
timestamp 1751740063
transform -1 0 27664 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _726_
timestamp 1751740063
transform 1 0 30688 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _727_
timestamp 1753960525
transform 1 0 29568 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _728_
timestamp 1751740063
transform 1 0 31472 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _729_
timestamp 1751889808
transform -1 0 36400 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _730_
timestamp 1751740063
transform 1 0 18928 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _731_
timestamp 1753441877
transform 1 0 20608 0 -1 29792
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _732_
timestamp 1753441877
transform 1 0 35952 0 -1 39200
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _733_
timestamp 1751534193
transform 1 0 36848 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _734_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751632746
transform 1 0 18368 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _735_
timestamp 1751632746
transform -1 0 14560 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _736_
timestamp 1751632746
transform 1 0 21840 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _737_
timestamp 1751632746
transform 1 0 25984 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _738_
timestamp 1751632746
transform 1 0 29680 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _739_
timestamp 1751632746
transform 1 0 33264 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _740_
timestamp 1751632746
transform -1 0 18592 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _741_
timestamp 1751632746
transform 1 0 17696 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _742_
timestamp 1751632746
transform 1 0 17360 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _743_
timestamp 1751632746
transform 1 0 16464 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _744_
timestamp 1751632746
transform 1 0 17584 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _745_
timestamp 1751632746
transform -1 0 25984 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _746_
timestamp 1751632746
transform -1 0 26544 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _747_
timestamp 1751632746
transform 1 0 26880 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _748_
timestamp 1751632746
transform -1 0 34944 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _749_
timestamp 1751632746
transform -1 0 36288 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _750_
timestamp 1751632746
transform 1 0 27440 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _751_
timestamp 1751632746
transform -1 0 33824 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _752_
timestamp 1751632746
transform 1 0 28560 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _753_
timestamp 1751632746
transform 1 0 21840 0 -1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _754_
timestamp 1751632746
transform -1 0 36176 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _755_
timestamp 1751632746
transform -1 0 34160 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _756_
timestamp 1751632746
transform -1 0 37632 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _757_
timestamp 1751632746
transform 1 0 40768 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _758_
timestamp 1751632746
transform 1 0 41104 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _759_
timestamp 1751632746
transform 1 0 33600 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _760_
timestamp 1751632746
transform 1 0 36848 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _761_
timestamp 1751632746
transform 1 0 40992 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _762_
timestamp 1751632746
transform 1 0 40880 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _763_
timestamp 1751632746
transform 1 0 40880 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _764_
timestamp 1751632746
transform 1 0 41104 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _765_
timestamp 1751632746
transform 1 0 41104 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _766_
timestamp 1751632746
transform 1 0 41104 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _767_
timestamp 1751632746
transform 1 0 39648 0 1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _768_
timestamp 1751632746
transform 1 0 33936 0 -1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _769_
timestamp 1751632746
transform 1 0 33600 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _770_
timestamp 1751632746
transform 1 0 7952 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _771_
timestamp 1751632746
transform 1 0 1792 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _772_
timestamp 1751632746
transform 1 0 1904 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _773_
timestamp 1751632746
transform 1 0 1792 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _774_
timestamp 1751632746
transform 1 0 6496 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _775_
timestamp 1751632746
transform 1 0 1792 0 1 32928
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _776_
timestamp 1751632746
transform 1 0 5712 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _777_
timestamp 1751632746
transform 1 0 2128 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _778_
timestamp 1751632746
transform 1 0 14000 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _779_
timestamp 1751632746
transform 1 0 10416 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _780_
timestamp 1751632746
transform 1 0 4480 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _781_
timestamp 1751632746
transform 1 0 2240 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _782_
timestamp 1751632746
transform 1 0 2240 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _783_
timestamp 1751632746
transform 1 0 10080 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _784_
timestamp 1751632746
transform -1 0 16800 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _785_
timestamp 1751632746
transform 1 0 6496 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _786_
timestamp 1751632746
transform -1 0 24640 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _787_
timestamp 1751632746
transform -1 0 24752 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _788_
timestamp 1751632746
transform -1 0 20944 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _789_
timestamp 1751632746
transform 1 0 7952 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _790_
timestamp 1751632746
transform -1 0 12656 0 1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _791_
timestamp 1751632746
transform -1 0 21392 0 -1 37632
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _792_
timestamp 1751632746
transform -1 0 12880 0 1 36064
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _793_
timestamp 1751632746
transform -1 0 13104 0 1 39200
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _794_
timestamp 1751632746
transform 1 0 25088 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _795_
timestamp 1751632746
transform 1 0 25088 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _796_
timestamp 1751632746
transform -1 0 32816 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _797_
timestamp 1751632746
transform 1 0 36288 0 -1 40768
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _798_
timestamp 1751534193
transform 1 0 39312 0 -1 40768
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _799_
timestamp 1751534193
transform -1 0 43008 0 1 39200
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__367__A dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform 1 0 21168 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__385__A
timestamp 1751532392
transform 1 0 12544 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__399__A
timestamp 1751532392
transform -1 0 22400 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__400__A
timestamp 1751532392
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__406__B
timestamp 1751532392
transform 1 0 15232 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__409__D
timestamp 1751532392
transform -1 0 17696 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__429__A
timestamp 1751532392
transform 1 0 23184 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__432__B
timestamp 1751532392
transform 1 0 19376 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__434__B
timestamp 1751532392
transform 1 0 31136 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__436__B
timestamp 1751532392
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__442__A
timestamp 1751532392
transform 1 0 22960 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__447__C
timestamp 1751532392
transform -1 0 24976 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__452__A
timestamp 1751532392
transform 1 0 22512 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__456__A
timestamp 1751532392
transform -1 0 27440 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__471__A
timestamp 1751532392
transform -1 0 25760 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__472__B
timestamp 1751532392
transform 1 0 20272 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__474__A
timestamp 1751532392
transform -1 0 23184 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__476__A
timestamp 1751532392
transform 1 0 21392 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__480__A
timestamp 1751532392
transform 1 0 20720 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__484__A
timestamp 1751532392
transform 1 0 20272 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__494__C
timestamp 1751532392
transform -1 0 26656 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__498__A
timestamp 1751532392
transform -1 0 27328 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__502__A
timestamp 1751532392
transform -1 0 30912 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__510__A
timestamp 1751532392
transform 1 0 27328 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__512__A
timestamp 1751532392
transform 1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__514__B
timestamp 1751532392
transform 1 0 36624 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__519__A
timestamp 1751532392
transform 1 0 37408 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__521__D
timestamp 1751532392
transform 1 0 35280 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__525__A
timestamp 1751532392
transform -1 0 36736 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__526__D
timestamp 1751532392
transform -1 0 35280 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__529__A
timestamp 1751532392
transform -1 0 40544 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__530__A
timestamp 1751532392
transform 1 0 23296 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__531__A
timestamp 1751532392
transform 1 0 37856 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__536__A
timestamp 1751532392
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__542__A
timestamp 1751532392
transform 1 0 24864 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__546__B
timestamp 1751532392
transform 1 0 34160 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__547__A
timestamp 1751532392
transform -1 0 33936 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__564__A
timestamp 1751532392
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__565__A
timestamp 1751532392
transform 1 0 39984 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__573__A
timestamp 1751532392
transform -1 0 38976 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__577__A
timestamp 1751532392
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__584__D
timestamp 1751532392
transform 1 0 34832 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__588__B
timestamp 1751532392
transform 1 0 12432 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__589__A
timestamp 1751532392
transform 1 0 15008 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__593__A
timestamp 1751532392
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__598__A
timestamp 1751532392
transform 1 0 17472 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__602__A
timestamp 1751532392
transform -1 0 5712 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__606__A
timestamp 1751532392
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__608__A
timestamp 1751532392
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__610__B
timestamp 1751532392
transform 1 0 18704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__611__B
timestamp 1751532392
transform 1 0 6048 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__611__D
timestamp 1751532392
transform -1 0 5824 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__618__A
timestamp 1751532392
transform 1 0 6944 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__620__B
timestamp 1751532392
transform 1 0 7168 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__620__C
timestamp 1751532392
transform 1 0 5824 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__625__C
timestamp 1751532392
transform -1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__628__B
timestamp 1751532392
transform -1 0 5264 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__634__D
timestamp 1751532392
transform -1 0 14336 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__635__C
timestamp 1751532392
transform 1 0 14000 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__641__B
timestamp 1751532392
transform 1 0 21392 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__641__D
timestamp 1751532392
transform 1 0 21616 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__642__C
timestamp 1751532392
transform 1 0 15568 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__644__A
timestamp 1751532392
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__660__D
timestamp 1751532392
transform 1 0 11424 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__664__B
timestamp 1751532392
transform -1 0 14896 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__672__A
timestamp 1751532392
transform 1 0 22848 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__675__B
timestamp 1751532392
transform -1 0 23072 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__676__C
timestamp 1751532392
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__682__B
timestamp 1751532392
transform 1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__682__D
timestamp 1751532392
transform 1 0 25760 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__683__B
timestamp 1751532392
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__684__B
timestamp 1751532392
transform 1 0 18816 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__689__A
timestamp 1751532392
transform 1 0 21504 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__692__A
timestamp 1751532392
transform 1 0 21392 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__693__B
timestamp 1751532392
transform 1 0 15008 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__699__B
timestamp 1751532392
transform 1 0 17472 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__701__A
timestamp 1751532392
transform 1 0 16128 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__706__C
timestamp 1751532392
transform 1 0 19376 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__711__B
timestamp 1751532392
transform 1 0 15120 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__715__D
timestamp 1751532392
transform -1 0 20384 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__716__B
timestamp 1751532392
transform 1 0 18368 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__718__B
timestamp 1751532392
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__719__B
timestamp 1751532392
transform 1 0 28672 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__720__A
timestamp 1751532392
transform 1 0 26096 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__727__D
timestamp 1751532392
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__729__B
timestamp 1751532392
transform 1 0 35392 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__731__A
timestamp 1751532392
transform -1 0 20608 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__731__C
timestamp 1751532392
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__732__C
timestamp 1751532392
transform 1 0 35728 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__736__CLK
timestamp 1751532392
transform 1 0 25312 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__737__CLK
timestamp 1751532392
transform 1 0 29232 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__738__CLK
timestamp 1751532392
transform -1 0 32928 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__739__CLK
timestamp 1751532392
transform -1 0 36512 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__741__CLK
timestamp 1751532392
transform 1 0 17472 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__742__CLK
timestamp 1751532392
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__743__CLK
timestamp 1751532392
transform 1 0 16240 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__744__CLK
timestamp 1751532392
transform 1 0 17360 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__745__CLK
timestamp 1751532392
transform 1 0 26208 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__746__CLK
timestamp 1751532392
transform 1 0 26544 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__747__CLK
timestamp 1751532392
transform 1 0 30128 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__748__CLK
timestamp 1751532392
transform -1 0 35392 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__749__CLK
timestamp 1751532392
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__750__CLK
timestamp 1751532392
transform 1 0 30464 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__751__CLK
timestamp 1751532392
transform 1 0 34048 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__752__CLK
timestamp 1751532392
transform 1 0 31808 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__753__CLK
timestamp 1751532392
transform 1 0 25312 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__754__CLK
timestamp 1751532392
transform 1 0 36400 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__755__CLK
timestamp 1751532392
transform 1 0 34160 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__756__CLK
timestamp 1751532392
transform 1 0 37856 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__757__CLK
timestamp 1751532392
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__758__CLK
timestamp 1751532392
transform 1 0 40208 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__759__CLK
timestamp 1751532392
transform 1 0 36848 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__760__CLK
timestamp 1751532392
transform 1 0 36624 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__761__CLK
timestamp 1751532392
transform 1 0 40768 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__762__CLK
timestamp 1751532392
transform 1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__763__CLK
timestamp 1751532392
transform 1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__764__CLK
timestamp 1751532392
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__765__CLK
timestamp 1751532392
transform 1 0 40880 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__766__CLK
timestamp 1751532392
transform 1 0 41216 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__767__CLK
timestamp 1751532392
transform 1 0 39424 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__768__CLK
timestamp 1751532392
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__769__CLK
timestamp 1751532392
transform 1 0 33376 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__770__CLK
timestamp 1751532392
transform 1 0 11200 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__771__CLK
timestamp 1751532392
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__772__CLK
timestamp 1751532392
transform 1 0 5152 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__773__CLK
timestamp 1751532392
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__774__CLK
timestamp 1751532392
transform 1 0 9632 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__775__CLK
timestamp 1751532392
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__776__CLK
timestamp 1751532392
transform -1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__777__CLK
timestamp 1751532392
transform -1 0 5600 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__778__CLK
timestamp 1751532392
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__779__CLK
timestamp 1751532392
transform 1 0 14000 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__780__CLK
timestamp 1751532392
transform 1 0 7728 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__781__CLK
timestamp 1751532392
transform 1 0 5488 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__782__CLK
timestamp 1751532392
transform 1 0 5712 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__783__CLK
timestamp 1751532392
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__784__CLK
timestamp 1751532392
transform -1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__785__CLK
timestamp 1751532392
transform -1 0 9968 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__786__CLK
timestamp 1751532392
transform 1 0 24864 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__787__CLK
timestamp 1751532392
transform -1 0 25200 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__788__CLK
timestamp 1751532392
transform 1 0 17696 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__789__CLK
timestamp 1751532392
transform 1 0 11200 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__791__CLK
timestamp 1751532392
transform 1 0 21616 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__794__CLK
timestamp 1751532392
transform 1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__795__CLK
timestamp 1751532392
transform 1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__796__CLK
timestamp 1751532392
transform 1 0 33040 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__797__CLK
timestamp 1751532392
transform 1 0 36064 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__799__A
timestamp 1751532392
transform 1 0 43232 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 21280 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_0__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 12880 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_1__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 17472 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_2__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_3__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 16352 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_4__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 27776 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_5__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 33040 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_6__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 28112 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_7__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload0_A
timestamp 1751532392
transform 1 0 9856 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload1_A
timestamp 1751532392
transform 1 0 13776 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload2_A
timestamp 1751532392
transform 1 0 8064 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload4_A
timestamp 1751532392
transform 1 0 29456 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload5_A
timestamp 1751532392
transform 1 0 27664 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input2_A
timestamp 1751532392
transform -1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0_wb_clk_i dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751661108
transform 1 0 21504 0 -1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_0__f_wb_clk_i
timestamp 1751661108
transform 1 0 9856 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_1__f_wb_clk_i
timestamp 1751661108
transform 1 0 14224 0 1 14112
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_2__f_wb_clk_i
timestamp 1751661108
transform -1 0 11872 0 1 29792
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_3__f_wb_clk_i
timestamp 1751661108
transform 1 0 13328 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_4__f_wb_clk_i
timestamp 1751661108
transform 1 0 29008 0 1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_5__f_wb_clk_i
timestamp 1751661108
transform 1 0 33264 0 1 17248
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_6__f_wb_clk_i
timestamp 1751661108
transform 1 0 29008 0 1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_7__f_wb_clk_i
timestamp 1751661108
transform 1 0 32928 0 -1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload0
timestamp 1751532043
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751633659
transform -1 0 14224 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload2
timestamp 1751633659
transform 1 0 8288 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload3
timestamp 1751661108
transform -1 0 15456 0 -1 31360
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload4
timestamp 1751532043
transform 1 0 29008 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  clkload5
timestamp 1751532043
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_18
timestamp 1751532351
transform 1 0 3360 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_36
timestamp 1751532351
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_52
timestamp 1751532351
transform 1 0 7168 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_70
timestamp 1751532351
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_86
timestamp 1751532351
transform 1 0 10976 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_104
timestamp 1751532351
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_120
timestamp 1751532351
transform 1 0 14784 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_138
timestamp 1751532351
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_154
timestamp 1751532351
transform 1 0 18592 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_172
timestamp 1751532351
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_188
timestamp 1751532351
transform 1 0 22400 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_206
timestamp 1751532351
transform 1 0 24416 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_222
timestamp 1751532351
transform 1 0 26208 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_240
timestamp 1751532351
transform 1 0 28224 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_256
timestamp 1751532351
transform 1 0 30016 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_274
timestamp 1751532351
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_290
timestamp 1751532351
transform 1 0 33824 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_308
timestamp 1751532351
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_324
timestamp 1751532351
transform 1 0 37632 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_342
timestamp 1751532351
transform 1 0 39648 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_358
timestamp 1751532351
transform 1 0 41440 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_376 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 43456 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_2
timestamp 1751532351
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_18
timestamp 1751532351
transform 1 0 3360 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_34
timestamp 1751532351
transform 1 0 5152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_50 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 6944 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_52 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 7168 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_59
timestamp 1751532312
transform 1 0 7952 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_67
timestamp 1751532440
transform 1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_69
timestamp 1751532423
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_72
timestamp 1751532351
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_88
timestamp 1751532351
transform 1 0 11200 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_104
timestamp 1751532351
transform 1 0 12992 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_120
timestamp 1751532351
transform 1 0 14784 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_136
timestamp 1751532440
transform 1 0 16576 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_142
timestamp 1751532351
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 19040 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_162
timestamp 1751532440
transform 1 0 19488 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_164
timestamp 1751532423
transform 1 0 19712 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_172
timestamp 1751532351
transform 1 0 20608 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_188
timestamp 1751532312
transform 1 0 22400 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_196
timestamp 1751532246
transform 1 0 23296 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_200
timestamp 1751532423
transform 1 0 23744 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_207
timestamp 1751532440
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_209
timestamp 1751532423
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_212
timestamp 1751532351
transform 1 0 25088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_255
timestamp 1751532440
transform 1 0 29904 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_259
timestamp 1751532351
transform 1 0 30352 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_275
timestamp 1751532246
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_279
timestamp 1751532423
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_282
timestamp 1751532351
transform 1 0 32928 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_298
timestamp 1751532351
transform 1 0 34720 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_314
timestamp 1751532351
transform 1 0 36512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_330
timestamp 1751532351
transform 1 0 38304 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_346
timestamp 1751532246
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_352
timestamp 1751532351
transform 1 0 40768 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_368
timestamp 1751532351
transform 1 0 42560 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_2
timestamp 1751532351
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_18
timestamp 1751532351
transform 1 0 3360 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_34
timestamp 1751532423
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_37
timestamp 1751532312
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_45
timestamp 1751532423
transform 1 0 6384 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_73
timestamp 1751532440
transform 1 0 9520 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_77
timestamp 1751532423
transform 1 0 9968 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_107
timestamp 1751532440
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_138
timestamp 1751532246
transform 1 0 16800 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_142
timestamp 1751532423
transform 1 0 17248 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_172
timestamp 1751532440
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_174
timestamp 1751532423
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_177
timestamp 1751532351
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_220
timestamp 1751532440
transform 1 0 25984 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_224
timestamp 1751532312
transform 1 0 26432 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_232
timestamp 1751532246
transform 1 0 27328 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_236
timestamp 1751532423
transform 1 0 27776 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_243
timestamp 1751532440
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_247
timestamp 1751532351
transform 1 0 29008 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_263
timestamp 1751532440
transform 1 0 30800 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_272
timestamp 1751532423
transform 1 0 31808 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_300
timestamp 1751532440
transform 1 0 34944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_304
timestamp 1751532312
transform 1 0 35392 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_312
timestamp 1751532440
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_314
timestamp 1751532423
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_317
timestamp 1751532351
transform 1 0 36848 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_333
timestamp 1751532351
transform 1 0 38640 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_349
timestamp 1751532351
transform 1 0 40432 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_365
timestamp 1751532351
transform 1 0 42224 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_381
timestamp 1751532440
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_383
timestamp 1751532423
transform 1 0 44240 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_2
timestamp 1751532351
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_18
timestamp 1751532351
transform 1 0 3360 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_34
timestamp 1751532351
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_50
timestamp 1751532246
transform 1 0 6944 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_54
timestamp 1751532440
transform 1 0 7392 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_76
timestamp 1751532351
transform 1 0 9856 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_92
timestamp 1751532440
transform 1 0 11648 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_105
timestamp 1751532246
transform 1 0 13104 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_115
timestamp 1751532351
transform 1 0 14224 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_131
timestamp 1751532312
transform 1 0 16016 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_139
timestamp 1751532423
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_142
timestamp 1751532351
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_158
timestamp 1751532246
transform 1 0 19040 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_183
timestamp 1751532246
transform 1 0 21840 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_194
timestamp 1751532246
transform 1 0 23072 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_205
timestamp 1751532246
transform 1 0 24304 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_209
timestamp 1751532423
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_212
timestamp 1751532351
transform 1 0 25088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_228
timestamp 1751532440
transform 1 0 26880 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_257
timestamp 1751532246
transform 1 0 30128 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_261
timestamp 1751532423
transform 1 0 30576 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_275
timestamp 1751532246
transform 1 0 32144 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_279
timestamp 1751532423
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_288
timestamp 1751532351
transform 1 0 33600 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_304
timestamp 1751532351
transform 1 0 35392 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_320
timestamp 1751532351
transform 1 0 37184 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_336
timestamp 1751532312
transform 1 0 38976 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_344
timestamp 1751532246
transform 1 0 39872 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_348
timestamp 1751532440
transform 1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_352
timestamp 1751532351
transform 1 0 40768 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_368
timestamp 1751532351
transform 1 0 42560 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_2
timestamp 1751532351
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_18
timestamp 1751532351
transform 1 0 3360 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_34
timestamp 1751532423
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_37
timestamp 1751532351
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_53
timestamp 1751532423
transform 1 0 7280 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_64
timestamp 1751532351
transform 1 0 8512 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_80
timestamp 1751532351
transform 1 0 10304 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_96
timestamp 1751532440
transform 1 0 12096 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_98
timestamp 1751532423
transform 1 0 12320 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_107
timestamp 1751532351
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_123
timestamp 1751532351
transform 1 0 15120 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_139
timestamp 1751532351
transform 1 0 16912 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_155
timestamp 1751532312
transform 1 0 18704 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_163
timestamp 1751532246
transform 1 0 19600 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_167
timestamp 1751532440
transform 1 0 20048 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_171
timestamp 1751532246
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_177
timestamp 1751532351
transform 1 0 21168 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_193
timestamp 1751532351
transform 1 0 22960 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_209
timestamp 1751532351
transform 1 0 24752 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_225
timestamp 1751532351
transform 1 0 26544 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_241
timestamp 1751532246
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_247
timestamp 1751532312
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_255
timestamp 1751532246
transform 1 0 29904 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_259
timestamp 1751532440
transform 1 0 30352 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_261
timestamp 1751532423
transform 1 0 30576 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_276
timestamp 1751532351
transform 1 0 32256 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_292
timestamp 1751532351
transform 1 0 34048 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_308
timestamp 1751532246
transform 1 0 35840 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_312
timestamp 1751532440
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_314
timestamp 1751532423
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_317
timestamp 1751532351
transform 1 0 36848 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_333
timestamp 1751532351
transform 1 0 38640 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_349
timestamp 1751532351
transform 1 0 40432 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_365
timestamp 1751532351
transform 1 0 42224 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_381
timestamp 1751532440
transform 1 0 44016 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_383
timestamp 1751532423
transform 1 0 44240 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_2
timestamp 1751532351
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_18
timestamp 1751532351
transform 1 0 3360 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_34
timestamp 1751532351
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_50
timestamp 1751532351
transform 1 0 6944 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_66
timestamp 1751532246
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_72
timestamp 1751532351
transform 1 0 9408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_88
timestamp 1751532351
transform 1 0 11200 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_104
timestamp 1751532312
transform 1 0 12992 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_112
timestamp 1751532440
transform 1 0 13888 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_121
timestamp 1751532351
transform 1 0 14896 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_137
timestamp 1751532440
transform 1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_139
timestamp 1751532423
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_142
timestamp 1751532246
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_146
timestamp 1751532423
transform 1 0 17696 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_153
timestamp 1751532312
transform 1 0 18480 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_161
timestamp 1751532246
transform 1 0 19376 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_165
timestamp 1751532440
transform 1 0 19824 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_174
timestamp 1751532246
transform 1 0 20832 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_178
timestamp 1751532440
transform 1 0 21280 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_180
timestamp 1751532423
transform 1 0 21504 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_188
timestamp 1751532351
transform 1 0 22400 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_204
timestamp 1751532246
transform 1 0 24192 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_208
timestamp 1751532440
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_212
timestamp 1751532351
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_228
timestamp 1751532351
transform 1 0 26880 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_244
timestamp 1751532351
transform 1 0 28672 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_260
timestamp 1751532351
transform 1 0 30464 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_276
timestamp 1751532246
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_282
timestamp 1751532351
transform 1 0 32928 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_298
timestamp 1751532351
transform 1 0 34720 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_314
timestamp 1751532351
transform 1 0 36512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_330
timestamp 1751532351
transform 1 0 38304 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_346
timestamp 1751532246
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_352
timestamp 1751532351
transform 1 0 40768 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_368
timestamp 1751532351
transform 1 0 42560 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_2
timestamp 1751532351
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_18
timestamp 1751532351
transform 1 0 3360 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_34
timestamp 1751532423
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_37
timestamp 1751532351
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_53
timestamp 1751532351
transform 1 0 7280 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_69
timestamp 1751532312
transform 1 0 9072 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_77
timestamp 1751532246
transform 1 0 9968 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_81
timestamp 1751532423
transform 1 0 10416 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_89
timestamp 1751532351
transform 1 0 11312 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_117
timestamp 1751532440
transform 1 0 14448 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_121
timestamp 1751532312
transform 1 0 14896 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_129
timestamp 1751532246
transform 1 0 15792 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_173
timestamp 1751532440
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_191
timestamp 1751532312
transform 1 0 22736 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_199
timestamp 1751532423
transform 1 0 23632 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_207
timestamp 1751532351
transform 1 0 24528 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_223
timestamp 1751532351
transform 1 0 26320 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_239
timestamp 1751532246
transform 1 0 28112 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_243
timestamp 1751532440
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_247
timestamp 1751532351
transform 1 0 29008 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_263
timestamp 1751532351
transform 1 0 30800 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_279
timestamp 1751532351
transform 1 0 32592 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_295
timestamp 1751532351
transform 1 0 34384 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_311
timestamp 1751532246
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_317
timestamp 1751532351
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_333
timestamp 1751532351
transform 1 0 38640 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_349
timestamp 1751532351
transform 1 0 40432 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_365
timestamp 1751532351
transform 1 0 42224 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_381
timestamp 1751532440
transform 1 0 44016 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_383
timestamp 1751532423
transform 1 0 44240 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_2
timestamp 1751532351
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_18
timestamp 1751532246
transform 1 0 3360 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_22
timestamp 1751532423
transform 1 0 3808 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_29
timestamp 1751532351
transform 1 0 4592 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_45
timestamp 1751532246
transform 1 0 6384 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_49
timestamp 1751532440
transform 1 0 6832 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_62
timestamp 1751532312
transform 1 0 8288 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_72
timestamp 1751532423
transform 1 0 9408 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_114
timestamp 1751532351
transform 1 0 14112 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_130
timestamp 1751532312
transform 1 0 15904 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_138
timestamp 1751532440
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_142
timestamp 1751532351
transform 1 0 17248 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_158
timestamp 1751532246
transform 1 0 19040 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_169
timestamp 1751532246
transform 1 0 20272 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_175
timestamp 1751532351
transform 1 0 20944 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_191
timestamp 1751532351
transform 1 0 22736 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_207
timestamp 1751532440
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_209
timestamp 1751532423
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_219
timestamp 1751532246
transform 1 0 25872 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_223
timestamp 1751532440
transform 1 0 26320 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_227
timestamp 1751532246
transform 1 0 26768 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_231
timestamp 1751532423
transform 1 0 27216 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_234
timestamp 1751532351
transform 1 0 27552 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_250
timestamp 1751532351
transform 1 0 29344 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_266
timestamp 1751532246
transform 1 0 31136 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_270
timestamp 1751532440
transform 1 0 31584 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_272
timestamp 1751532423
transform 1 0 31808 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_295
timestamp 1751532351
transform 1 0 34384 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_311
timestamp 1751532351
transform 1 0 36176 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_327
timestamp 1751532351
transform 1 0 37968 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_343
timestamp 1751532246
transform 1 0 39760 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_347
timestamp 1751532440
transform 1 0 40208 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_349
timestamp 1751532423
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_352
timestamp 1751532351
transform 1 0 40768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_368
timestamp 1751532351
transform 1 0 42560 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_2
timestamp 1751532246
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_6
timestamp 1751532440
transform 1 0 2016 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_37
timestamp 1751532440
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_41
timestamp 1751532312
transform 1 0 5936 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_49
timestamp 1751532440
transform 1 0 6832 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_71
timestamp 1751532351
transform 1 0 9296 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_87
timestamp 1751532440
transform 1 0 11088 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_89
timestamp 1751532423
transform 1 0 11312 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_92
timestamp 1751532312
transform 1 0 11648 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_100
timestamp 1751532246
transform 1 0 12544 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_104
timestamp 1751532423
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_107
timestamp 1751532351
transform 1 0 13328 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_123
timestamp 1751532351
transform 1 0 15120 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_139
timestamp 1751532351
transform 1 0 16912 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_155
timestamp 1751532351
transform 1 0 18704 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_171
timestamp 1751532246
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_177
timestamp 1751532351
transform 1 0 21168 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_193
timestamp 1751532246
transform 1 0 22960 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_197
timestamp 1751532423
transform 1 0 23408 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_232
timestamp 1751532440
transform 1 0 27328 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_241
timestamp 1751532246
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_247
timestamp 1751532312
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_255
timestamp 1751532246
transform 1 0 29904 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_259
timestamp 1751532423
transform 1 0 30352 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_262
timestamp 1751532423
transform 1 0 30688 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_281
timestamp 1751532246
transform 1 0 32816 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_312
timestamp 1751532440
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_314
timestamp 1751532423
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_317
timestamp 1751532440
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_321
timestamp 1751532351
transform 1 0 37296 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_337
timestamp 1751532351
transform 1 0 39088 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_353
timestamp 1751532351
transform 1 0 40880 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_369
timestamp 1751532312
transform 1 0 42672 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_377
timestamp 1751532246
transform 1 0 43568 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_381
timestamp 1751532440
transform 1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_383
timestamp 1751532423
transform 1 0 44240 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_2
timestamp 1751532351
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_18
timestamp 1751532351
transform 1 0 3360 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_34
timestamp 1751532351
transform 1 0 5152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_50
timestamp 1751532351
transform 1 0 6944 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_66
timestamp 1751532246
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_78
timestamp 1751532440
transform 1 0 10080 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_82
timestamp 1751532312
transform 1 0 10528 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_90
timestamp 1751532246
transform 1 0 11424 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_94
timestamp 1751532440
transform 1 0 11872 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_106
timestamp 1751532351
transform 1 0 13216 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_122
timestamp 1751532351
transform 1 0 15008 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_138
timestamp 1751532440
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_142
timestamp 1751532351
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_158
timestamp 1751532351
transform 1 0 19040 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_174
timestamp 1751532312
transform 1 0 20832 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_182
timestamp 1751532440
transform 1 0 21728 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_191
timestamp 1751532312
transform 1 0 22736 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_199
timestamp 1751532246
transform 1 0 23632 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_203
timestamp 1751532440
transform 1 0 24080 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_205
timestamp 1751532423
transform 1 0 24304 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_222
timestamp 1751532440
transform 1 0 26208 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_226
timestamp 1751532246
transform 1 0 26656 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_230
timestamp 1751532440
transform 1 0 27104 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_232
timestamp 1751532423
transform 1 0 27328 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_274
timestamp 1751532246
transform 1 0 32032 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_278
timestamp 1751532440
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_289
timestamp 1751532351
transform 1 0 33712 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_305
timestamp 1751532312
transform 1 0 35504 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_313
timestamp 1751532440
transform 1 0 36400 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_344
timestamp 1751532246
transform 1 0 39872 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_348
timestamp 1751532440
transform 1 0 40320 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_352
timestamp 1751532351
transform 1 0 40768 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_368
timestamp 1751532351
transform 1 0 42560 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_2
timestamp 1751532351
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_18
timestamp 1751532423
transform 1 0 3360 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_25
timestamp 1751532312
transform 1 0 4144 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_33
timestamp 1751532440
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_37
timestamp 1751532312
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_45
timestamp 1751532440
transform 1 0 6384 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_58
timestamp 1751532351
transform 1 0 7840 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_74
timestamp 1751532351
transform 1 0 9632 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_90
timestamp 1751532312
transform 1 0 11424 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_98
timestamp 1751532246
transform 1 0 12320 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_102
timestamp 1751532440
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_104
timestamp 1751532423
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_107
timestamp 1751532351
transform 1 0 13328 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_123
timestamp 1751532351
transform 1 0 15120 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_139
timestamp 1751532351
transform 1 0 16912 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_155
timestamp 1751532312
transform 1 0 18704 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_170
timestamp 1751532246
transform 1 0 20384 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_174
timestamp 1751532423
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_177
timestamp 1751532351
transform 1 0 21168 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_193
timestamp 1751532351
transform 1 0 22960 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_209
timestamp 1751532351
transform 1 0 24752 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_225
timestamp 1751532312
transform 1 0 26544 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_233
timestamp 1751532246
transform 1 0 27440 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_243
timestamp 1751532440
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_247
timestamp 1751532351
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_263
timestamp 1751532351
transform 1 0 30800 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_279
timestamp 1751532351
transform 1 0 32592 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_295
timestamp 1751532351
transform 1 0 34384 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_311
timestamp 1751532246
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_317
timestamp 1751532312
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_325
timestamp 1751532246
transform 1 0 37744 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_329
timestamp 1751532423
transform 1 0 38192 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_336
timestamp 1751532351
transform 1 0 38976 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_381
timestamp 1751532440
transform 1 0 44016 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_383
timestamp 1751532423
transform 1 0 44240 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_2
timestamp 1751532246
transform 1 0 1568 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_6
timestamp 1751532440
transform 1 0 2016 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_35
timestamp 1751532440
transform 1 0 5264 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_39
timestamp 1751532351
transform 1 0 5712 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_55
timestamp 1751532312
transform 1 0 7504 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_63
timestamp 1751532246
transform 1 0 8400 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_67
timestamp 1751532440
transform 1 0 8848 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_69
timestamp 1751532423
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_72
timestamp 1751532351
transform 1 0 9408 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_88
timestamp 1751532312
transform 1 0 11200 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_96
timestamp 1751532440
transform 1 0 12096 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_98
timestamp 1751532423
transform 1 0 12320 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_113
timestamp 1751532351
transform 1 0 14000 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_129
timestamp 1751532312
transform 1 0 15792 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_137
timestamp 1751532423
transform 1 0 16688 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_142
timestamp 1751532423
transform 1 0 17248 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_177
timestamp 1751532440
transform 1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_181
timestamp 1751532351
transform 1 0 21616 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_197
timestamp 1751532312
transform 1 0 23408 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_205
timestamp 1751532246
transform 1 0 24304 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_209
timestamp 1751532423
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_212
timestamp 1751532351
transform 1 0 25088 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_228
timestamp 1751532351
transform 1 0 26880 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_244
timestamp 1751532351
transform 1 0 28672 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_260
timestamp 1751532351
transform 1 0 30464 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_276
timestamp 1751532246
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_282
timestamp 1751532351
transform 1 0 32928 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_298
timestamp 1751532351
transform 1 0 34720 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_314
timestamp 1751532351
transform 1 0 36512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_330
timestamp 1751532440
transform 1 0 38304 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_342
timestamp 1751532312
transform 1 0 39648 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_352
timestamp 1751532440
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_354
timestamp 1751532423
transform 1 0 40992 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_361
timestamp 1751532351
transform 1 0 41776 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_377
timestamp 1751532246
transform 1 0 43568 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_381
timestamp 1751532440
transform 1 0 44016 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_383
timestamp 1751532423
transform 1 0 44240 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_2
timestamp 1751532351
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_18
timestamp 1751532351
transform 1 0 3360 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_34
timestamp 1751532423
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_37
timestamp 1751532312
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_45
timestamp 1751532246
transform 1 0 6384 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_49
timestamp 1751532423
transform 1 0 6832 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_74
timestamp 1751532312
transform 1 0 9632 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_82
timestamp 1751532246
transform 1 0 10528 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_86
timestamp 1751532423
transform 1 0 10976 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_111
timestamp 1751532440
transform 1 0 13776 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_115
timestamp 1751532351
transform 1 0 14224 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_131
timestamp 1751532312
transform 1 0 16016 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_139
timestamp 1751532246
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_143
timestamp 1751532423
transform 1 0 17360 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_173
timestamp 1751532440
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_188
timestamp 1751532351
transform 1 0 22400 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_204
timestamp 1751532351
transform 1 0 24192 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_220
timestamp 1751532351
transform 1 0 25984 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_236
timestamp 1751532312
transform 1 0 27776 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_244
timestamp 1751532423
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_247
timestamp 1751532351
transform 1 0 29008 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_263
timestamp 1751532351
transform 1 0 30800 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_279
timestamp 1751532312
transform 1 0 32592 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_287
timestamp 1751532246
transform 1 0 33488 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_291
timestamp 1751532440
transform 1 0 33936 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_293
timestamp 1751532423
transform 1 0 34160 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_300
timestamp 1751532312
transform 1 0 34944 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_308
timestamp 1751532246
transform 1 0 35840 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_312
timestamp 1751532440
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_314
timestamp 1751532423
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_317
timestamp 1751532312
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_325
timestamp 1751532440
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_327
timestamp 1751532423
transform 1 0 37968 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_335
timestamp 1751532312
transform 1 0 38864 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_12_353
timestamp 1751532351
transform 1 0 40880 0 1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_369
timestamp 1751532312
transform 1 0 42672 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_377
timestamp 1751532246
transform 1 0 43568 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_381
timestamp 1751532440
transform 1 0 44016 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_383
timestamp 1751532423
transform 1 0 44240 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_2
timestamp 1751532351
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_18
timestamp 1751532351
transform 1 0 3360 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_34
timestamp 1751532351
transform 1 0 5152 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_50
timestamp 1751532351
transform 1 0 6944 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_66
timestamp 1751532246
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_72
timestamp 1751532312
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_80
timestamp 1751532423
transform 1 0 10304 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_125
timestamp 1751532440
transform 1 0 15344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_129
timestamp 1751532312
transform 1 0 15792 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_137
timestamp 1751532440
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_139
timestamp 1751532423
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_142
timestamp 1751532351
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_158
timestamp 1751532246
transform 1 0 19040 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_183
timestamp 1751532351
transform 1 0 21840 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_199
timestamp 1751532312
transform 1 0 23632 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_207
timestamp 1751532440
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_209
timestamp 1751532423
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_212
timestamp 1751532351
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_228
timestamp 1751532351
transform 1 0 26880 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_244
timestamp 1751532351
transform 1 0 28672 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_260
timestamp 1751532351
transform 1 0 30464 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_276
timestamp 1751532246
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_282
timestamp 1751532246
transform 1 0 32928 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_286
timestamp 1751532440
transform 1 0 33376 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_315
timestamp 1751532440
transform 1 0 36624 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_319
timestamp 1751532351
transform 1 0 37072 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_335
timestamp 1751532312
transform 1 0 38864 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_343
timestamp 1751532246
transform 1 0 39760 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_347
timestamp 1751532440
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_349
timestamp 1751532423
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_352
timestamp 1751532351
transform 1 0 40768 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_368
timestamp 1751532351
transform 1 0 42560 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_2
timestamp 1751532351
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_18
timestamp 1751532351
transform 1 0 3360 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_34
timestamp 1751532423
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_37
timestamp 1751532440
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_60
timestamp 1751532351
transform 1 0 8064 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_78
timestamp 1751532351
transform 1 0 10080 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_101
timestamp 1751532246
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_107
timestamp 1751532423
transform 1 0 13328 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_140
timestamp 1751532440
transform 1 0 17024 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_144
timestamp 1751532351
transform 1 0 17472 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_160
timestamp 1751532312
transform 1 0 19264 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_168
timestamp 1751532423
transform 1 0 20160 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_171
timestamp 1751532246
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_177
timestamp 1751532351
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_193
timestamp 1751532312
transform 1 0 22960 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_201
timestamp 1751532246
transform 1 0 23856 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_205
timestamp 1751532440
transform 1 0 24304 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_207
timestamp 1751532423
transform 1 0 24528 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_214
timestamp 1751532440
transform 1 0 25312 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_218
timestamp 1751532312
transform 1 0 25760 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_226
timestamp 1751532440
transform 1 0 26656 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_235
timestamp 1751532246
transform 1 0 27664 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_241
timestamp 1751532246
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_247
timestamp 1751532246
transform 1 0 29008 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_253
timestamp 1751532423
transform 1 0 29680 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_281
timestamp 1751532440
transform 1 0 32816 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_285
timestamp 1751532246
transform 1 0 33264 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_302
timestamp 1751532312
transform 1 0 35168 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_310
timestamp 1751532246
transform 1 0 36064 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_314
timestamp 1751532423
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_317
timestamp 1751532312
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_325
timestamp 1751532246
transform 1 0 37744 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_329
timestamp 1751532440
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_341
timestamp 1751532246
transform 1 0 39536 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_345
timestamp 1751532440
transform 1 0 39984 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_382
timestamp 1751532440
transform 1 0 44128 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_2
timestamp 1751532351
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_18
timestamp 1751532312
transform 1 0 3360 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_26
timestamp 1751532440
transform 1 0 4256 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_55
timestamp 1751532440
transform 1 0 7504 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_59
timestamp 1751532312
transform 1 0 7952 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_67
timestamp 1751532440
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_69
timestamp 1751532423
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_101
timestamp 1751532440
transform 1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_105
timestamp 1751532246
transform 1 0 13104 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_109
timestamp 1751532440
transform 1 0 13552 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_142
timestamp 1751532440
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_146
timestamp 1751532351
transform 1 0 17696 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_162
timestamp 1751532351
transform 1 0 19488 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_178
timestamp 1751532351
transform 1 0 21280 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_194
timestamp 1751532246
transform 1 0 23072 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_246
timestamp 1751532423
transform 1 0 28896 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_251
timestamp 1751532423
transform 1 0 29456 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_276
timestamp 1751532440
transform 1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_282
timestamp 1751532312
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_290
timestamp 1751532440
transform 1 0 33824 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_292
timestamp 1751532423
transform 1 0 34048 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_302
timestamp 1751532351
transform 1 0 35168 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_318
timestamp 1751532312
transform 1 0 36960 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_336
timestamp 1751532246
transform 1 0 38976 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_352
timestamp 1751532351
transform 1 0 40768 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_368
timestamp 1751532351
transform 1 0 42560 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_2
timestamp 1751532351
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_18
timestamp 1751532351
transform 1 0 3360 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_34
timestamp 1751532423
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_37
timestamp 1751532351
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_53
timestamp 1751532351
transform 1 0 7280 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_69
timestamp 1751532351
transform 1 0 9072 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_85
timestamp 1751532351
transform 1 0 10864 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_101
timestamp 1751532246
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_107
timestamp 1751532312
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_115
timestamp 1751532246
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_119
timestamp 1751532440
transform 1 0 14672 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_127
timestamp 1751532351
transform 1 0 15568 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_143
timestamp 1751532351
transform 1 0 17360 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_159
timestamp 1751532351
transform 1 0 19152 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_177
timestamp 1751532440
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_181
timestamp 1751532312
transform 1 0 21616 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_189
timestamp 1751532246
transform 1 0 22512 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_201
timestamp 1751532312
transform 1 0 23856 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_209
timestamp 1751532423
transform 1 0 24752 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_212
timestamp 1751532351
transform 1 0 25088 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_228
timestamp 1751532312
transform 1 0 26880 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_272
timestamp 1751532351
transform 1 0 31808 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_288
timestamp 1751532351
transform 1 0 33600 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_304
timestamp 1751532312
transform 1 0 35392 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_312
timestamp 1751532440
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_314
timestamp 1751532423
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_317
timestamp 1751532351
transform 1 0 36848 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_333
timestamp 1751532440
transform 1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_335
timestamp 1751532423
transform 1 0 38864 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_342
timestamp 1751532351
transform 1 0 39648 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_358
timestamp 1751532351
transform 1 0 41440 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_374
timestamp 1751532312
transform 1 0 43232 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_382
timestamp 1751532440
transform 1 0 44128 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_2
timestamp 1751532351
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_18
timestamp 1751532351
transform 1 0 3360 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_34
timestamp 1751532351
transform 1 0 5152 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_50
timestamp 1751532351
transform 1 0 6944 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_66
timestamp 1751532246
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_72
timestamp 1751532351
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_88
timestamp 1751532351
transform 1 0 11200 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_104
timestamp 1751532312
transform 1 0 12992 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_112
timestamp 1751532246
transform 1 0 13888 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_116
timestamp 1751532423
transform 1 0 14336 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_124
timestamp 1751532351
transform 1 0 15232 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_142
timestamp 1751532351
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_158
timestamp 1751532312
transform 1 0 19040 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_166
timestamp 1751532440
transform 1 0 19936 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_168
timestamp 1751532423
transform 1 0 20160 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_179
timestamp 1751532440
transform 1 0 21392 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_189
timestamp 1751532351
transform 1 0 22512 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_205
timestamp 1751532246
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_209
timestamp 1751532423
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_212
timestamp 1751532351
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_228
timestamp 1751532312
transform 1 0 26880 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_236
timestamp 1751532440
transform 1 0 27776 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_251
timestamp 1751532351
transform 1 0 29456 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_267
timestamp 1751532312
transform 1 0 31248 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_275
timestamp 1751532246
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_279
timestamp 1751532423
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_282
timestamp 1751532246
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_286
timestamp 1751532440
transform 1 0 33376 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_296
timestamp 1751532351
transform 1 0 34496 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_312
timestamp 1751532312
transform 1 0 36288 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_320
timestamp 1751532440
transform 1 0 37184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_324
timestamp 1751532312
transform 1 0 37632 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_332
timestamp 1751532440
transform 1 0 38528 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_334
timestamp 1751532423
transform 1 0 38752 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_345
timestamp 1751532246
transform 1 0 39984 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_349
timestamp 1751532423
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_352
timestamp 1751532351
transform 1 0 40768 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_368
timestamp 1751532351
transform 1 0 42560 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_2
timestamp 1751532351
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_18
timestamp 1751532351
transform 1 0 3360 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_34
timestamp 1751532423
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_37
timestamp 1751532351
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_53
timestamp 1751532246
transform 1 0 7280 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_57
timestamp 1751532440
transform 1 0 7728 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_86
timestamp 1751532440
transform 1 0 10976 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_90
timestamp 1751532312
transform 1 0 11424 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_98
timestamp 1751532246
transform 1 0 12320 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_102
timestamp 1751532440
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_104
timestamp 1751532423
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_107
timestamp 1751532246
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_111
timestamp 1751532440
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_113
timestamp 1751532423
transform 1 0 14000 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_130
timestamp 1751532312
transform 1 0 15904 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_138
timestamp 1751532246
transform 1 0 16800 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_142
timestamp 1751532423
transform 1 0 17248 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_149
timestamp 1751532351
transform 1 0 18032 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_165
timestamp 1751532312
transform 1 0 19824 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_173
timestamp 1751532440
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_184
timestamp 1751532440
transform 1 0 21952 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_188
timestamp 1751532351
transform 1 0 22400 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_204
timestamp 1751532351
transform 1 0 24192 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_220
timestamp 1751532312
transform 1 0 25984 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_228
timestamp 1751532246
transform 1 0 26880 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_234
timestamp 1751532312
transform 1 0 27552 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_242
timestamp 1751532440
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_244
timestamp 1751532423
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_247
timestamp 1751532351
transform 1 0 29008 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_263
timestamp 1751532351
transform 1 0 30800 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_279
timestamp 1751532246
transform 1 0 32592 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_310
timestamp 1751532246
transform 1 0 36064 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_314
timestamp 1751532423
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_317
timestamp 1751532423
transform 1 0 36848 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_330
timestamp 1751532351
transform 1 0 38304 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_346
timestamp 1751532246
transform 1 0 40096 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_350
timestamp 1751532423
transform 1 0 40544 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_380
timestamp 1751532246
transform 1 0 43904 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_2
timestamp 1751532351
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_18
timestamp 1751532351
transform 1 0 3360 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_34
timestamp 1751532351
transform 1 0 5152 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_50
timestamp 1751532351
transform 1 0 6944 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_66
timestamp 1751532246
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_78
timestamp 1751532440
transform 1 0 10080 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_82
timestamp 1751532351
transform 1 0 10528 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_98
timestamp 1751532312
transform 1 0 12320 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_106
timestamp 1751532246
transform 1 0 13216 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_110
timestamp 1751532440
transform 1 0 13664 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_112
timestamp 1751532423
transform 1 0 13888 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_139
timestamp 1751532423
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_148
timestamp 1751532351
transform 1 0 17920 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_164
timestamp 1751532423
transform 1 0 19712 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_178
timestamp 1751532440
transform 1 0 21280 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_182
timestamp 1751532351
transform 1 0 21728 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_198
timestamp 1751532312
transform 1 0 23520 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_206
timestamp 1751532246
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_212
timestamp 1751532312
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_220
timestamp 1751532423
transform 1 0 25984 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_241
timestamp 1751532440
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_243
timestamp 1751532423
transform 1 0 28560 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_253
timestamp 1751532440
transform 1 0 29680 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_255
timestamp 1751532423
transform 1 0 29904 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_270
timestamp 1751532312
transform 1 0 31584 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_278
timestamp 1751532440
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_282
timestamp 1751532440
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_311
timestamp 1751532440
transform 1 0 36176 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_315
timestamp 1751532351
transform 1 0 36624 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_343
timestamp 1751532246
transform 1 0 39760 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_347
timestamp 1751532440
transform 1 0 40208 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_349
timestamp 1751532423
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_352
timestamp 1751532440
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_358
timestamp 1751532351
transform 1 0 41440 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_374
timestamp 1751532312
transform 1 0 43232 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_382
timestamp 1751532440
transform 1 0 44128 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_2
timestamp 1751532440
transform 1 0 1568 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_31
timestamp 1751532440
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_37
timestamp 1751532440
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_53
timestamp 1751532351
transform 1 0 7280 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_80
timestamp 1751532440
transform 1 0 10304 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_82
timestamp 1751532423
transform 1 0 10528 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_89
timestamp 1751532351
transform 1 0 11312 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_107
timestamp 1751532351
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_123
timestamp 1751532351
transform 1 0 15120 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_139
timestamp 1751532246
transform 1 0 16912 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_143
timestamp 1751532440
transform 1 0 17360 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_145
timestamp 1751532423
transform 1 0 17584 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_177
timestamp 1751532351
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_193
timestamp 1751532351
transform 1 0 22960 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_209
timestamp 1751532312
transform 1 0 24752 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_223
timestamp 1751532351
transform 1 0 26320 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_239
timestamp 1751532246
transform 1 0 28112 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_243
timestamp 1751532440
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_247
timestamp 1751532351
transform 1 0 29008 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_263
timestamp 1751532351
transform 1 0 30800 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_279
timestamp 1751532351
transform 1 0 32592 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_295
timestamp 1751532246
transform 1 0 34384 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_309
timestamp 1751532246
transform 1 0 35952 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_313
timestamp 1751532440
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_317
timestamp 1751532351
transform 1 0 36848 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_333
timestamp 1751532246
transform 1 0 38640 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_337
timestamp 1751532423
transform 1 0 39088 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_344
timestamp 1751532246
transform 1 0 39872 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_348
timestamp 1751532440
transform 1 0 40320 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_350
timestamp 1751532423
transform 1 0 40544 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_20_361
timestamp 1751532351
transform 1 0 41776 0 1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_377
timestamp 1751532246
transform 1 0 43568 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_381
timestamp 1751532440
transform 1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_383
timestamp 1751532423
transform 1 0 44240 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_2
timestamp 1751532312
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_10
timestamp 1751532246
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_20
timestamp 1751532246
transform 1 0 3584 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_35
timestamp 1751532440
transform 1 0 5264 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_46
timestamp 1751532351
transform 1 0 6496 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_62
timestamp 1751532312
transform 1 0 8288 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_72
timestamp 1751532312
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_80
timestamp 1751532246
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_98
timestamp 1751532440
transform 1 0 12320 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_102
timestamp 1751532351
transform 1 0 12768 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_118
timestamp 1751532351
transform 1 0 14560 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_134
timestamp 1751532246
transform 1 0 16352 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_138
timestamp 1751532440
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_142
timestamp 1751532351
transform 1 0 17248 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_158
timestamp 1751532351
transform 1 0 19040 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_174
timestamp 1751532351
transform 1 0 20832 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_190
timestamp 1751532351
transform 1 0 22624 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_206
timestamp 1751532246
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_245
timestamp 1751532440
transform 1 0 28784 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_249
timestamp 1751532351
transform 1 0 29232 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_265
timestamp 1751532312
transform 1 0 31024 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_273
timestamp 1751532423
transform 1 0 31920 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_278
timestamp 1751532440
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_286
timestamp 1751532351
transform 1 0 33376 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_302
timestamp 1751532423
transform 1 0 35168 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_315
timestamp 1751532351
transform 1 0 36624 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_331
timestamp 1751532351
transform 1 0 38416 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_347
timestamp 1751532440
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_349
timestamp 1751532423
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_352
timestamp 1751532351
transform 1 0 40768 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_368
timestamp 1751532351
transform 1 0 42560 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_2
timestamp 1751532351
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_18
timestamp 1751532351
transform 1 0 3360 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_34
timestamp 1751532423
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_44
timestamp 1751532351
transform 1 0 6272 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_60
timestamp 1751532351
transform 1 0 8064 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_76
timestamp 1751532312
transform 1 0 9856 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_84
timestamp 1751532246
transform 1 0 10752 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_88
timestamp 1751532440
transform 1 0 11200 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_97
timestamp 1751532312
transform 1 0 12208 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_114
timestamp 1751532351
transform 1 0 14112 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_130
timestamp 1751532351
transform 1 0 15904 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_146
timestamp 1751532351
transform 1 0 17696 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_162
timestamp 1751532312
transform 1 0 19488 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_170
timestamp 1751532246
transform 1 0 20384 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_174
timestamp 1751532423
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_177
timestamp 1751532246
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_208
timestamp 1751532440
transform 1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_212
timestamp 1751532351
transform 1 0 25088 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_228
timestamp 1751532351
transform 1 0 26880 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_244
timestamp 1751532423
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_254
timestamp 1751532351
transform 1 0 29792 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_270
timestamp 1751532351
transform 1 0 31584 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_286
timestamp 1751532351
transform 1 0 33376 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_302
timestamp 1751532312
transform 1 0 35168 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_310
timestamp 1751532246
transform 1 0 36064 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_314
timestamp 1751532423
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_317
timestamp 1751532351
transform 1 0 36848 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_333
timestamp 1751532351
transform 1 0 38640 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_349
timestamp 1751532440
transform 1 0 40432 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_361
timestamp 1751532351
transform 1 0 41776 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_377
timestamp 1751532246
transform 1 0 43568 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_381
timestamp 1751532440
transform 1 0 44016 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_383
timestamp 1751532423
transform 1 0 44240 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_2
timestamp 1751532351
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_18
timestamp 1751532351
transform 1 0 3360 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_34
timestamp 1751532351
transform 1 0 5152 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_50
timestamp 1751532351
transform 1 0 6944 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_66
timestamp 1751532246
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_72
timestamp 1751532423
transform 1 0 9408 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_97
timestamp 1751532440
transform 1 0 12208 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_101
timestamp 1751532351
transform 1 0 12656 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_117
timestamp 1751532312
transform 1 0 14448 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_125
timestamp 1751532423
transform 1 0 15344 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_142
timestamp 1751532351
transform 1 0 17248 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_158
timestamp 1751532440
transform 1 0 19040 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_160
timestamp 1751532423
transform 1 0 19264 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_170
timestamp 1751532351
transform 1 0 20384 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_186
timestamp 1751532312
transform 1 0 22176 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_194
timestamp 1751532423
transform 1 0 23072 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_201
timestamp 1751532312
transform 1 0 23856 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_209
timestamp 1751532423
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_212
timestamp 1751532351
transform 1 0 25088 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_228
timestamp 1751532312
transform 1 0 26880 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_236
timestamp 1751532246
transform 1 0 27776 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_240
timestamp 1751532440
transform 1 0 28224 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_254
timestamp 1751532351
transform 1 0 29792 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_270
timestamp 1751532312
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_278
timestamp 1751532440
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_282
timestamp 1751532312
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_290
timestamp 1751532423
transform 1 0 33824 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_324
timestamp 1751532440
transform 1 0 37632 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_328
timestamp 1751532312
transform 1 0 38080 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_336
timestamp 1751532246
transform 1 0 38976 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_362
timestamp 1751532246
transform 1 0 41888 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_366
timestamp 1751532423
transform 1 0 42336 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_371
timestamp 1751532312
transform 1 0 42896 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_379
timestamp 1751532246
transform 1 0 43792 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_383
timestamp 1751532423
transform 1 0 44240 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_2
timestamp 1751532351
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_18
timestamp 1751532312
transform 1 0 3360 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_26
timestamp 1751532440
transform 1 0 4256 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_44
timestamp 1751532312
transform 1 0 6272 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_52
timestamp 1751532246
transform 1 0 7168 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_56
timestamp 1751532440
transform 1 0 7616 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_58
timestamp 1751532423
transform 1 0 7840 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_86
timestamp 1751532440
transform 1 0 10976 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_90
timestamp 1751532312
transform 1 0 11424 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_98
timestamp 1751532246
transform 1 0 12320 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_102
timestamp 1751532440
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_104
timestamp 1751532423
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_107
timestamp 1751532423
transform 1 0 13328 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_115
timestamp 1751532246
transform 1 0 14224 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_119
timestamp 1751532423
transform 1 0 14672 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_137
timestamp 1751532440
transform 1 0 16688 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_141
timestamp 1751532440
transform 1 0 17136 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_143
timestamp 1751532423
transform 1 0 17360 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_167
timestamp 1751532312
transform 1 0 20048 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_177
timestamp 1751532351
transform 1 0 21168 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_193
timestamp 1751532246
transform 1 0 22960 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_197
timestamp 1751532440
transform 1 0 23408 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_199
timestamp 1751532423
transform 1 0 23632 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_207
timestamp 1751532351
transform 1 0 24528 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_223
timestamp 1751532312
transform 1 0 26320 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_247
timestamp 1751532440
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_263
timestamp 1751532312
transform 1 0 30800 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_303
timestamp 1751532423
transform 1 0 35280 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_314
timestamp 1751532423
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_317
timestamp 1751532351
transform 1 0 36848 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_333
timestamp 1751532440
transform 1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_345
timestamp 1751532246
transform 1 0 39984 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_349
timestamp 1751532440
transform 1 0 40432 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_380
timestamp 1751532246
transform 1 0 43904 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_2
timestamp 1751532351
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_18
timestamp 1751532440
transform 1 0 3360 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_31
timestamp 1751532440
transform 1 0 4816 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_33
timestamp 1751532423
transform 1 0 5040 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_48
timestamp 1751532351
transform 1 0 6720 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_64
timestamp 1751532246
transform 1 0 8512 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_68
timestamp 1751532440
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_72
timestamp 1751532351
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_88
timestamp 1751532351
transform 1 0 11200 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_104
timestamp 1751532312
transform 1 0 12992 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_112
timestamp 1751532246
transform 1 0 13888 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_116
timestamp 1751532423
transform 1 0 14336 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_127
timestamp 1751532440
transform 1 0 15568 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_131
timestamp 1751532440
transform 1 0 16016 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_139
timestamp 1751532423
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_142
timestamp 1751532246
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_146
timestamp 1751532440
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_148
timestamp 1751532423
transform 1 0 17920 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_156
timestamp 1751532351
transform 1 0 18816 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_172
timestamp 1751532246
transform 1 0 20608 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_176
timestamp 1751532440
transform 1 0 21056 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_205
timestamp 1751532246
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_209
timestamp 1751532423
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_212
timestamp 1751532351
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_228
timestamp 1751532351
transform 1 0 26880 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_244
timestamp 1751532246
transform 1 0 28672 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_262
timestamp 1751532351
transform 1 0 30688 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_278
timestamp 1751532440
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_282
timestamp 1751532351
transform 1 0 32928 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_298
timestamp 1751532351
transform 1 0 34720 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_314
timestamp 1751532423
transform 1 0 36512 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_317
timestamp 1751532351
transform 1 0 36848 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_333
timestamp 1751532351
transform 1 0 38640 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_349
timestamp 1751532423
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_352
timestamp 1751532351
transform 1 0 40768 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_25_368
timestamp 1751532351
transform 1 0 42560 0 -1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_2
timestamp 1751532312
transform 1 0 1568 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_10
timestamp 1751532246
transform 1 0 2464 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_20
timestamp 1751532312
transform 1 0 3584 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_28
timestamp 1751532440
transform 1 0 4480 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_30
timestamp 1751532423
transform 1 0 4704 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_33
timestamp 1751532440
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_37
timestamp 1751532351
transform 1 0 5488 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_53
timestamp 1751532351
transform 1 0 7280 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_69
timestamp 1751532246
transform 1 0 9072 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_79
timestamp 1751532312
transform 1 0 10192 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_87
timestamp 1751532246
transform 1 0 11088 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_97
timestamp 1751532312
transform 1 0 12208 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_107
timestamp 1751532312
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_115
timestamp 1751532246
transform 1 0 14224 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_119
timestamp 1751532440
transform 1 0 14672 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_121
timestamp 1751532423
transform 1 0 14896 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_130
timestamp 1751532351
transform 1 0 15904 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_146
timestamp 1751532351
transform 1 0 17696 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_162
timestamp 1751532312
transform 1 0 19488 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_170
timestamp 1751532246
transform 1 0 20384 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_174
timestamp 1751532423
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_177
timestamp 1751532312
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_185
timestamp 1751532246
transform 1 0 22064 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_189
timestamp 1751532440
transform 1 0 22512 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_191
timestamp 1751532423
transform 1 0 22736 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_211
timestamp 1751532440
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_215
timestamp 1751532351
transform 1 0 25424 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_231
timestamp 1751532312
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_239
timestamp 1751532246
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_243
timestamp 1751532440
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_247
timestamp 1751532351
transform 1 0 29008 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_263
timestamp 1751532351
transform 1 0 30800 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_279
timestamp 1751532351
transform 1 0 32592 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_295
timestamp 1751532312
transform 1 0 34384 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_303
timestamp 1751532423
transform 1 0 35280 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_313
timestamp 1751532440
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_330
timestamp 1751532312
transform 1 0 38304 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_338
timestamp 1751532246
transform 1 0 39200 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_346
timestamp 1751532440
transform 1 0 40096 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_350
timestamp 1751532351
transform 1 0 40544 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_366
timestamp 1751532351
transform 1 0 42336 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_382
timestamp 1751532440
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_2
timestamp 1751532440
transform 1 0 1568 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_4
timestamp 1751532423
transform 1 0 1792 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_32
timestamp 1751532440
transform 1 0 4928 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_36
timestamp 1751532440
transform 1 0 5376 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_38
timestamp 1751532423
transform 1 0 5600 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_52
timestamp 1751532351
transform 1 0 7168 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_68
timestamp 1751532440
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_72
timestamp 1751532351
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_88
timestamp 1751532351
transform 1 0 11200 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_104
timestamp 1751532246
transform 1 0 12992 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_108
timestamp 1751532423
transform 1 0 13440 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_120
timestamp 1751532440
transform 1 0 14784 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_124
timestamp 1751532351
transform 1 0 15232 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_142
timestamp 1751532351
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_158
timestamp 1751532440
transform 1 0 19040 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_170
timestamp 1751532351
transform 1 0 20384 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_186
timestamp 1751532246
transform 1 0 22176 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_190
timestamp 1751532440
transform 1 0 22624 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_204
timestamp 1751532246
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_208
timestamp 1751532440
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_212
timestamp 1751532351
transform 1 0 25088 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_228
timestamp 1751532351
transform 1 0 26880 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_244
timestamp 1751532351
transform 1 0 28672 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_260
timestamp 1751532351
transform 1 0 30464 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_276
timestamp 1751532246
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_282
timestamp 1751532312
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_290
timestamp 1751532440
transform 1 0 33824 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_292
timestamp 1751532423
transform 1 0 34048 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_299
timestamp 1751532351
transform 1 0 34832 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_315
timestamp 1751532351
transform 1 0 36624 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_331
timestamp 1751532351
transform 1 0 38416 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_347
timestamp 1751532440
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_349
timestamp 1751532423
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_352
timestamp 1751532351
transform 1 0 40768 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_368
timestamp 1751532351
transform 1 0 42560 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_2
timestamp 1751532351
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_18
timestamp 1751532351
transform 1 0 3360 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_34
timestamp 1751532423
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_37
timestamp 1751532351
transform 1 0 5488 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_53
timestamp 1751532351
transform 1 0 7280 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_79
timestamp 1751532423
transform 1 0 10192 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_86
timestamp 1751532351
transform 1 0 10976 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_102
timestamp 1751532440
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_104
timestamp 1751532423
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_107
timestamp 1751532440
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_109
timestamp 1751532423
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_124
timestamp 1751532351
transform 1 0 15232 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_28_140
timestamp 1751532312
transform 1 0 17024 0 1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_148
timestamp 1751532440
transform 1 0 17920 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_157
timestamp 1751532423
transform 1 0 18928 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_169
timestamp 1751532246
transform 1 0 20272 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_173
timestamp 1751532440
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_28_177
timestamp 1751532312
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_185
timestamp 1751532246
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_189
timestamp 1751532440
transform 1 0 22512 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_191
timestamp 1751532423
transform 1 0 22736 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_216
timestamp 1751532440
transform 1 0 25536 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_220
timestamp 1751532351
transform 1 0 25984 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_28_236
timestamp 1751532312
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_244
timestamp 1751532423
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_247
timestamp 1751532246
transform 1 0 29008 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_251
timestamp 1751532423
transform 1 0 29456 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_266
timestamp 1751532351
transform 1 0 31136 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_282
timestamp 1751532351
transform 1 0 32928 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_298
timestamp 1751532351
transform 1 0 34720 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_314
timestamp 1751532423
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_317
timestamp 1751532351
transform 1 0 36848 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_333
timestamp 1751532351
transform 1 0 38640 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_349
timestamp 1751532351
transform 1 0 40432 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_365
timestamp 1751532440
transform 1 0 42224 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_28_371
timestamp 1751532312
transform 1 0 42896 0 1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_28_379
timestamp 1751532246
transform 1 0 43792 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_383
timestamp 1751532423
transform 1 0 44240 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_2
timestamp 1751532351
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_18
timestamp 1751532351
transform 1 0 3360 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_34
timestamp 1751532351
transform 1 0 5152 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_50
timestamp 1751532351
transform 1 0 6944 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_66
timestamp 1751532246
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_82
timestamp 1751532351
transform 1 0 10528 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_98
timestamp 1751532312
transform 1 0 12320 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_106
timestamp 1751532440
transform 1 0 13216 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_115
timestamp 1751532440
transform 1 0 14224 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_127
timestamp 1751532312
transform 1 0 15568 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_135
timestamp 1751532246
transform 1 0 16464 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_139
timestamp 1751532423
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_142
timestamp 1751532246
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_146
timestamp 1751532440
transform 1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_148
timestamp 1751532423
transform 1 0 17920 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_166
timestamp 1751532351
transform 1 0 19936 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_182
timestamp 1751532246
transform 1 0 21728 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_186
timestamp 1751532440
transform 1 0 22176 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_188
timestamp 1751532423
transform 1 0 22400 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_193
timestamp 1751532312
transform 1 0 22960 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_201
timestamp 1751532440
transform 1 0 23856 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_203
timestamp 1751532423
transform 1 0 24080 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_206
timestamp 1751532246
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_212
timestamp 1751532351
transform 1 0 25088 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_228
timestamp 1751532312
transform 1 0 26880 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_236
timestamp 1751532440
transform 1 0 27776 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_238
timestamp 1751532423
transform 1 0 28000 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_264
timestamp 1751532440
transform 1 0 30912 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_268
timestamp 1751532312
transform 1 0 31360 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_276
timestamp 1751532246
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_282
timestamp 1751532312
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_290
timestamp 1751532423
transform 1 0 33824 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_297
timestamp 1751532312
transform 1 0 34608 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_305
timestamp 1751532246
transform 1 0 35504 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_309
timestamp 1751532440
transform 1 0 35952 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_311
timestamp 1751532423
transform 1 0 36176 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_318
timestamp 1751532423
transform 1 0 36960 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_325
timestamp 1751532351
transform 1 0 37744 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_341
timestamp 1751532246
transform 1 0 39536 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_345
timestamp 1751532440
transform 1 0 39984 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_347
timestamp 1751532423
transform 1 0 40208 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_352
timestamp 1751532440
transform 1 0 40768 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_354
timestamp 1751532423
transform 1 0 40992 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_382
timestamp 1751532440
transform 1 0 44128 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_2
timestamp 1751532351
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_18
timestamp 1751532351
transform 1 0 3360 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_34
timestamp 1751532423
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_37
timestamp 1751532246
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_41
timestamp 1751532423
transform 1 0 5936 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_56
timestamp 1751532351
transform 1 0 7616 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_72
timestamp 1751532351
transform 1 0 9408 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_88
timestamp 1751532351
transform 1 0 11200 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_104
timestamp 1751532423
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_107
timestamp 1751532312
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_122
timestamp 1751532440
transform 1 0 15008 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_126
timestamp 1751532351
transform 1 0 15456 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_142
timestamp 1751532312
transform 1 0 17248 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_150
timestamp 1751532246
transform 1 0 18144 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_154
timestamp 1751532440
transform 1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_158
timestamp 1751532351
transform 1 0 19040 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_174
timestamp 1751532423
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_183
timestamp 1751532246
transform 1 0 21840 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_187
timestamp 1751532440
transform 1 0 22288 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_201
timestamp 1751532351
transform 1 0 23856 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_217
timestamp 1751532351
transform 1 0 25648 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_233
timestamp 1751532246
transform 1 0 27440 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_237
timestamp 1751532423
transform 1 0 27888 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_247
timestamp 1751532440
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_260
timestamp 1751532351
transform 1 0 30464 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_276
timestamp 1751532351
transform 1 0 32256 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_292
timestamp 1751532246
transform 1 0 34048 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_296
timestamp 1751532440
transform 1 0 34496 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_298
timestamp 1751532423
transform 1 0 34720 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_311
timestamp 1751532440
transform 1 0 36176 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_329
timestamp 1751532246
transform 1 0 38192 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_333
timestamp 1751532440
transform 1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_335
timestamp 1751532423
transform 1 0 38864 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_352
timestamp 1751532440
transform 1 0 40768 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_364
timestamp 1751532351
transform 1 0 42112 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_380
timestamp 1751532246
transform 1 0 43904 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_2
timestamp 1751532351
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_18
timestamp 1751532246
transform 1 0 3360 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_36
timestamp 1751532440
transform 1 0 5376 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_40
timestamp 1751532440
transform 1 0 5824 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_44
timestamp 1751532351
transform 1 0 6272 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_60
timestamp 1751532312
transform 1 0 8064 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_68
timestamp 1751532440
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_72
timestamp 1751532246
transform 1 0 9408 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_87
timestamp 1751532351
transform 1 0 11088 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_103
timestamp 1751532246
transform 1 0 12880 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_107
timestamp 1751532440
transform 1 0 13328 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_123
timestamp 1751532351
transform 1 0 15120 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_139
timestamp 1751532423
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_153
timestamp 1751532440
transform 1 0 18480 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_157
timestamp 1751532351
transform 1 0 18928 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_173
timestamp 1751532351
transform 1 0 20720 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_189
timestamp 1751532351
transform 1 0 22512 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_205
timestamp 1751532440
transform 1 0 24304 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_207
timestamp 1751532423
transform 1 0 24528 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_212
timestamp 1751532440
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_214
timestamp 1751532423
transform 1 0 25312 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_229
timestamp 1751532351
transform 1 0 26992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_259
timestamp 1751532351
transform 1 0 30352 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_275
timestamp 1751532246
transform 1 0 32144 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_279
timestamp 1751532423
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_282
timestamp 1751532312
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_290
timestamp 1751532440
transform 1 0 33824 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_292
timestamp 1751532423
transform 1 0 34048 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_295
timestamp 1751532246
transform 1 0 34384 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_299
timestamp 1751532440
transform 1 0 34832 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_303
timestamp 1751532312
transform 1 0 35280 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_311
timestamp 1751532440
transform 1 0 36176 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_313
timestamp 1751532423
transform 1 0 36400 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_322
timestamp 1751532246
transform 1 0 37408 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_334
timestamp 1751532423
transform 1 0 38752 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_341
timestamp 1751532312
transform 1 0 39536 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_349
timestamp 1751532423
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_362
timestamp 1751532351
transform 1 0 41888 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_378
timestamp 1751532246
transform 1 0 43680 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_382
timestamp 1751532440
transform 1 0 44128 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_2
timestamp 1751532440
transform 1 0 1568 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_31
timestamp 1751532440
transform 1 0 4816 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_37
timestamp 1751532351
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_53
timestamp 1751532440
transform 1 0 7280 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_55
timestamp 1751532423
transform 1 0 7504 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_63
timestamp 1751532312
transform 1 0 8400 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_71
timestamp 1751532440
transform 1 0 9296 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_95
timestamp 1751532312
transform 1 0 11984 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_103
timestamp 1751532440
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_107
timestamp 1751532351
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_123
timestamp 1751532351
transform 1 0 15120 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_139
timestamp 1751532351
transform 1 0 16912 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_155
timestamp 1751532440
transform 1 0 18704 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_164
timestamp 1751532246
transform 1 0 19712 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_168
timestamp 1751532423
transform 1 0 20160 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_177
timestamp 1751532246
transform 1 0 21168 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_181
timestamp 1751532423
transform 1 0 21616 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_209
timestamp 1751532440
transform 1 0 24752 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_213
timestamp 1751532312
transform 1 0 25200 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_221
timestamp 1751532440
transform 1 0 26096 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_233
timestamp 1751532312
transform 1 0 27440 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_241
timestamp 1751532246
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_257
timestamp 1751532312
transform 1 0 30128 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_265
timestamp 1751532423
transform 1 0 31024 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_313
timestamp 1751532440
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_317
timestamp 1751532351
transform 1 0 36848 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_333
timestamp 1751532351
transform 1 0 38640 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_349
timestamp 1751532351
transform 1 0 40432 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_365
timestamp 1751532351
transform 1 0 42224 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_381
timestamp 1751532440
transform 1 0 44016 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_383
timestamp 1751532423
transform 1 0 44240 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_2
timestamp 1751532351
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_18
timestamp 1751532423
transform 1 0 3360 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_26
timestamp 1751532312
transform 1 0 4256 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_34
timestamp 1751532246
transform 1 0 5152 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_38
timestamp 1751532440
transform 1 0 5600 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_40
timestamp 1751532423
transform 1 0 5824 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_55
timestamp 1751532312
transform 1 0 7504 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_63
timestamp 1751532246
transform 1 0 8400 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_67
timestamp 1751532440
transform 1 0 8848 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_69
timestamp 1751532423
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_72
timestamp 1751532246
transform 1 0 9408 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_76
timestamp 1751532423
transform 1 0 9856 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_87
timestamp 1751532440
transform 1 0 11088 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_95
timestamp 1751532351
transform 1 0 11984 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_111
timestamp 1751532312
transform 1 0 13776 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_119
timestamp 1751532246
transform 1 0 14672 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_130
timestamp 1751532440
transform 1 0 15904 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_134
timestamp 1751532246
transform 1 0 16352 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_138
timestamp 1751532440
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_142
timestamp 1751532351
transform 1 0 17248 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_158
timestamp 1751532312
transform 1 0 19040 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_166
timestamp 1751532246
transform 1 0 19936 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_182
timestamp 1751532440
transform 1 0 21728 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_186
timestamp 1751532351
transform 1 0 22176 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_202
timestamp 1751532312
transform 1 0 23968 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_212
timestamp 1751532351
transform 1 0 25088 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_234
timestamp 1751532351
transform 1 0 27552 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_250
timestamp 1751532351
transform 1 0 29344 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_266
timestamp 1751532312
transform 1 0 31136 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_274
timestamp 1751532246
transform 1 0 32032 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_278
timestamp 1751532440
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_282
timestamp 1751532423
transform 1 0 32928 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_289
timestamp 1751532351
transform 1 0 33712 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_305
timestamp 1751532351
transform 1 0 35504 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_321
timestamp 1751532351
transform 1 0 37296 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_337
timestamp 1751532312
transform 1 0 39088 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_347
timestamp 1751532440
transform 1 0 40208 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_349
timestamp 1751532423
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_352
timestamp 1751532351
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_368
timestamp 1751532351
transform 1 0 42560 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_2
timestamp 1751532351
transform 1 0 1568 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_18
timestamp 1751532351
transform 1 0 3360 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_34
timestamp 1751532423
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_37
timestamp 1751532351
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_53
timestamp 1751532246
transform 1 0 7280 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_57
timestamp 1751532440
transform 1 0 7728 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_59
timestamp 1751532423
transform 1 0 7952 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_100
timestamp 1751532440
transform 1 0 12544 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_104
timestamp 1751532423
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_34_107
timestamp 1751532312
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_115
timestamp 1751532246
transform 1 0 14224 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_119
timestamp 1751532423
transform 1 0 14672 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_131
timestamp 1751532423
transform 1 0 16016 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_142
timestamp 1751532440
transform 1 0 17248 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_146
timestamp 1751532351
transform 1 0 17696 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_162
timestamp 1751532440
transform 1 0 19488 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_164
timestamp 1751532423
transform 1 0 19712 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_172
timestamp 1751532440
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_174
timestamp 1751532423
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_177
timestamp 1751532440
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_181
timestamp 1751532351
transform 1 0 21616 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_197
timestamp 1751532351
transform 1 0 23408 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_34_213
timestamp 1751532312
transform 1 0 25200 0 1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_221
timestamp 1751532440
transform 1 0 26096 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_223
timestamp 1751532423
transform 1 0 26320 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_34_235
timestamp 1751532312
transform 1 0 27664 0 1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_243
timestamp 1751532440
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_247
timestamp 1751532351
transform 1 0 29008 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_263
timestamp 1751532351
transform 1 0 30800 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_279
timestamp 1751532351
transform 1 0 32592 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_295
timestamp 1751532351
transform 1 0 34384 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_311
timestamp 1751532246
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_317
timestamp 1751532351
transform 1 0 36848 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_333
timestamp 1751532246
transform 1 0 38640 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_365
timestamp 1751532351
transform 1 0 42224 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_381
timestamp 1751532440
transform 1 0 44016 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_383
timestamp 1751532423
transform 1 0 44240 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_2
timestamp 1751532351
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_18
timestamp 1751532351
transform 1 0 3360 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_34
timestamp 1751532351
transform 1 0 5152 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_50
timestamp 1751532351
transform 1 0 6944 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_66
timestamp 1751532246
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_72
timestamp 1751532246
transform 1 0 9408 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_86
timestamp 1751532246
transform 1 0 10976 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_90
timestamp 1751532423
transform 1 0 11424 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_126
timestamp 1751532246
transform 1 0 15456 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_130
timestamp 1751532423
transform 1 0 15904 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_138
timestamp 1751532440
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_142
timestamp 1751532440
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_146
timestamp 1751532440
transform 1 0 17696 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_161
timestamp 1751532351
transform 1 0 19376 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_177
timestamp 1751532351
transform 1 0 21168 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_193
timestamp 1751532351
transform 1 0 22960 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_209
timestamp 1751532423
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_212
timestamp 1751532312
transform 1 0 25088 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_220
timestamp 1751532440
transform 1 0 25984 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_222
timestamp 1751532423
transform 1 0 26208 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_249
timestamp 1751532351
transform 1 0 29232 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_265
timestamp 1751532312
transform 1 0 31024 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_273
timestamp 1751532246
transform 1 0 31920 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_277
timestamp 1751532423
transform 1 0 32368 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_317
timestamp 1751532351
transform 1 0 36848 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_333
timestamp 1751532312
transform 1 0 38640 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_341
timestamp 1751532246
transform 1 0 39536 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_345
timestamp 1751532440
transform 1 0 39984 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_349
timestamp 1751532423
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_352
timestamp 1751532440
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_354
timestamp 1751532423
transform 1 0 40992 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_382
timestamp 1751532440
transform 1 0 44128 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_2
timestamp 1751532351
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_18
timestamp 1751532351
transform 1 0 3360 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_34
timestamp 1751532423
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_37
timestamp 1751532440
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_39
timestamp 1751532423
transform 1 0 5712 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_42
timestamp 1751532440
transform 1 0 6048 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_44
timestamp 1751532423
transform 1 0 6272 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_59
timestamp 1751532312
transform 1 0 7952 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_67
timestamp 1751532246
transform 1 0 8848 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_71
timestamp 1751532440
transform 1 0 9296 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_73
timestamp 1751532423
transform 1 0 9520 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_101
timestamp 1751532246
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_139
timestamp 1751532440
transform 1 0 16912 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_147
timestamp 1751532351
transform 1 0 17808 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_163
timestamp 1751532312
transform 1 0 19600 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_171
timestamp 1751532246
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_177
timestamp 1751532312
transform 1 0 21168 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_185
timestamp 1751532440
transform 1 0 22064 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_187
timestamp 1751532423
transform 1 0 22288 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_194
timestamp 1751532440
transform 1 0 23072 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_198
timestamp 1751532351
transform 1 0 23520 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_214
timestamp 1751532246
transform 1 0 25312 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_222
timestamp 1751532312
transform 1 0 26208 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_230
timestamp 1751532246
transform 1 0 27104 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_234
timestamp 1751532423
transform 1 0 27552 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_237
timestamp 1751532440
transform 1 0 27888 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_36_272
timestamp 1751532312
transform 1 0 31808 0 1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_280
timestamp 1751532246
transform 1 0 32704 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_284
timestamp 1751532440
transform 1 0 33152 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_321
timestamp 1751532351
transform 1 0 37296 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_337
timestamp 1751532351
transform 1 0 39088 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_365
timestamp 1751532351
transform 1 0 42224 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_381
timestamp 1751532440
transform 1 0 44016 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_383
timestamp 1751532423
transform 1 0 44240 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_2
timestamp 1751532351
transform 1 0 1568 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_18
timestamp 1751532246
transform 1 0 3360 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_22
timestamp 1751532440
transform 1 0 3808 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_38
timestamp 1751532423
transform 1 0 5600 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_50
timestamp 1751532440
transform 1 0 6944 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_54
timestamp 1751532351
transform 1 0 7392 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_72
timestamp 1751532351
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_88
timestamp 1751532351
transform 1 0 11200 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_104
timestamp 1751532351
transform 1 0 12992 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_120
timestamp 1751532312
transform 1 0 14784 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_128
timestamp 1751532246
transform 1 0 15680 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_134
timestamp 1751532246
transform 1 0 16352 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_138
timestamp 1751532440
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_142
timestamp 1751532351
transform 1 0 17248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_158
timestamp 1751532351
transform 1 0 19040 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_174
timestamp 1751532312
transform 1 0 20832 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_182
timestamp 1751532423
transform 1 0 21728 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_212
timestamp 1751532440
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_216
timestamp 1751532351
transform 1 0 25536 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_232
timestamp 1751532312
transform 1 0 27328 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_240
timestamp 1751532440
transform 1 0 28224 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_242
timestamp 1751532423
transform 1 0 28448 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_270
timestamp 1751532440
transform 1 0 31584 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_274
timestamp 1751532246
transform 1 0 32032 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_278
timestamp 1751532440
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_282
timestamp 1751532351
transform 1 0 32928 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_37_298
timestamp 1751532312
transform 1 0 34720 0 -1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_306
timestamp 1751532246
transform 1 0 35616 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_310
timestamp 1751532423
transform 1 0 36064 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_327
timestamp 1751532351
transform 1 0 37968 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_343
timestamp 1751532246
transform 1 0 39760 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_347
timestamp 1751532440
transform 1 0 40208 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_37_349
timestamp 1751532423
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_37_362
timestamp 1751532351
transform 1 0 41888 0 -1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_37_378
timestamp 1751532246
transform 1 0 43680 0 -1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_37_382
timestamp 1751532440
transform 1 0 44128 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_2
timestamp 1751532440
transform 1 0 1568 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_31
timestamp 1751532440
transform 1 0 4816 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_38_51
timestamp 1751532312
transform 1 0 7056 0 1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_59
timestamp 1751532440
transform 1 0 7952 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_67
timestamp 1751532351
transform 1 0 8848 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_83
timestamp 1751532351
transform 1 0 10640 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_99
timestamp 1751532246
transform 1 0 12432 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_103
timestamp 1751532440
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_107
timestamp 1751532351
transform 1 0 13328 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_123
timestamp 1751532351
transform 1 0 15120 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_38_139
timestamp 1751532312
transform 1 0 16912 0 1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_147
timestamp 1751532440
transform 1 0 17808 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_159
timestamp 1751532440
transform 1 0 19152 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_38_163
timestamp 1751532312
transform 1 0 19600 0 1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_171
timestamp 1751532246
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_177
timestamp 1751532246
transform 1 0 21168 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_187
timestamp 1751532440
transform 1 0 22288 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_191
timestamp 1751532246
transform 1 0 22736 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_210
timestamp 1751532351
transform 1 0 24864 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_226
timestamp 1751532351
transform 1 0 26656 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_242
timestamp 1751532440
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_244
timestamp 1751532423
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_247
timestamp 1751532440
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_256
timestamp 1751532351
transform 1 0 30016 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_272
timestamp 1751532246
transform 1 0 31808 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_276
timestamp 1751532440
transform 1 0 32256 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_284
timestamp 1751532351
transform 1 0 33152 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_38_300
timestamp 1751532312
transform 1 0 34944 0 1 32928
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_38_308
timestamp 1751532246
transform 1 0 35840 0 1 32928
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_312
timestamp 1751532440
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_314
timestamp 1751532423
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_317
timestamp 1751532351
transform 1 0 36848 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_333
timestamp 1751532351
transform 1 0 38640 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_349
timestamp 1751532351
transform 1 0 40432 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_38_365
timestamp 1751532351
transform 1 0 42224 0 1 32928
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_38_381
timestamp 1751532440
transform 1 0 44016 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_38_383
timestamp 1751532423
transform 1 0 44240 0 1 32928
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_2
timestamp 1751532312
transform 1 0 1568 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_10
timestamp 1751532246
transform 1 0 2464 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_14
timestamp 1751532423
transform 1 0 2912 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_22
timestamp 1751532312
transform 1 0 3808 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_44
timestamp 1751532351
transform 1 0 6272 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_60
timestamp 1751532312
transform 1 0 8064 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_68
timestamp 1751532440
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_72
timestamp 1751532351
transform 1 0 9408 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_88
timestamp 1751532351
transform 1 0 11200 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_104
timestamp 1751532246
transform 1 0 12992 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_108
timestamp 1751532440
transform 1 0 13440 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_121
timestamp 1751532440
transform 1 0 14896 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_125
timestamp 1751532246
transform 1 0 15344 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_129
timestamp 1751532423
transform 1 0 15792 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_166
timestamp 1751532440
transform 1 0 19936 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_170
timestamp 1751532246
transform 1 0 20384 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_174
timestamp 1751532440
transform 1 0 20832 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_176
timestamp 1751532423
transform 1 0 21056 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_185
timestamp 1751532440
transform 1 0 22064 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_191
timestamp 1751532440
transform 1 0 22736 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_195
timestamp 1751532423
transform 1 0 23184 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_202
timestamp 1751532312
transform 1 0 23968 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_212
timestamp 1751532351
transform 1 0 25088 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_228
timestamp 1751532440
transform 1 0 26880 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_230
timestamp 1751532423
transform 1 0 27104 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_244
timestamp 1751532312
transform 1 0 28672 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_252
timestamp 1751532440
transform 1 0 29568 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_254
timestamp 1751532423
transform 1 0 29792 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_39_265
timestamp 1751532312
transform 1 0 31024 0 -1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_273
timestamp 1751532246
transform 1 0 31920 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_39_277
timestamp 1751532440
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_279
timestamp 1751532423
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_282
timestamp 1751532351
transform 1 0 32928 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_298
timestamp 1751532246
transform 1 0 34720 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_302
timestamp 1751532423
transform 1 0 35168 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_313
timestamp 1751532351
transform 1 0 36400 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_329
timestamp 1751532351
transform 1 0 38192 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_39_345
timestamp 1751532246
transform 1 0 39984 0 -1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_39_349
timestamp 1751532423
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_352
timestamp 1751532351
transform 1 0 40768 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_39_368
timestamp 1751532351
transform 1 0 42560 0 -1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_2
timestamp 1751532351
transform 1 0 1568 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_18
timestamp 1751532351
transform 1 0 3360 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_34
timestamp 1751532423
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_48
timestamp 1751532440
transform 1 0 6720 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_52
timestamp 1751532351
transform 1 0 7168 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_68
timestamp 1751532351
transform 1 0 8960 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_84
timestamp 1751532351
transform 1 0 10752 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_100
timestamp 1751532246
transform 1 0 12544 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_104
timestamp 1751532423
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_107
timestamp 1751532246
transform 1 0 13328 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_111
timestamp 1751532423
transform 1 0 13776 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_126
timestamp 1751532312
transform 1 0 15456 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_134
timestamp 1751532423
transform 1 0 16352 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_149
timestamp 1751532440
transform 1 0 18032 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_151
timestamp 1751532423
transform 1 0 18256 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_162
timestamp 1751532312
transform 1 0 19488 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_170
timestamp 1751532246
transform 1 0 20384 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_174
timestamp 1751532423
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_177
timestamp 1751532351
transform 1 0 21168 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_193
timestamp 1751532351
transform 1 0 22960 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_221
timestamp 1751532246
transform 1 0 26096 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_225
timestamp 1751532423
transform 1 0 26544 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_230
timestamp 1751532423
transform 1 0 27104 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_261
timestamp 1751532351
transform 1 0 30576 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_277
timestamp 1751532351
transform 1 0 32368 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_40_293
timestamp 1751532351
transform 1 0 34160 0 1 34496
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_309
timestamp 1751532423
transform 1 0 35952 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_314
timestamp 1751532423
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_317
timestamp 1751532440
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_321
timestamp 1751532312
transform 1 0 37296 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_329
timestamp 1751532423
transform 1 0 38192 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_340
timestamp 1751532423
transform 1 0 39424 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_40_351
timestamp 1751532440
transform 1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_363
timestamp 1751532246
transform 1 0 42000 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_40_371
timestamp 1751532312
transform 1 0 42896 0 1 34496
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_40_379
timestamp 1751532246
transform 1 0 43792 0 1 34496
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_40_383
timestamp 1751532423
transform 1 0 44240 0 1 34496
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_2
timestamp 1751532351
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_18
timestamp 1751532351
transform 1 0 3360 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_34
timestamp 1751532312
transform 1 0 5152 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_42
timestamp 1751532440
transform 1 0 6048 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_50
timestamp 1751532351
transform 1 0 6944 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_66
timestamp 1751532246
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_86
timestamp 1751532246
transform 1 0 10976 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_96
timestamp 1751532312
transform 1 0 12096 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_104
timestamp 1751532440
transform 1 0 12992 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_122
timestamp 1751532351
transform 1 0 15008 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_138
timestamp 1751532440
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_142
timestamp 1751532312
transform 1 0 17248 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_150
timestamp 1751532440
transform 1 0 18144 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_158
timestamp 1751532351
transform 1 0 19040 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_174
timestamp 1751532351
transform 1 0 20832 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_190
timestamp 1751532351
transform 1 0 22624 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_206
timestamp 1751532246
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_212
timestamp 1751532351
transform 1 0 25088 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_228
timestamp 1751532312
transform 1 0 26880 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_236
timestamp 1751532246
transform 1 0 27776 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_240
timestamp 1751532440
transform 1 0 28224 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_242
timestamp 1751532423
transform 1 0 28448 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_41_260
timestamp 1751532351
transform 1 0 30464 0 -1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_41_276
timestamp 1751532246
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_41_282
timestamp 1751532312
transform 1 0 32928 0 -1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_290
timestamp 1751532423
transform 1 0 33824 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_332
timestamp 1751532440
transform 1 0 38528 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_352
timestamp 1751532440
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_41_354
timestamp 1751532423
transform 1 0 40992 0 -1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_41_382
timestamp 1751532440
transform 1 0 44128 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_2
timestamp 1751532351
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_18
timestamp 1751532351
transform 1 0 3360 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_34
timestamp 1751532423
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_37
timestamp 1751532312
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_45
timestamp 1751532423
transform 1 0 6384 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_73
timestamp 1751532440
transform 1 0 9520 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_75
timestamp 1751532423
transform 1 0 9744 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_103
timestamp 1751532440
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_107
timestamp 1751532351
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_123
timestamp 1751532351
transform 1 0 15120 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_139
timestamp 1751532312
transform 1 0 16912 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_147
timestamp 1751532246
transform 1 0 17808 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_151
timestamp 1751532423
transform 1 0 18256 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_154
timestamp 1751532246
transform 1 0 18592 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_158
timestamp 1751532423
transform 1 0 19040 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_165
timestamp 1751532312
transform 1 0 19824 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_173
timestamp 1751532440
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_177
timestamp 1751532351
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_193
timestamp 1751532351
transform 1 0 22960 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_219
timestamp 1751532351
transform 1 0 25872 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_235
timestamp 1751532312
transform 1 0 27664 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_243
timestamp 1751532440
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_247
timestamp 1751532351
transform 1 0 29008 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_290
timestamp 1751532440
transform 1 0 33824 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_294
timestamp 1751532351
transform 1 0 34272 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_310
timestamp 1751532246
transform 1 0 36064 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_314
timestamp 1751532423
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_317
timestamp 1751532440
transform 1 0 36848 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_321
timestamp 1751532351
transform 1 0 37296 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_42_337
timestamp 1751532246
transform 1 0 39088 0 1 36064
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_341
timestamp 1751532440
transform 1 0 39536 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_42_343
timestamp 1751532423
transform 1 0 39760 0 1 36064
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_354
timestamp 1751532440
transform 1 0 40992 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_42_358
timestamp 1751532351
transform 1 0 41440 0 1 36064
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_42_374
timestamp 1751532312
transform 1 0 43232 0 1 36064
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_42_382
timestamp 1751532440
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_2
timestamp 1751532351
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_18
timestamp 1751532440
transform 1 0 3360 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_20
timestamp 1751532423
transform 1 0 3584 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_31
timestamp 1751532440
transform 1 0 4816 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_35
timestamp 1751532351
transform 1 0 5264 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_51
timestamp 1751532351
transform 1 0 7056 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_67
timestamp 1751532440
transform 1 0 8848 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_69
timestamp 1751532423
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_72
timestamp 1751532440
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_76
timestamp 1751532351
transform 1 0 9856 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_92
timestamp 1751532351
transform 1 0 11648 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_108
timestamp 1751532351
transform 1 0 13440 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_124
timestamp 1751532351
transform 1 0 15232 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_179
timestamp 1751532440
transform 1 0 21392 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_183
timestamp 1751532351
transform 1 0 21840 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_43_199
timestamp 1751532312
transform 1 0 23632 0 -1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_207
timestamp 1751532440
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_209
timestamp 1751532423
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_43_212
timestamp 1751532440
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_228
timestamp 1751532246
transform 1 0 26880 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_43_232
timestamp 1751532423
transform 1 0 27328 0 -1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_240
timestamp 1751532351
transform 1 0 28224 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_256
timestamp 1751532351
transform 1 0 30016 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_43_272
timestamp 1751532312
transform 1 0 31808 0 -1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_282
timestamp 1751532351
transform 1 0 32928 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_298
timestamp 1751532351
transform 1 0 34720 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_314
timestamp 1751532351
transform 1 0 36512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_330
timestamp 1751532351
transform 1 0 38304 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_346
timestamp 1751532246
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_43_356
timestamp 1751532351
transform 1 0 41216 0 -1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_43_372
timestamp 1751532312
transform 1 0 43008 0 -1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_43_380
timestamp 1751532246
transform 1 0 43904 0 -1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_2
timestamp 1751532351
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_18
timestamp 1751532440
transform 1 0 3360 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_20
timestamp 1751532423
transform 1 0 3584 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_31
timestamp 1751532440
transform 1 0 4816 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_37
timestamp 1751532351
transform 1 0 5488 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_53
timestamp 1751532351
transform 1 0 7280 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_69
timestamp 1751532351
transform 1 0 9072 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_85
timestamp 1751532351
transform 1 0 10864 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_101
timestamp 1751532246
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_107
timestamp 1751532351
transform 1 0 13328 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_123
timestamp 1751532351
transform 1 0 15120 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_139
timestamp 1751532351
transform 1 0 16912 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_155
timestamp 1751532351
transform 1 0 18704 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_171
timestamp 1751532246
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_177
timestamp 1751532351
transform 1 0 21168 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_193
timestamp 1751532440
transform 1 0 22960 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_205
timestamp 1751532351
transform 1 0 24304 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_221
timestamp 1751532351
transform 1 0 26096 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_44_237
timestamp 1751532312
transform 1 0 27888 0 1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_260
timestamp 1751532351
transform 1 0 30464 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_276
timestamp 1751532351
transform 1 0 32256 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_292
timestamp 1751532351
transform 1 0 34048 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_308
timestamp 1751532246
transform 1 0 35840 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_312
timestamp 1751532440
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_314
timestamp 1751532423
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_44_317
timestamp 1751532351
transform 1 0 36848 0 1 37632
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_333
timestamp 1751532246
transform 1 0 38640 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_337
timestamp 1751532440
transform 1 0 39088 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_339
timestamp 1751532423
transform 1 0 39312 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_44_369
timestamp 1751532312
transform 1 0 42672 0 1 37632
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_44_377
timestamp 1751532246
transform 1 0 43568 0 1 37632
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_44_381
timestamp 1751532440
transform 1 0 44016 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_44_383
timestamp 1751532423
transform 1 0 44240 0 1 37632
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_2
timestamp 1751532312
transform 1 0 1568 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_10
timestamp 1751532423
transform 1 0 2464 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_38
timestamp 1751532351
transform 1 0 5600 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_54
timestamp 1751532423
transform 1 0 7392 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_61
timestamp 1751532312
transform 1 0 8176 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_69
timestamp 1751532423
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_72
timestamp 1751532351
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_88
timestamp 1751532351
transform 1 0 11200 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_104
timestamp 1751532246
transform 1 0 12992 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_114
timestamp 1751532312
transform 1 0 14112 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_122
timestamp 1751532246
transform 1 0 15008 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_126
timestamp 1751532440
transform 1 0 15456 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_128
timestamp 1751532423
transform 1 0 15680 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_135
timestamp 1751532246
transform 1 0 16464 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_139
timestamp 1751532423
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_142
timestamp 1751532351
transform 1 0 17248 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_158
timestamp 1751532351
transform 1 0 19040 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_174
timestamp 1751532351
transform 1 0 20832 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_190
timestamp 1751532312
transform 1 0 22624 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_208
timestamp 1751532440
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_212
timestamp 1751532351
transform 1 0 25088 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_228
timestamp 1751532312
transform 1 0 26880 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_236
timestamp 1751532246
transform 1 0 27776 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_247
timestamp 1751532351
transform 1 0 29008 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_263
timestamp 1751532351
transform 1 0 30800 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_279
timestamp 1751532423
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_282
timestamp 1751532351
transform 1 0 32928 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_298
timestamp 1751532312
transform 1 0 34720 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_306
timestamp 1751532423
transform 1 0 35616 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_319
timestamp 1751532351
transform 1 0 37072 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_45_335
timestamp 1751532312
transform 1 0 38864 0 -1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_45_343
timestamp 1751532246
transform 1 0 39760 0 -1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_45_347
timestamp 1751532440
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_45_349
timestamp 1751532423
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_352
timestamp 1751532351
transform 1 0 40768 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_45_368
timestamp 1751532351
transform 1 0 42560 0 -1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_2
timestamp 1751532351
transform 1 0 1568 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_18
timestamp 1751532312
transform 1 0 3360 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_26
timestamp 1751532440
transform 1 0 4256 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_37
timestamp 1751532351
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_53
timestamp 1751532312
transform 1 0 7280 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_61
timestamp 1751532440
transform 1 0 8176 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_63
timestamp 1751532423
transform 1 0 8400 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_107
timestamp 1751532440
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_109
timestamp 1751532423
transform 1 0 13552 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_116
timestamp 1751532312
transform 1 0 14336 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_124
timestamp 1751532440
transform 1 0 15232 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_126
timestamp 1751532423
transform 1 0 15456 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_154
timestamp 1751532312
transform 1 0 18592 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_162
timestamp 1751532246
transform 1 0 19488 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_172
timestamp 1751532440
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_174
timestamp 1751532423
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_177
timestamp 1751532351
transform 1 0 21168 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_193
timestamp 1751532440
transform 1 0 22960 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_195
timestamp 1751532423
transform 1 0 23184 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_209
timestamp 1751532351
transform 1 0 24752 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_225
timestamp 1751532351
transform 1 0 26544 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_241
timestamp 1751532246
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_254
timestamp 1751532423
transform 1 0 29792 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_261
timestamp 1751532351
transform 1 0 30576 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_277
timestamp 1751532423
transform 1 0 32368 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_284
timestamp 1751532351
transform 1 0 33152 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_300
timestamp 1751532312
transform 1 0 34944 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_308
timestamp 1751532440
transform 1 0 35840 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_312
timestamp 1751532440
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_314
timestamp 1751532423
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_46_323
timestamp 1751532351
transform 1 0 37520 0 1 39200
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_339
timestamp 1751532312
transform 1 0 39312 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_46_347
timestamp 1751532246
transform 1 0 40208 0 1 39200
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_357
timestamp 1751532312
transform 1 0 41328 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_46_365
timestamp 1751532423
transform 1 0 42224 0 1 39200
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_46_372
timestamp 1751532440
transform 1 0 43008 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_46_376
timestamp 1751532312
transform 1 0 43456 0 1 39200
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_2
timestamp 1751532246
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_6
timestamp 1751532423
transform 1 0 2016 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_34
timestamp 1751532440
transform 1 0 5152 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_38
timestamp 1751532423
transform 1 0 5600 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_66
timestamp 1751532440
transform 1 0 8736 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_72
timestamp 1751532351
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_88
timestamp 1751532440
transform 1 0 11200 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_90
timestamp 1751532423
transform 1 0 11424 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_47_118
timestamp 1751532351
transform 1 0 14560 0 -1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_134
timestamp 1751532246
transform 1 0 16352 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_138
timestamp 1751532440
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_47_142
timestamp 1751532312
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_150
timestamp 1751532440
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_179
timestamp 1751532246
transform 1 0 21392 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_212
timestamp 1751532440
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_216
timestamp 1751532246
transform 1 0 25536 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_247
timestamp 1751532440
transform 1 0 29008 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_251
timestamp 1751532440
transform 1 0 29456 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_282
timestamp 1751532440
transform 1 0 32928 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_284
timestamp 1751532423
transform 1 0 33152 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_47_345
timestamp 1751532440
transform 1 0 39984 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_347
timestamp 1751532423
transform 1 0 40208 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_47_379
timestamp 1751532246
transform 1 0 43792 0 -1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_47_383
timestamp 1751532423
transform 1 0 44240 0 -1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_2
timestamp 1751532351
transform 1 0 1568 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_18
timestamp 1751532351
transform 1 0 3360 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_34
timestamp 1751532423
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_37
timestamp 1751532351
transform 1 0 5488 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_53
timestamp 1751532351
transform 1 0 7280 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_69
timestamp 1751532351
transform 1 0 9072 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_85
timestamp 1751532351
transform 1 0 10864 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_101
timestamp 1751532246
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_107
timestamp 1751532351
transform 1 0 13328 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_123
timestamp 1751532351
transform 1 0 15120 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_139
timestamp 1751532351
transform 1 0 16912 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_155
timestamp 1751532351
transform 1 0 18704 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_171
timestamp 1751532246
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_177
timestamp 1751532351
transform 1 0 21168 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_193
timestamp 1751532351
transform 1 0 22960 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_209
timestamp 1751532351
transform 1 0 24752 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_225
timestamp 1751532351
transform 1 0 26544 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_241
timestamp 1751532246
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_247
timestamp 1751532351
transform 1 0 29008 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_263
timestamp 1751532351
transform 1 0 30800 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_279
timestamp 1751532423
transform 1 0 32592 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_282
timestamp 1751532351
transform 1 0 32928 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_48_298
timestamp 1751532312
transform 1 0 34720 0 1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_48_306
timestamp 1751532246
transform 1 0 35616 0 1 40768
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_310
timestamp 1751532440
transform 1 0 36064 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_48_314
timestamp 1751532423
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_317
timestamp 1751532351
transform 1 0 36848 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_48_333
timestamp 1751532351
transform 1 0 38640 0 1 40768
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_48_349
timestamp 1751532312
transform 1 0 40432 0 1 40768
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_48_357
timestamp 1751532440
transform 1 0 41328 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_2
timestamp 1751532351
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_49_18
timestamp 1751532312
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_26
timestamp 1751532246
transform 1 0 4256 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_30
timestamp 1751532440
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_36
timestamp 1751532440
transform 1 0 5376 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_38
timestamp 1751532423
transform 1 0 5600 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_45
timestamp 1751532351
transform 1 0 6384 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_61
timestamp 1751532246
transform 1 0 8176 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_65
timestamp 1751532423
transform 1 0 8624 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_70
timestamp 1751532440
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_72
timestamp 1751532423
transform 1 0 9408 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_49_79
timestamp 1751532351
transform 1 0 10192 0 -1 42336
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_95
timestamp 1751532246
transform 1 0 11984 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_99
timestamp 1751532440
transform 1 0 12432 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_101
timestamp 1751532423
transform 1 0 12656 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_104
timestamp 1751532440
transform 1 0 12992 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_106
timestamp 1751532423
transform 1 0 13216 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_132
timestamp 1751532246
transform 1 0 16128 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_138
timestamp 1751532440
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_140
timestamp 1751532423
transform 1 0 17024 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_166
timestamp 1751532246
transform 1 0 19936 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_172
timestamp 1751532440
transform 1 0 20608 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_174
timestamp 1751532423
transform 1 0 20832 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_200
timestamp 1751532246
transform 1 0 23744 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_206
timestamp 1751532440
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_208
timestamp 1751532423
transform 1 0 24640 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_234
timestamp 1751532246
transform 1 0 27552 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_240
timestamp 1751532440
transform 1 0 28224 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_242
timestamp 1751532423
transform 1 0 28448 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_268
timestamp 1751532246
transform 1 0 31360 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_274
timestamp 1751532440
transform 1 0 32032 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_276
timestamp 1751532423
transform 1 0 32256 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_302
timestamp 1751532246
transform 1 0 35168 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_308
timestamp 1751532440
transform 1 0 35840 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_310
timestamp 1751532423
transform 1 0 36064 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_336
timestamp 1751532246
transform 1 0 38976 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_49_342
timestamp 1751532440
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_49_344
timestamp 1751532423
transform 1 0 39872 0 -1 42336
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_49_370
timestamp 1751532246
transform 1 0 42784 0 -1 42336
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_49_376
timestamp 1751532312
transform 1 0 43456 0 -1 42336
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform 1 0 9520 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input2
timestamp 1751534193
transform 1 0 5712 0 -1 42336
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output3
timestamp 1751661108
transform 1 0 13328 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output4
timestamp 1751661108
transform 1 0 17136 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output5
timestamp 1751661108
transform 1 0 20944 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output6
timestamp 1751661108
transform 1 0 24752 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output7
timestamp 1751661108
transform 1 0 28560 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output8
timestamp 1751661108
transform 1 0 32368 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output9
timestamp 1751661108
transform 1 0 36176 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output10
timestamp 1751661108
transform 1 0 39984 0 -1 42336
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output11
timestamp 1751661108
transform 1 0 41552 0 1 40768
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_50 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 44576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_51
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 44576 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_52
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 44576 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_53
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_54
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 44576 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_55
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_56
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 44576 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_57
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_58
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 44576 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_59
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_60
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 44576 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_61
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 44576 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_62
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 44576 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_63
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 44576 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_64
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 44576 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_65
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_66
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 44576 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_67
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_68
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 44576 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_69
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_70
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 44576 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_71
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Left_72
timestamp 1751532504
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Right_22
timestamp 1751532504
transform -1 0 44576 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Left_73
timestamp 1751532504
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Right_23
timestamp 1751532504
transform -1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Left_74
timestamp 1751532504
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Right_24
timestamp 1751532504
transform -1 0 44576 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Left_75
timestamp 1751532504
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Right_25
timestamp 1751532504
transform -1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Left_76
timestamp 1751532504
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Right_26
timestamp 1751532504
transform -1 0 44576 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Left_77
timestamp 1751532504
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Right_27
timestamp 1751532504
transform -1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Left_78
timestamp 1751532504
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Right_28
timestamp 1751532504
transform -1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Left_79
timestamp 1751532504
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Right_29
timestamp 1751532504
transform -1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Left_80
timestamp 1751532504
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Right_30
timestamp 1751532504
transform -1 0 44576 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Left_81
timestamp 1751532504
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Right_31
timestamp 1751532504
transform -1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Left_82
timestamp 1751532504
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Right_32
timestamp 1751532504
transform -1 0 44576 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Left_83
timestamp 1751532504
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Right_33
timestamp 1751532504
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Left_84
timestamp 1751532504
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Right_34
timestamp 1751532504
transform -1 0 44576 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Left_85
timestamp 1751532504
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Right_35
timestamp 1751532504
transform -1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Left_86
timestamp 1751532504
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Right_36
timestamp 1751532504
transform -1 0 44576 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Left_87
timestamp 1751532504
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_37_Right_37
timestamp 1751532504
transform -1 0 44576 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Left_88
timestamp 1751532504
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_38_Right_38
timestamp 1751532504
transform -1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Left_89
timestamp 1751532504
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_39_Right_39
timestamp 1751532504
transform -1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Left_90
timestamp 1751532504
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_40_Right_40
timestamp 1751532504
transform -1 0 44576 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Left_91
timestamp 1751532504
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_41_Right_41
timestamp 1751532504
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Left_92
timestamp 1751532504
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_42_Right_42
timestamp 1751532504
transform -1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Left_93
timestamp 1751532504
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_43_Right_43
timestamp 1751532504
transform -1 0 44576 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Left_94
timestamp 1751532504
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_44_Right_44
timestamp 1751532504
transform -1 0 44576 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Left_95
timestamp 1751532504
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_45_Right_45
timestamp 1751532504
transform -1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Left_96
timestamp 1751532504
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_46_Right_46
timestamp 1751532504
transform -1 0 44576 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Left_97
timestamp 1751532504
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_47_Right_47
timestamp 1751532504
transform -1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Left_98
timestamp 1751532504
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_48_Right_48
timestamp 1751532504
transform -1 0 44576 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Left_99
timestamp 1751532504
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_49_Right_49
timestamp 1751532504
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_100
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_101
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_102
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_103
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_104
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_105
timestamp 1751532504
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_106
timestamp 1751532504
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_107
timestamp 1751532504
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_108
timestamp 1751532504
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_109
timestamp 1751532504
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_110
timestamp 1751532504
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_111
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_112
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_113
timestamp 1751532504
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_114
timestamp 1751532504
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_115
timestamp 1751532504
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_116
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_117
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_118
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_119
timestamp 1751532504
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_120
timestamp 1751532504
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_121
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_122
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_123
timestamp 1751532504
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_124
timestamp 1751532504
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_125
timestamp 1751532504
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_126
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_127
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_128
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_129
timestamp 1751532504
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_130
timestamp 1751532504
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_131
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_132
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_133
timestamp 1751532504
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_134
timestamp 1751532504
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_135
timestamp 1751532504
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_136
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_137
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_138
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_139
timestamp 1751532504
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_140
timestamp 1751532504
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_141
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_142
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_143
timestamp 1751532504
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_144
timestamp 1751532504
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_145
timestamp 1751532504
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_146
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_147
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_148
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_149
timestamp 1751532504
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_150
timestamp 1751532504
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_151
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_152
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_153
timestamp 1751532504
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_154
timestamp 1751532504
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_155
timestamp 1751532504
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_156
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_157
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_158
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_159
timestamp 1751532504
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_160
timestamp 1751532504
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_161
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_162
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_163
timestamp 1751532504
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_164
timestamp 1751532504
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_165
timestamp 1751532504
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_166
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_167
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_168
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_169
timestamp 1751532504
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_170
timestamp 1751532504
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_171
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_172
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_173
timestamp 1751532504
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_174
timestamp 1751532504
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_175
timestamp 1751532504
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_176
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_177
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_178
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_179
timestamp 1751532504
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_180
timestamp 1751532504
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_181
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_182
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_183
timestamp 1751532504
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_184
timestamp 1751532504
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_185
timestamp 1751532504
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_186
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_187
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_188
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_189
timestamp 1751532504
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_190
timestamp 1751532504
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_191
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_192
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_193
timestamp 1751532504
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_194
timestamp 1751532504
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_195
timestamp 1751532504
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_196
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_197
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_198
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_199
timestamp 1751532504
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_200
timestamp 1751532504
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_201
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_202
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_203
timestamp 1751532504
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_204
timestamp 1751532504
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_205
timestamp 1751532504
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_206
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_207
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_208
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_209
timestamp 1751532504
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_210
timestamp 1751532504
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_211
timestamp 1751532504
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_212
timestamp 1751532504
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_213
timestamp 1751532504
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_214
timestamp 1751532504
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_215
timestamp 1751532504
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_216
timestamp 1751532504
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_217
timestamp 1751532504
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_218
timestamp 1751532504
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_219
timestamp 1751532504
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_220
timestamp 1751532504
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_221
timestamp 1751532504
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_222
timestamp 1751532504
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_223
timestamp 1751532504
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_224
timestamp 1751532504
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_225
timestamp 1751532504
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_226
timestamp 1751532504
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_227
timestamp 1751532504
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_228
timestamp 1751532504
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_229
timestamp 1751532504
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_230
timestamp 1751532504
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_231
timestamp 1751532504
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_232
timestamp 1751532504
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_233
timestamp 1751532504
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_234
timestamp 1751532504
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_235
timestamp 1751532504
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_236
timestamp 1751532504
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_237
timestamp 1751532504
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_238
timestamp 1751532504
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_239
timestamp 1751532504
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_240
timestamp 1751532504
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_241
timestamp 1751532504
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_242
timestamp 1751532504
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_243
timestamp 1751532504
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_244
timestamp 1751532504
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_245
timestamp 1751532504
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_246
timestamp 1751532504
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_247
timestamp 1751532504
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_248
timestamp 1751532504
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_249
timestamp 1751532504
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_250
timestamp 1751532504
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_251
timestamp 1751532504
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_252
timestamp 1751532504
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_253
timestamp 1751532504
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_254
timestamp 1751532504
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_255
timestamp 1751532504
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_256
timestamp 1751532504
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_257
timestamp 1751532504
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_258
timestamp 1751532504
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_259
timestamp 1751532504
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_260
timestamp 1751532504
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_261
timestamp 1751532504
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_262
timestamp 1751532504
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_263
timestamp 1751532504
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_264
timestamp 1751532504
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_265
timestamp 1751532504
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_266
timestamp 1751532504
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_267
timestamp 1751532504
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_268
timestamp 1751532504
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_269
timestamp 1751532504
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_270
timestamp 1751532504
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_271
timestamp 1751532504
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_272
timestamp 1751532504
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_273
timestamp 1751532504
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_274
timestamp 1751532504
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_275
timestamp 1751532504
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_276
timestamp 1751532504
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_277
timestamp 1751532504
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_278
timestamp 1751532504
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_279
timestamp 1751532504
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_280
timestamp 1751532504
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_281
timestamp 1751532504
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_282
timestamp 1751532504
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_283
timestamp 1751532504
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_284
timestamp 1751532504
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_285
timestamp 1751532504
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_286
timestamp 1751532504
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_287
timestamp 1751532504
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_288
timestamp 1751532504
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_289
timestamp 1751532504
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_290
timestamp 1751532504
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_291
timestamp 1751532504
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_292
timestamp 1751532504
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_293
timestamp 1751532504
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_294
timestamp 1751532504
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_37_295
timestamp 1751532504
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_296
timestamp 1751532504
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_297
timestamp 1751532504
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_298
timestamp 1751532504
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_299
timestamp 1751532504
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_38_300
timestamp 1751532504
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_301
timestamp 1751532504
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_302
timestamp 1751532504
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_303
timestamp 1751532504
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_304
timestamp 1751532504
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_39_305
timestamp 1751532504
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_306
timestamp 1751532504
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_307
timestamp 1751532504
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_308
timestamp 1751532504
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_309
timestamp 1751532504
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_40_310
timestamp 1751532504
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_311
timestamp 1751532504
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_312
timestamp 1751532504
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_313
timestamp 1751532504
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_314
timestamp 1751532504
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_41_315
timestamp 1751532504
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_316
timestamp 1751532504
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_317
timestamp 1751532504
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_318
timestamp 1751532504
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_319
timestamp 1751532504
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_42_320
timestamp 1751532504
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_321
timestamp 1751532504
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_322
timestamp 1751532504
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_323
timestamp 1751532504
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_324
timestamp 1751532504
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_43_325
timestamp 1751532504
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_326
timestamp 1751532504
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_327
timestamp 1751532504
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_328
timestamp 1751532504
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_329
timestamp 1751532504
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_44_330
timestamp 1751532504
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_331
timestamp 1751532504
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_332
timestamp 1751532504
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_333
timestamp 1751532504
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_334
timestamp 1751532504
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_45_335
timestamp 1751532504
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_336
timestamp 1751532504
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_337
timestamp 1751532504
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_338
timestamp 1751532504
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_339
timestamp 1751532504
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_46_340
timestamp 1751532504
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_341
timestamp 1751532504
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_342
timestamp 1751532504
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_343
timestamp 1751532504
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_344
timestamp 1751532504
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_47_345
timestamp 1751532504
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_346
timestamp 1751532504
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_347
timestamp 1751532504
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_348
timestamp 1751532504
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_349
timestamp 1751532504
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_48_350
timestamp 1751532504
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_351
timestamp 1751532504
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_352
timestamp 1751532504
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_353
timestamp 1751532504
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_354
timestamp 1751532504
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_355
timestamp 1751532504
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_356
timestamp 1751532504
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_357
timestamp 1751532504
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_358
timestamp 1751532504
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_359
timestamp 1751532504
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_360
timestamp 1751532504
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_49_361
timestamp 1751532504
transform 1 0 43232 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal2 s 9408 45200 9520 46000 0 FreeSans 448 90 0 0 io_in
port 0 nsew signal input
flabel metal2 s 13216 45200 13328 46000 0 FreeSans 448 90 0 0 io_out[0]
port 1 nsew signal output
flabel metal2 s 17024 45200 17136 46000 0 FreeSans 448 90 0 0 io_out[1]
port 2 nsew signal output
flabel metal2 s 20832 45200 20944 46000 0 FreeSans 448 90 0 0 io_out[2]
port 3 nsew signal output
flabel metal2 s 24640 45200 24752 46000 0 FreeSans 448 90 0 0 io_out[3]
port 4 nsew signal output
flabel metal2 s 28448 45200 28560 46000 0 FreeSans 448 90 0 0 io_out[4]
port 5 nsew signal output
flabel metal2 s 32256 45200 32368 46000 0 FreeSans 448 90 0 0 io_out[5]
port 6 nsew signal output
flabel metal2 s 36064 45200 36176 46000 0 FreeSans 448 90 0 0 io_out[6]
port 7 nsew signal output
flabel metal2 s 39872 45200 39984 46000 0 FreeSans 448 90 0 0 io_out[7]
port 8 nsew signal output
flabel metal2 s 43680 45200 43792 46000 0 FreeSans 448 90 0 0 io_out[8]
port 9 nsew signal output
flabel metal2 s 5600 45200 5712 46000 0 FreeSans 448 90 0 0 rst_n
port 10 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal2 s 1792 45200 1904 46000 0 FreeSans 448 90 0 0 wb_clk_i
port 13 nsew signal input
rlabel metal1 22960 41552 22960 41552 0 vdd
rlabel metal1 22960 42336 22960 42336 0 vss
rlabel metal2 13944 40040 13944 40040 0 _000_
rlabel metal3 23576 39816 23576 39816 0 _001_
rlabel metal2 26768 40264 26768 40264 0 _002_
rlabel metal2 30296 40040 30296 40040 0 _003_
rlabel metal3 33488 39816 33488 39816 0 _004_
rlabel metal2 19208 40040 19208 40040 0 _005_
rlabel metal2 23688 39732 23688 39732 0 _006_
rlabel metal2 18536 13328 18536 13328 0 _007_
rlabel metal2 18200 11760 18200 11760 0 _008_
rlabel metal2 18088 7728 18088 7728 0 _009_
rlabel metal3 19208 4200 19208 4200 0 _010_
rlabel metal2 24248 4592 24248 4592 0 _011_
rlabel metal2 25592 9492 25592 9492 0 _012_
rlabel metal2 27720 4592 27720 4592 0 _013_
rlabel metal2 34104 5432 34104 5432 0 _014_
rlabel metal3 34776 9240 34776 9240 0 _015_
rlabel metal2 28280 10864 28280 10864 0 _016_
rlabel metal2 26532 37200 26532 37200 0 _017_
rlabel metal2 29624 33684 29624 33684 0 _018_
rlabel metal2 24584 35784 24584 35784 0 _019_
rlabel metal2 35336 18536 35336 18536 0 _020_
rlabel metal2 33320 28952 33320 28952 0 _021_
rlabel metal2 36792 21728 36792 21728 0 _022_
rlabel metal2 41048 40040 41048 40040 0 _023_
rlabel metal2 41944 14840 41944 14840 0 _024_
rlabel metal2 34664 13384 34664 13384 0 _025_
rlabel metal2 37688 10864 37688 10864 0 _026_
rlabel metal2 41832 11704 41832 11704 0 _027_
rlabel metal2 41720 17976 41720 17976 0 _028_
rlabel metal2 41496 21616 41496 21616 0 _029_
rlabel metal2 41888 26264 41888 26264 0 _030_
rlabel metal2 41944 31304 41944 31304 0 _031_
rlabel metal2 41216 34888 41216 34888 0 _032_
rlabel metal2 40152 37296 40152 37296 0 _033_
rlabel metal3 35448 34216 35448 34216 0 _034_
rlabel metal3 35224 31080 35224 31080 0 _035_
rlabel metal2 8792 17976 8792 17976 0 _036_
rlabel metal2 2632 19544 2632 19544 0 _037_
rlabel metal2 3192 24192 3192 24192 0 _038_
rlabel metal2 2632 29008 2632 29008 0 _039_
rlabel metal3 7000 35896 7000 35896 0 _040_
rlabel metal2 2632 33712 2632 33712 0 _041_
rlabel metal3 5824 40264 5824 40264 0 _042_
rlabel metal2 2912 38920 2912 38920 0 _043_
rlabel metal2 14840 15568 14840 15568 0 _044_
rlabel metal2 11256 13328 11256 13328 0 _045_
rlabel metal2 5320 14896 5320 14896 0 _046_
rlabel metal3 3416 11592 3416 11592 0 _047_
rlabel metal3 3640 9240 3640 9240 0 _048_
rlabel metal2 10920 6636 10920 6636 0 _049_
rlabel metal2 13832 5432 13832 5432 0 _050_
rlabel metal2 7560 4816 7560 4816 0 _051_
rlabel metal2 23800 21112 23800 21112 0 _052_
rlabel metal2 23576 27440 23576 27440 0 _053_
rlabel metal3 20608 18200 20608 18200 0 _054_
rlabel metal2 8792 23072 8792 23072 0 _055_
rlabel metal2 12152 31080 12152 31080 0 _056_
rlabel metal2 20552 37072 20552 37072 0 _057_
rlabel metal2 11760 35896 11760 35896 0 _058_
rlabel metal3 14168 39032 14168 39032 0 _059_
rlabel metal2 25928 19656 25928 19656 0 _060_
rlabel metal2 25928 14896 25928 14896 0 _061_
rlabel metal2 32032 14616 32032 14616 0 _062_
rlabel metal2 37184 39816 37184 39816 0 _063_
rlabel metal2 23156 16072 23156 16072 0 _064_
rlabel metal2 26488 31276 26488 31276 0 _065_
rlabel metal2 10696 25760 10696 25760 0 _066_
rlabel metal2 10360 26740 10360 26740 0 _067_
rlabel metal3 11200 29400 11200 29400 0 _068_
rlabel metal2 10304 28532 10304 28532 0 _069_
rlabel metal2 9856 28616 9856 28616 0 _070_
rlabel metal2 10024 28280 10024 28280 0 _071_
rlabel metal2 6328 28000 6328 28000 0 _072_
rlabel metal2 8120 28728 8120 28728 0 _073_
rlabel metal2 8232 28532 8232 28532 0 _074_
rlabel metal2 5768 24052 5768 24052 0 _075_
rlabel metal2 9352 26852 9352 26852 0 _076_
rlabel metal2 10808 30268 10808 30268 0 _077_
rlabel metal2 11032 31192 11032 31192 0 _078_
rlabel metal2 10864 27832 10864 27832 0 _079_
rlabel metal2 13608 22456 13608 22456 0 _080_
rlabel metal3 10696 20776 10696 20776 0 _081_
rlabel metal3 11480 20440 11480 20440 0 _082_
rlabel metal2 12040 20860 12040 20860 0 _083_
rlabel metal2 12992 11032 12992 11032 0 _084_
rlabel metal2 12152 7224 12152 7224 0 _085_
rlabel metal2 9464 12600 9464 12600 0 _086_
rlabel metal3 14224 12152 14224 12152 0 _087_
rlabel metal2 13692 20664 13692 20664 0 _088_
rlabel metal2 13944 21616 13944 21616 0 _089_
rlabel metal2 31248 6776 31248 6776 0 _090_
rlabel metal2 31864 13888 31864 13888 0 _091_
rlabel metal2 21336 13216 21336 13216 0 _092_
rlabel metal3 22148 10696 22148 10696 0 _093_
rlabel metal2 22148 7560 22148 7560 0 _094_
rlabel metal2 21840 16856 21840 16856 0 _095_
rlabel metal2 20328 20860 20328 20860 0 _096_
rlabel metal3 16352 22344 16352 22344 0 _097_
rlabel metal2 13720 28224 13720 28224 0 _098_
rlabel metal2 13832 25312 13832 25312 0 _099_
rlabel metal2 14056 27005 14056 27005 0 _100_
rlabel metal2 13440 35672 13440 35672 0 _101_
rlabel metal2 14392 29876 14392 29876 0 _102_
rlabel metal2 14728 27496 14728 27496 0 _103_
rlabel metal3 16688 27720 16688 27720 0 _104_
rlabel metal2 20216 21952 20216 21952 0 _105_
rlabel metal2 20384 28616 20384 28616 0 _106_
rlabel metal2 27552 29176 27552 29176 0 _107_
rlabel metal2 29288 17640 29288 17640 0 _108_
rlabel metal2 31060 18788 31060 18788 0 _109_
rlabel metal2 27384 22288 27384 22288 0 _110_
rlabel metal2 29064 21295 29064 21295 0 _111_
rlabel metal2 28672 27048 28672 27048 0 _112_
rlabel metal2 29456 22344 29456 22344 0 _113_
rlabel metal2 31976 22848 31976 22848 0 _114_
rlabel metal2 29960 26964 29960 26964 0 _115_
rlabel metal2 28168 29120 28168 29120 0 _116_
rlabel metal2 35056 22260 35056 22260 0 _117_
rlabel metal3 31098 22344 31098 22344 0 _118_
rlabel metal2 28616 26165 28616 26165 0 _119_
rlabel metal2 29736 24752 29736 24752 0 _120_
rlabel metal2 35560 25928 35560 25928 0 _121_
rlabel metal2 28952 25984 28952 25984 0 _122_
rlabel metal2 26264 27384 26264 27384 0 _123_
rlabel metal2 27160 30282 27160 30282 0 _124_
rlabel metal3 25424 33320 25424 33320 0 _125_
rlabel metal2 24108 33320 24108 33320 0 _126_
rlabel metal2 25200 25844 25200 25844 0 _127_
rlabel metal2 25032 26600 25032 26600 0 _128_
rlabel metal2 30388 26208 30388 26208 0 _129_
rlabel metal2 29848 27552 29848 27552 0 _130_
rlabel metal2 29064 27748 29064 27748 0 _131_
rlabel metal2 25704 29820 25704 29820 0 _132_
rlabel metal2 27832 34776 27832 34776 0 _133_
rlabel metal3 28560 38024 28560 38024 0 _134_
rlabel metal2 29512 28280 29512 28280 0 _135_
rlabel metal2 29624 28392 29624 28392 0 _136_
rlabel metal2 29876 28840 29876 28840 0 _137_
rlabel metal2 30016 33964 30016 33964 0 _138_
rlabel metal2 30184 34832 30184 34832 0 _139_
rlabel metal2 29904 38024 29904 38024 0 _140_
rlabel metal2 24024 37968 24024 37968 0 _141_
rlabel metal3 21476 17080 21476 17080 0 _142_
rlabel metal2 25312 35112 25312 35112 0 _143_
rlabel metal2 23858 37912 23858 37912 0 _144_
rlabel metal2 23464 38920 23464 38920 0 _145_
rlabel metal3 21756 30072 21756 30072 0 _146_
rlabel metal3 23464 29960 23464 29960 0 _147_
rlabel metal2 27440 30296 27440 30296 0 _148_
rlabel metal2 27888 34104 27888 34104 0 _149_
rlabel metal3 23968 38808 23968 38808 0 _150_
rlabel metal2 23856 38696 23856 38696 0 _151_
rlabel metal2 28840 39144 28840 39144 0 _152_
rlabel metal2 29764 39592 29764 39592 0 _153_
rlabel metal2 29400 36456 29400 36456 0 _154_
rlabel metal2 20552 39536 20552 39536 0 _155_
rlabel metal3 34328 26264 34328 26264 0 _156_
rlabel metal2 25312 24248 25312 24248 0 _157_
rlabel metal2 27244 6104 27244 6104 0 _158_
rlabel metal2 20216 11424 20216 11424 0 _159_
rlabel metal2 28616 13048 28616 13048 0 _160_
rlabel metal2 23912 15904 23912 15904 0 _161_
rlabel metal2 19880 11584 19880 11584 0 _162_
rlabel metal2 20104 8548 20104 8548 0 _163_
rlabel metal2 20580 7560 20580 7560 0 _164_
rlabel metal2 18424 7728 18424 7728 0 _165_
rlabel metal3 21028 5656 21028 5656 0 _166_
rlabel metal3 20244 5880 20244 5880 0 _167_
rlabel metal2 20104 5292 20104 5292 0 _168_
rlabel metal3 23212 5880 23212 5880 0 _169_
rlabel via2 27048 9792 27048 9792 0 _170_
rlabel metal2 23800 7000 23800 7000 0 _171_
rlabel metal2 23912 4984 23912 4984 0 _172_
rlabel metal3 25340 10584 25340 10584 0 _173_
rlabel metal2 27608 6126 27608 6126 0 _174_
rlabel metal2 25368 25424 25368 25424 0 _175_
rlabel metal2 25424 9100 25424 9100 0 _176_
rlabel metal3 28056 5768 28056 5768 0 _177_
rlabel metal2 31584 5025 31584 5025 0 _178_
rlabel metal2 28504 5572 28504 5572 0 _179_
rlabel metal2 31528 5563 31528 5563 0 _180_
rlabel metal2 31864 6552 31864 6552 0 _181_
rlabel metal2 31864 5964 31864 5964 0 _182_
rlabel metal2 32312 9240 32312 9240 0 _183_
rlabel metal2 33152 9464 33152 9464 0 _184_
rlabel metal2 32592 10080 32592 10080 0 _185_
rlabel metal2 33768 9464 33768 9464 0 _186_
rlabel metal2 27832 10080 27832 10080 0 _187_
rlabel metal2 28084 10024 28084 10024 0 _188_
rlabel metal2 36960 26264 36960 26264 0 _189_
rlabel metal3 36932 23016 36932 23016 0 _190_
rlabel metal3 37016 23912 37016 23912 0 _191_
rlabel metal3 38640 23688 38640 23688 0 _192_
rlabel metal2 35616 20888 35616 20888 0 _193_
rlabel metal2 39032 18368 39032 18368 0 _194_
rlabel metal3 37352 20216 37352 20216 0 _195_
rlabel metal2 38304 17864 38304 17864 0 _196_
rlabel metal3 37632 20328 37632 20328 0 _197_
rlabel metal2 35840 19516 35840 19516 0 _198_
rlabel metal2 36456 30590 36456 30590 0 _199_
rlabel metal2 36624 26488 36624 26488 0 _200_
rlabel metal2 37128 28336 37128 28336 0 _201_
rlabel metal3 35477 28616 35477 28616 0 _202_
rlabel metal2 33656 29288 33656 29288 0 _203_
rlabel metal2 39648 22652 39648 22652 0 _204_
rlabel metal2 22736 31528 22736 31528 0 _205_
rlabel metal2 39816 22736 39816 22736 0 _206_
rlabel metal3 37744 22344 37744 22344 0 _207_
rlabel metal2 39032 24472 39032 24472 0 _208_
rlabel metal2 39844 27272 39844 27272 0 _209_
rlabel metal2 40544 30632 40544 30632 0 _210_
rlabel metal2 39704 15568 39704 15568 0 _211_
rlabel via2 39850 15306 39850 15306 0 _212_
rlabel metal2 40488 14784 40488 14784 0 _213_
rlabel metal3 25340 18312 25340 18312 0 _214_
rlabel via1 34440 14490 34440 14490 0 _215_
rlabel metal2 15792 18228 15792 18228 0 _216_
rlabel metal2 20776 27832 20776 27832 0 _217_
rlabel metal2 34776 14840 34776 14840 0 _218_
rlabel metal2 34328 13636 34328 13636 0 _219_
rlabel metal2 39182 12227 39182 12227 0 _220_
rlabel metal2 38920 11648 38920 11648 0 _221_
rlabel metal2 40179 12936 40179 12936 0 _222_
rlabel metal3 40880 12152 40880 12152 0 _223_
rlabel metal2 41188 18648 41188 18648 0 _224_
rlabel metal2 41272 21056 41272 21056 0 _225_
rlabel metal2 40292 21336 40292 21336 0 _226_
rlabel metal3 41972 25256 41972 25256 0 _227_
rlabel metal2 41664 21084 41664 21084 0 _228_
rlabel metal2 41608 34930 41608 34930 0 _229_
rlabel metal2 35560 27160 35560 27160 0 _230_
rlabel metal2 37912 27496 37912 27496 0 _231_
rlabel metal2 41384 28168 41384 28168 0 _232_
rlabel metal2 42000 27356 42000 27356 0 _233_
rlabel metal2 42000 30576 42000 30576 0 _234_
rlabel metal2 41384 34048 41384 34048 0 _235_
rlabel metal3 37408 32536 37408 32536 0 _236_
rlabel metal2 42112 31836 42112 31836 0 _237_
rlabel metal2 40208 34888 40208 34888 0 _238_
rlabel metal3 40712 34888 40712 34888 0 _239_
rlabel metal2 40824 36764 40824 36764 0 _240_
rlabel metal2 38248 35168 38248 35168 0 _241_
rlabel metal2 39200 35168 39200 35168 0 _242_
rlabel metal2 36288 34608 36288 34608 0 _243_
rlabel metal3 36652 31528 36652 31528 0 _244_
rlabel metal2 36372 32648 36372 32648 0 _245_
rlabel metal2 35980 27272 35980 27272 0 _246_
rlabel metal2 13720 22484 13720 22484 0 _247_
rlabel metal2 6272 23128 6272 23128 0 _248_
rlabel metal3 10584 20552 10584 20552 0 _249_
rlabel metal2 21056 18536 21056 18536 0 _250_
rlabel metal2 15652 21336 15652 21336 0 _251_
rlabel metal2 7000 19096 7000 19096 0 _252_
rlabel metal3 6244 19208 6244 19208 0 _253_
rlabel metal2 10024 18732 10024 18732 0 _254_
rlabel metal2 6440 23464 6440 23464 0 _255_
rlabel metal2 16408 22400 16408 22400 0 _256_
rlabel metal2 18424 25312 18424 25312 0 _257_
rlabel metal3 5236 24024 5236 24024 0 _258_
rlabel metal3 5152 20888 5152 20888 0 _259_
rlabel metal2 6216 19488 6216 19488 0 _260_
rlabel metal2 4816 22260 4816 22260 0 _261_
rlabel metal2 3528 20076 3528 20076 0 _262_
rlabel metal2 4312 25508 4312 25508 0 _263_
rlabel metal2 3976 22792 3976 22792 0 _264_
rlabel metal2 3528 23744 3528 23744 0 _265_
rlabel metal2 14952 23128 14952 23128 0 _266_
rlabel metal3 5516 28056 5516 28056 0 _267_
rlabel metal2 4088 27888 4088 27888 0 _268_
rlabel metal2 4088 28952 4088 28952 0 _269_
rlabel metal2 5992 27070 5992 27070 0 _270_
rlabel via2 3752 29407 3752 29407 0 _271_
rlabel metal2 6552 32816 6552 32816 0 _272_
rlabel metal2 6104 34412 6104 34412 0 _273_
rlabel metal2 6048 33600 6048 33600 0 _274_
rlabel metal2 6328 35196 6328 35196 0 _275_
rlabel metal2 3696 34104 3696 34104 0 _276_
rlabel metal2 6496 33320 6496 33320 0 _277_
rlabel metal2 3304 33999 3304 33999 0 _278_
rlabel metal2 4648 37744 4648 37744 0 _279_
rlabel metal2 3080 39200 3080 39200 0 _280_
rlabel metal2 4984 39122 4984 39122 0 _281_
rlabel metal2 3304 38710 3304 38710 0 _282_
rlabel metal3 3612 38808 3612 38808 0 _283_
rlabel metal2 6300 29512 6300 29512 0 _284_
rlabel metal3 6776 29400 6776 29400 0 _285_
rlabel metal2 7476 29176 7476 29176 0 _286_
rlabel metal2 14504 17304 14504 17304 0 _287_
rlabel metal3 14980 18424 14980 18424 0 _288_
rlabel metal2 14672 16856 14672 16856 0 _289_
rlabel metal2 14952 16352 14952 16352 0 _290_
rlabel metal2 13608 14112 13608 14112 0 _291_
rlabel metal2 7672 13034 7672 13034 0 _292_
rlabel metal2 20356 16632 20356 16632 0 _293_
rlabel metal2 11368 13208 11368 13208 0 _294_
rlabel metal2 6720 11368 6720 11368 0 _295_
rlabel via2 5992 14496 5992 14496 0 _296_
rlabel metal2 7224 12076 7224 12076 0 _297_
rlabel metal2 8680 13076 8680 13076 0 _298_
rlabel metal2 12600 10584 12600 10584 0 _299_
rlabel metal2 7448 10696 7448 10696 0 _300_
rlabel metal3 5488 11368 5488 11368 0 _301_
rlabel metal3 7840 9800 7840 9800 0 _302_
rlabel metal2 7784 9912 7784 9912 0 _303_
rlabel metal2 7896 9352 7896 9352 0 _304_
rlabel metal3 5936 9016 5936 9016 0 _305_
rlabel metal2 12600 6664 12600 6664 0 _306_
rlabel metal3 10192 8232 10192 8232 0 _307_
rlabel metal2 11032 8308 11032 8308 0 _308_
rlabel metal2 7672 7093 7672 7093 0 _309_
rlabel metal3 13664 8232 13664 8232 0 _310_
rlabel metal2 14336 7448 14336 7448 0 _311_
rlabel metal2 14168 6272 14168 6272 0 _312_
rlabel metal2 7784 6272 7784 6272 0 _313_
rlabel metal2 8316 5880 8316 5880 0 _314_
rlabel metal2 8232 6384 8232 6384 0 _315_
rlabel metal2 8232 4592 8232 4592 0 _316_
rlabel metal2 20216 25088 20216 25088 0 _317_
rlabel metal2 23800 24192 23800 24192 0 _318_
rlabel metal2 23016 27141 23016 27141 0 _319_
rlabel metal2 23800 22792 23800 22792 0 _320_
rlabel metal2 24024 22680 24024 22680 0 _321_
rlabel metal2 23800 21728 23800 21728 0 _322_
rlabel metal2 20328 25032 20328 25032 0 _323_
rlabel metal2 22736 26544 22736 26544 0 _324_
rlabel metal2 24920 25536 24920 25536 0 _325_
rlabel metal2 24332 25368 24332 25368 0 _326_
rlabel metal2 18228 26376 18228 26376 0 _327_
rlabel metal2 15176 25872 15176 25872 0 _328_
rlabel metal2 19544 25424 19544 25424 0 _329_
rlabel metal2 18732 25704 18732 25704 0 _330_
rlabel metal3 19292 26040 19292 26040 0 _331_
rlabel metal2 20524 18424 20524 18424 0 _332_
rlabel metal2 14280 24892 14280 24892 0 _333_
rlabel metal3 13832 28952 13832 28952 0 _334_
rlabel metal3 11956 23912 11956 23912 0 _335_
rlabel via1 15568 29414 15568 29414 0 _336_
rlabel metal2 16660 31864 16660 31864 0 _337_
rlabel metal3 18200 31528 18200 31528 0 _338_
rlabel metal2 17136 30268 17136 30268 0 _339_
rlabel metal2 15400 30100 15400 30100 0 _340_
rlabel metal2 15736 29736 15736 29736 0 _341_
rlabel metal2 12488 30128 12488 30128 0 _342_
rlabel metal2 18424 34608 18424 34608 0 _343_
rlabel metal2 18900 34216 18900 34216 0 _344_
rlabel metal2 18984 34720 18984 34720 0 _345_
rlabel metal2 18536 34216 18536 34216 0 _346_
rlabel metal2 19236 35112 19236 35112 0 _347_
rlabel metal3 15008 34888 15008 34888 0 _348_
rlabel metal2 14336 34188 14336 34188 0 _349_
rlabel metal3 12964 34216 12964 34216 0 _350_
rlabel metal3 17332 34104 17332 34104 0 _351_
rlabel metal2 17024 35000 17024 35000 0 _352_
rlabel metal2 17500 34216 17500 34216 0 _353_
rlabel metal3 17248 37128 17248 37128 0 _354_
rlabel metal2 26936 18508 26936 18508 0 _355_
rlabel metal3 28308 18312 28308 18312 0 _356_
rlabel metal2 26264 19040 26264 19040 0 _357_
rlabel metal2 28896 16800 28896 16800 0 _358_
rlabel metal2 28392 15624 28392 15624 0 _359_
rlabel metal2 27160 14202 27160 14202 0 _360_
rlabel metal2 31640 15232 31640 15232 0 _361_
rlabel via2 31976 15295 31976 15295 0 _362_
rlabel metal2 35840 24304 35840 24304 0 _363_
rlabel metal2 19544 29064 19544 29064 0 _364_
rlabel metal3 29008 29176 29008 29176 0 _365_
rlabel metal2 36792 39144 36792 39144 0 _366_
rlabel metal2 30856 35252 30856 35252 0 bcd\[0\]
rlabel metal3 30576 33320 30576 33320 0 bcd\[1\]
rlabel metal3 25200 31752 25200 31752 0 bcd\[2\]
rlabel metal2 23044 24696 23044 24696 0 clkdiv\[0\]
rlabel metal2 22008 27832 22008 27832 0 clkdiv\[1\]
rlabel via2 13944 26271 13944 26271 0 clkdiv\[2\]
rlabel metal2 10696 23184 10696 23184 0 clkdiv\[3\]
rlabel metal2 12264 30184 12264 30184 0 clkdiv\[4\]
rlabel metal2 7784 31360 7784 31360 0 clkdiv\[5\]
rlabel metal2 10808 36008 10808 36008 0 clkdiv\[6\]
rlabel metal2 10360 39144 10360 39144 0 clkdiv\[7\]
rlabel metal2 22456 26544 22456 26544 0 clknet_0_wb_clk_i
rlabel metal3 6216 5096 6216 5096 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 17612 15512 17612 15512 0 clknet_3_1__leaf_wb_clk_i
rlabel metal3 6636 24584 6636 24584 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 14952 31261 14952 31261 0 clknet_3_3__leaf_wb_clk_i
rlabel metal3 28588 4312 28588 4312 0 clknet_3_4__leaf_wb_clk_i
rlabel metal3 35756 5208 35756 5208 0 clknet_3_5__leaf_wb_clk_i
rlabel metal3 23632 31864 23632 31864 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 40796 26264 40796 26264 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 10696 18480 10696 18480 0 counter\[0\]
rlabel metal2 7896 13720 7896 13720 0 counter\[10\]
rlabel metal2 7056 12796 7056 12796 0 counter\[11\]
rlabel metal2 7112 9856 7112 9856 0 counter\[12\]
rlabel metal2 12768 5880 12768 5880 0 counter\[13\]
rlabel via2 12488 5899 12488 5899 0 counter\[14\]
rlabel metal3 10920 5880 10920 5880 0 counter\[15\]
rlabel metal2 6048 23128 6048 23128 0 counter\[1\]
rlabel metal3 5880 24696 5880 24696 0 counter\[2\]
rlabel metal2 5432 22456 5432 22456 0 counter\[3\]
rlabel metal3 9744 30968 9744 30968 0 counter\[4\]
rlabel metal2 6907 31836 6907 31836 0 counter\[5\]
rlabel metal2 9912 37520 9912 37520 0 counter\[6\]
rlabel metal2 4716 37203 4716 37203 0 counter\[7\]
rlabel metal3 15904 15176 15904 15176 0 counter\[8\]
rlabel metal3 13944 13720 13944 13720 0 counter\[9\]
rlabel metal3 37576 40488 37576 40488 0 dp
rlabel metal2 9464 44478 9464 44478 0 io_in
rlabel metal3 13888 41832 13888 41832 0 io_out[0]
rlabel metal3 17696 41832 17696 41832 0 io_out[1]
rlabel metal3 21504 41832 21504 41832 0 io_out[2]
rlabel metal3 25312 41832 25312 41832 0 io_out[3]
rlabel metal3 29120 41832 29120 41832 0 io_out[4]
rlabel metal3 32928 41832 32928 41832 0 io_out[5]
rlabel metal3 36736 41832 36736 41832 0 io_out[6]
rlabel metal3 40544 41832 40544 41832 0 io_out[7]
rlabel metal2 43736 43218 43736 43218 0 io_out[8]
rlabel metal3 33992 21560 33992 21560 0 lfsr\[0\]
rlabel metal2 43848 25816 43848 25816 0 lfsr\[10\]
rlabel metal2 42168 30520 42168 30520 0 lfsr\[11\]
rlabel metal2 42840 35112 42840 35112 0 lfsr\[12\]
rlabel metal2 41160 36792 41160 36792 0 lfsr\[13\]
rlabel metal3 37342 35672 37342 35672 0 lfsr\[14\]
rlabel metal3 36624 31752 36624 31752 0 lfsr\[15\]
rlabel metal2 28840 21644 28840 21644 0 lfsr\[1\]
rlabel metal2 34888 22624 34888 22624 0 lfsr\[2\]
rlabel metal2 40236 23912 40236 23912 0 lfsr\[3\]
rlabel metal2 43848 15064 43848 15064 0 lfsr\[4\]
rlabel metal3 36596 15288 36596 15288 0 lfsr\[5\]
rlabel metal2 39536 12152 39536 12152 0 lfsr\[6\]
rlabel metal2 43736 12208 43736 12208 0 lfsr\[7\]
rlabel metal3 40208 18424 40208 18424 0 lfsr\[8\]
rlabel metal2 42840 21896 42840 21896 0 lfsr\[9\]
rlabel metal3 20944 13720 20944 13720 0 m_clkdiv\[0\]
rlabel metal2 20328 13608 20328 13608 0 m_clkdiv\[1\]
rlabel metal2 21784 8436 21784 8436 0 m_clkdiv\[2\]
rlabel metal2 20888 5544 20888 5544 0 m_clkdiv\[3\]
rlabel metal2 22456 5544 22456 5544 0 m_clkdiv\[4\]
rlabel metal2 23800 10248 23800 10248 0 m_clkdiv\[5\]
rlabel metal2 29512 5936 29512 5936 0 m_clkdiv\[6\]
rlabel metal2 31472 6664 31472 6664 0 m_clkdiv\[7\]
rlabel metal2 31416 9380 31416 9380 0 m_clkdiv\[8\]
rlabel metal2 30184 10304 30184 10304 0 m_clkdiv\[9\]
rlabel metal3 12068 24024 12068 24024 0 net1
rlabel metal3 39928 40600 39928 40600 0 net10
rlabel metal3 42224 39816 42224 39816 0 net11
rlabel metal2 6216 37856 6216 37856 0 net2
rlabel metal2 11816 40544 11816 40544 0 net3
rlabel metal2 15848 40096 15848 40096 0 net4
rlabel metal2 21112 41229 21112 41229 0 net5
rlabel metal2 24584 40824 24584 40824 0 net6
rlabel metal2 28728 41229 28728 41229 0 net7
rlabel metal2 32480 40488 32480 40488 0 net8
rlabel metal2 36008 40824 36008 40824 0 net9
rlabel metal2 29064 20468 29064 20468 0 r_counter\[0\]
rlabel metal2 29316 21000 29316 21000 0 r_counter\[1\]
rlabel metal2 30968 15960 30968 15960 0 r_counter\[2\]
rlabel metal2 5656 44478 5656 44478 0 rst_n
rlabel metal2 21672 23197 21672 23197 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
