magic
tech gf180mcuD
magscale 1 10
timestamp 1702311871
<< metal1 >>
rect 1344 20410 22784 20444
rect 1344 20358 6534 20410
rect 6586 20358 6638 20410
rect 6690 20358 6742 20410
rect 6794 20358 11854 20410
rect 11906 20358 11958 20410
rect 12010 20358 12062 20410
rect 12114 20358 17174 20410
rect 17226 20358 17278 20410
rect 17330 20358 17382 20410
rect 17434 20358 22494 20410
rect 22546 20358 22598 20410
rect 22650 20358 22702 20410
rect 22754 20358 22784 20410
rect 1344 20324 22784 20358
rect 2034 20078 2046 20130
rect 2098 20078 2110 20130
rect 4274 20078 4286 20130
rect 4338 20078 4350 20130
rect 6514 20078 6526 20130
rect 6578 20078 6590 20130
rect 9314 20078 9326 20130
rect 9378 20078 9390 20130
rect 10994 20078 11006 20130
rect 11058 20078 11070 20130
rect 13234 20078 13246 20130
rect 13298 20078 13310 20130
rect 15474 20078 15486 20130
rect 15538 20078 15550 20130
rect 17714 20078 17726 20130
rect 17778 20078 17790 20130
rect 20178 20078 20190 20130
rect 20242 20078 20254 20130
rect 20738 20078 20750 20130
rect 20802 20078 20814 20130
rect 22194 20078 22206 20130
rect 22258 20078 22270 20130
rect 2382 20018 2434 20030
rect 13582 20018 13634 20030
rect 19854 20018 19906 20030
rect 21870 20018 21922 20030
rect 4498 19966 4510 20018
rect 4562 19966 4574 20018
rect 6738 19966 6750 20018
rect 6802 19966 6814 20018
rect 9538 19966 9550 20018
rect 9602 19966 9614 20018
rect 11218 19966 11230 20018
rect 11282 19966 11294 20018
rect 15698 19966 15710 20018
rect 15762 19966 15774 20018
rect 17938 19966 17950 20018
rect 18002 19966 18014 20018
rect 20962 19966 20974 20018
rect 21026 19966 21038 20018
rect 2382 19954 2434 19966
rect 13582 19954 13634 19966
rect 19854 19954 19906 19966
rect 21870 19954 21922 19966
rect 18846 19906 18898 19918
rect 18846 19842 18898 19854
rect 18734 19794 18786 19806
rect 18734 19730 18786 19742
rect 1344 19626 22624 19660
rect 1344 19574 3874 19626
rect 3926 19574 3978 19626
rect 4030 19574 4082 19626
rect 4134 19574 9194 19626
rect 9246 19574 9298 19626
rect 9350 19574 9402 19626
rect 9454 19574 14514 19626
rect 14566 19574 14618 19626
rect 14670 19574 14722 19626
rect 14774 19574 19834 19626
rect 19886 19574 19938 19626
rect 19990 19574 20042 19626
rect 20094 19574 22624 19626
rect 1344 19540 22624 19574
rect 4510 19458 4562 19470
rect 4510 19394 4562 19406
rect 6190 19346 6242 19358
rect 18510 19346 18562 19358
rect 5842 19294 5854 19346
rect 5906 19294 5918 19346
rect 6514 19294 6526 19346
rect 6578 19294 6590 19346
rect 7522 19294 7534 19346
rect 7586 19294 7598 19346
rect 11666 19294 11678 19346
rect 11730 19294 11742 19346
rect 13794 19294 13806 19346
rect 13858 19294 13870 19346
rect 6190 19282 6242 19294
rect 18510 19282 18562 19294
rect 3054 19234 3106 19246
rect 13470 19234 13522 19246
rect 17950 19234 18002 19246
rect 19294 19234 19346 19246
rect 3378 19182 3390 19234
rect 3442 19182 3454 19234
rect 15250 19182 15262 19234
rect 15314 19182 15326 19234
rect 18722 19182 18734 19234
rect 18786 19182 18798 19234
rect 3054 19170 3106 19182
rect 13470 19170 13522 19182
rect 17950 19170 18002 19182
rect 19294 19170 19346 19182
rect 21646 19234 21698 19246
rect 21646 19170 21698 19182
rect 4622 19122 4674 19134
rect 4622 19058 4674 19070
rect 6862 19122 6914 19134
rect 6862 19058 6914 19070
rect 7198 19122 7250 19134
rect 11454 19122 11506 19134
rect 18062 19122 18114 19134
rect 10098 19070 10110 19122
rect 10162 19070 10174 19122
rect 15474 19070 15486 19122
rect 15538 19070 15550 19122
rect 7198 19058 7250 19070
rect 11454 19058 11506 19070
rect 18062 19058 18114 19070
rect 18398 19122 18450 19134
rect 18398 19058 18450 19070
rect 19182 19122 19234 19134
rect 19182 19058 19234 19070
rect 19630 19122 19682 19134
rect 19630 19058 19682 19070
rect 3166 19010 3218 19022
rect 3166 18946 3218 18958
rect 3950 19010 4002 19022
rect 3950 18946 4002 18958
rect 5966 19010 6018 19022
rect 5966 18946 6018 18958
rect 6638 19010 6690 19022
rect 6638 18946 6690 18958
rect 7422 19010 7474 19022
rect 7422 18946 7474 18958
rect 9774 19010 9826 19022
rect 9774 18946 9826 18958
rect 11678 19010 11730 19022
rect 11678 18946 11730 18958
rect 13694 19010 13746 19022
rect 13694 18946 13746 18958
rect 19406 19010 19458 19022
rect 19406 18946 19458 18958
rect 21310 19010 21362 19022
rect 21310 18946 21362 18958
rect 1344 18842 22784 18876
rect 1344 18790 6534 18842
rect 6586 18790 6638 18842
rect 6690 18790 6742 18842
rect 6794 18790 11854 18842
rect 11906 18790 11958 18842
rect 12010 18790 12062 18842
rect 12114 18790 17174 18842
rect 17226 18790 17278 18842
rect 17330 18790 17382 18842
rect 17434 18790 22494 18842
rect 22546 18790 22598 18842
rect 22650 18790 22702 18842
rect 22754 18790 22784 18842
rect 1344 18756 22784 18790
rect 4062 18674 4114 18686
rect 4062 18610 4114 18622
rect 5966 18674 6018 18686
rect 5966 18610 6018 18622
rect 10894 18674 10946 18686
rect 10894 18610 10946 18622
rect 14030 18674 14082 18686
rect 18610 18622 18622 18674
rect 18674 18622 18686 18674
rect 14030 18610 14082 18622
rect 3838 18562 3890 18574
rect 3838 18498 3890 18510
rect 5854 18562 5906 18574
rect 5854 18498 5906 18510
rect 7086 18562 7138 18574
rect 7086 18498 7138 18510
rect 7982 18562 8034 18574
rect 7982 18498 8034 18510
rect 11790 18562 11842 18574
rect 21870 18562 21922 18574
rect 12786 18510 12798 18562
rect 12850 18510 12862 18562
rect 15586 18510 15598 18562
rect 15650 18510 15662 18562
rect 16594 18510 16606 18562
rect 16658 18510 16670 18562
rect 11790 18498 11842 18510
rect 21870 18498 21922 18510
rect 3950 18450 4002 18462
rect 3950 18386 4002 18398
rect 4510 18450 4562 18462
rect 6750 18450 6802 18462
rect 6178 18398 6190 18450
rect 6242 18398 6254 18450
rect 4510 18386 4562 18398
rect 6750 18386 6802 18398
rect 6974 18450 7026 18462
rect 6974 18386 7026 18398
rect 7534 18450 7586 18462
rect 7534 18386 7586 18398
rect 7646 18450 7698 18462
rect 7646 18386 7698 18398
rect 10334 18450 10386 18462
rect 11454 18450 11506 18462
rect 10658 18398 10670 18450
rect 10722 18398 10734 18450
rect 11218 18398 11230 18450
rect 11282 18398 11294 18450
rect 10334 18386 10386 18398
rect 11454 18386 11506 18398
rect 12462 18450 12514 18462
rect 12462 18386 12514 18398
rect 13246 18450 13298 18462
rect 14142 18450 14194 18462
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 13246 18386 13298 18398
rect 14142 18386 14194 18398
rect 14366 18450 14418 18462
rect 14366 18386 14418 18398
rect 15934 18450 15986 18462
rect 15934 18386 15986 18398
rect 16270 18450 16322 18462
rect 16270 18386 16322 18398
rect 18286 18450 18338 18462
rect 18286 18386 18338 18398
rect 21646 18450 21698 18462
rect 21646 18386 21698 18398
rect 22206 18450 22258 18462
rect 22206 18386 22258 18398
rect 2942 18338 2994 18350
rect 2942 18274 2994 18286
rect 8430 18338 8482 18350
rect 11678 18338 11730 18350
rect 10770 18286 10782 18338
rect 10834 18286 10846 18338
rect 8430 18274 8482 18286
rect 11678 18274 11730 18286
rect 3166 18226 3218 18238
rect 3166 18162 3218 18174
rect 3502 18226 3554 18238
rect 3502 18162 3554 18174
rect 6638 18226 6690 18238
rect 6638 18162 6690 18174
rect 7870 18226 7922 18238
rect 7870 18162 7922 18174
rect 13134 18226 13186 18238
rect 13134 18162 13186 18174
rect 1344 18058 22624 18092
rect 1344 18006 3874 18058
rect 3926 18006 3978 18058
rect 4030 18006 4082 18058
rect 4134 18006 9194 18058
rect 9246 18006 9298 18058
rect 9350 18006 9402 18058
rect 9454 18006 14514 18058
rect 14566 18006 14618 18058
rect 14670 18006 14722 18058
rect 14774 18006 19834 18058
rect 19886 18006 19938 18058
rect 19990 18006 20042 18058
rect 20094 18006 22624 18058
rect 1344 17972 22624 18006
rect 6862 17890 6914 17902
rect 6862 17826 6914 17838
rect 11006 17890 11058 17902
rect 19854 17890 19906 17902
rect 12002 17838 12014 17890
rect 12066 17838 12078 17890
rect 11006 17826 11058 17838
rect 19854 17826 19906 17838
rect 4510 17778 4562 17790
rect 4510 17714 4562 17726
rect 5070 17778 5122 17790
rect 5070 17714 5122 17726
rect 7086 17778 7138 17790
rect 7086 17714 7138 17726
rect 19518 17778 19570 17790
rect 19518 17714 19570 17726
rect 19966 17778 20018 17790
rect 19966 17714 20018 17726
rect 2942 17666 2994 17678
rect 2942 17602 2994 17614
rect 3166 17666 3218 17678
rect 3166 17602 3218 17614
rect 3390 17666 3442 17678
rect 3390 17602 3442 17614
rect 3502 17666 3554 17678
rect 3502 17602 3554 17614
rect 3950 17666 4002 17678
rect 20190 17666 20242 17678
rect 11218 17614 11230 17666
rect 11282 17614 11294 17666
rect 3950 17602 4002 17614
rect 20190 17602 20242 17614
rect 20302 17666 20354 17678
rect 20302 17602 20354 17614
rect 10446 17554 10498 17566
rect 10446 17490 10498 17502
rect 11454 17554 11506 17566
rect 11454 17490 11506 17502
rect 11566 17554 11618 17566
rect 11566 17490 11618 17502
rect 3614 17442 3666 17454
rect 3614 17378 3666 17390
rect 4398 17442 4450 17454
rect 4398 17378 4450 17390
rect 4622 17442 4674 17454
rect 10670 17442 10722 17454
rect 6514 17390 6526 17442
rect 6578 17390 6590 17442
rect 4622 17378 4674 17390
rect 10670 17378 10722 17390
rect 10894 17442 10946 17454
rect 10894 17378 10946 17390
rect 1344 17274 22784 17308
rect 1344 17222 6534 17274
rect 6586 17222 6638 17274
rect 6690 17222 6742 17274
rect 6794 17222 11854 17274
rect 11906 17222 11958 17274
rect 12010 17222 12062 17274
rect 12114 17222 17174 17274
rect 17226 17222 17278 17274
rect 17330 17222 17382 17274
rect 17434 17222 22494 17274
rect 22546 17222 22598 17274
rect 22650 17222 22702 17274
rect 22754 17222 22784 17274
rect 1344 17188 22784 17222
rect 3950 17106 4002 17118
rect 3950 17042 4002 17054
rect 11006 17106 11058 17118
rect 11006 17042 11058 17054
rect 11118 17106 11170 17118
rect 11118 17042 11170 17054
rect 11230 17106 11282 17118
rect 11230 17042 11282 17054
rect 20302 17106 20354 17118
rect 20302 17042 20354 17054
rect 3054 16994 3106 17006
rect 3054 16930 3106 16942
rect 9662 16994 9714 17006
rect 9662 16930 9714 16942
rect 11342 16994 11394 17006
rect 11342 16930 11394 16942
rect 15038 16994 15090 17006
rect 15038 16930 15090 16942
rect 20638 16994 20690 17006
rect 20638 16930 20690 16942
rect 21870 16994 21922 17006
rect 21870 16930 21922 16942
rect 3278 16882 3330 16894
rect 3278 16818 3330 16830
rect 3614 16882 3666 16894
rect 12238 16882 12290 16894
rect 19630 16882 19682 16894
rect 11778 16830 11790 16882
rect 11842 16830 11854 16882
rect 15586 16830 15598 16882
rect 15650 16830 15662 16882
rect 19394 16830 19406 16882
rect 19458 16830 19470 16882
rect 3614 16818 3666 16830
rect 12238 16818 12290 16830
rect 19630 16818 19682 16830
rect 19966 16882 20018 16894
rect 19966 16818 20018 16830
rect 20414 16882 20466 16894
rect 20414 16818 20466 16830
rect 20974 16882 21026 16894
rect 20974 16818 21026 16830
rect 21198 16882 21250 16894
rect 21198 16818 21250 16830
rect 21646 16882 21698 16894
rect 21646 16818 21698 16830
rect 22206 16882 22258 16894
rect 22206 16818 22258 16830
rect 15150 16770 15202 16782
rect 9538 16718 9550 16770
rect 9602 16718 9614 16770
rect 15150 16706 15202 16718
rect 21086 16770 21138 16782
rect 21086 16706 21138 16718
rect 3838 16658 3890 16670
rect 3838 16594 3890 16606
rect 9886 16658 9938 16670
rect 9886 16594 9938 16606
rect 15262 16658 15314 16670
rect 15262 16594 15314 16606
rect 15598 16658 15650 16670
rect 15598 16594 15650 16606
rect 15934 16658 15986 16670
rect 15934 16594 15986 16606
rect 19742 16658 19794 16670
rect 19742 16594 19794 16606
rect 1344 16490 22624 16524
rect 1344 16438 3874 16490
rect 3926 16438 3978 16490
rect 4030 16438 4082 16490
rect 4134 16438 9194 16490
rect 9246 16438 9298 16490
rect 9350 16438 9402 16490
rect 9454 16438 14514 16490
rect 14566 16438 14618 16490
rect 14670 16438 14722 16490
rect 14774 16438 19834 16490
rect 19886 16438 19938 16490
rect 19990 16438 20042 16490
rect 20094 16438 22624 16490
rect 1344 16404 22624 16438
rect 15038 16322 15090 16334
rect 15038 16258 15090 16270
rect 19406 16322 19458 16334
rect 19406 16258 19458 16270
rect 19742 16322 19794 16334
rect 19742 16258 19794 16270
rect 21310 16322 21362 16334
rect 21310 16258 21362 16270
rect 19630 16210 19682 16222
rect 19630 16146 19682 16158
rect 22318 16210 22370 16222
rect 22318 16146 22370 16158
rect 6190 16098 6242 16110
rect 4610 16046 4622 16098
rect 4674 16046 4686 16098
rect 6190 16034 6242 16046
rect 14926 16098 14978 16110
rect 14926 16034 14978 16046
rect 15262 16098 15314 16110
rect 20078 16098 20130 16110
rect 15474 16046 15486 16098
rect 15538 16046 15550 16098
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 15262 16034 15314 16046
rect 20078 16034 20130 16046
rect 21422 16098 21474 16110
rect 21422 16034 21474 16046
rect 4846 15986 4898 15998
rect 4846 15922 4898 15934
rect 20414 15986 20466 15998
rect 20414 15922 20466 15934
rect 20638 15986 20690 15998
rect 20638 15922 20690 15934
rect 20302 15874 20354 15886
rect 5842 15822 5854 15874
rect 5906 15822 5918 15874
rect 20302 15810 20354 15822
rect 1344 15706 22784 15740
rect 1344 15654 6534 15706
rect 6586 15654 6638 15706
rect 6690 15654 6742 15706
rect 6794 15654 11854 15706
rect 11906 15654 11958 15706
rect 12010 15654 12062 15706
rect 12114 15654 17174 15706
rect 17226 15654 17278 15706
rect 17330 15654 17382 15706
rect 17434 15654 22494 15706
rect 22546 15654 22598 15706
rect 22650 15654 22702 15706
rect 22754 15654 22784 15706
rect 1344 15620 22784 15654
rect 3390 15538 3442 15550
rect 3390 15474 3442 15486
rect 8878 15538 8930 15550
rect 8878 15474 8930 15486
rect 9662 15538 9714 15550
rect 9662 15474 9714 15486
rect 9774 15538 9826 15550
rect 19966 15538 20018 15550
rect 10434 15486 10446 15538
rect 10498 15486 10510 15538
rect 9774 15474 9826 15486
rect 19966 15474 20018 15486
rect 13918 15426 13970 15438
rect 13918 15362 13970 15374
rect 14478 15426 14530 15438
rect 14478 15362 14530 15374
rect 18174 15426 18226 15438
rect 18174 15362 18226 15374
rect 20526 15426 20578 15438
rect 20526 15362 20578 15374
rect 8654 15314 8706 15326
rect 8654 15250 8706 15262
rect 8990 15314 9042 15326
rect 8990 15250 9042 15262
rect 9550 15314 9602 15326
rect 9550 15250 9602 15262
rect 10222 15314 10274 15326
rect 10222 15250 10274 15262
rect 15822 15314 15874 15326
rect 15822 15250 15874 15262
rect 19182 15314 19234 15326
rect 19182 15250 19234 15262
rect 19518 15314 19570 15326
rect 19518 15250 19570 15262
rect 19630 15314 19682 15326
rect 20302 15314 20354 15326
rect 19730 15262 19742 15314
rect 19794 15262 19806 15314
rect 19630 15250 19682 15262
rect 20302 15250 20354 15262
rect 3502 15202 3554 15214
rect 3502 15138 3554 15150
rect 11006 15202 11058 15214
rect 11006 15138 11058 15150
rect 14814 15202 14866 15214
rect 14814 15138 14866 15150
rect 17502 15202 17554 15214
rect 17502 15138 17554 15150
rect 17614 15202 17666 15214
rect 17614 15138 17666 15150
rect 17838 15202 17890 15214
rect 17838 15138 17890 15150
rect 18062 15202 18114 15214
rect 20626 15150 20638 15202
rect 20690 15150 20702 15202
rect 18062 15138 18114 15150
rect 10782 15090 10834 15102
rect 10782 15026 10834 15038
rect 13806 15090 13858 15102
rect 13806 15026 13858 15038
rect 14142 15090 14194 15102
rect 14142 15026 14194 15038
rect 14590 15090 14642 15102
rect 14590 15026 14642 15038
rect 14926 15090 14978 15102
rect 14926 15026 14978 15038
rect 15374 15090 15426 15102
rect 15374 15026 15426 15038
rect 15486 15090 15538 15102
rect 15486 15026 15538 15038
rect 15710 15090 15762 15102
rect 15710 15026 15762 15038
rect 1344 14922 22624 14956
rect 1344 14870 3874 14922
rect 3926 14870 3978 14922
rect 4030 14870 4082 14922
rect 4134 14870 9194 14922
rect 9246 14870 9298 14922
rect 9350 14870 9402 14922
rect 9454 14870 14514 14922
rect 14566 14870 14618 14922
rect 14670 14870 14722 14922
rect 14774 14870 19834 14922
rect 19886 14870 19938 14922
rect 19990 14870 20042 14922
rect 20094 14870 22624 14922
rect 1344 14836 22624 14870
rect 9202 14590 9214 14642
rect 9266 14590 9278 14642
rect 3614 14530 3666 14542
rect 3614 14466 3666 14478
rect 3838 14530 3890 14542
rect 14702 14530 14754 14542
rect 4610 14478 4622 14530
rect 4674 14478 4686 14530
rect 9314 14478 9326 14530
rect 9378 14478 9390 14530
rect 14130 14478 14142 14530
rect 14194 14478 14206 14530
rect 3838 14466 3890 14478
rect 14702 14466 14754 14478
rect 8654 14418 8706 14430
rect 8654 14354 8706 14366
rect 8878 14306 8930 14318
rect 4162 14254 4174 14306
rect 4226 14254 4238 14306
rect 4834 14254 4846 14306
rect 4898 14254 4910 14306
rect 8878 14242 8930 14254
rect 9102 14306 9154 14318
rect 9102 14242 9154 14254
rect 10334 14306 10386 14318
rect 14354 14254 14366 14306
rect 14418 14254 14430 14306
rect 15026 14254 15038 14306
rect 15090 14254 15102 14306
rect 10334 14242 10386 14254
rect 1344 14138 22784 14172
rect 1344 14086 6534 14138
rect 6586 14086 6638 14138
rect 6690 14086 6742 14138
rect 6794 14086 11854 14138
rect 11906 14086 11958 14138
rect 12010 14086 12062 14138
rect 12114 14086 17174 14138
rect 17226 14086 17278 14138
rect 17330 14086 17382 14138
rect 17434 14086 22494 14138
rect 22546 14086 22598 14138
rect 22650 14086 22702 14138
rect 22754 14086 22784 14138
rect 1344 14052 22784 14086
rect 4174 13970 4226 13982
rect 4174 13906 4226 13918
rect 9662 13970 9714 13982
rect 9662 13906 9714 13918
rect 9886 13858 9938 13870
rect 9886 13794 9938 13806
rect 21870 13858 21922 13870
rect 21870 13794 21922 13806
rect 4062 13746 4114 13758
rect 3042 13694 3054 13746
rect 3106 13694 3118 13746
rect 3490 13694 3502 13746
rect 3554 13694 3566 13746
rect 4062 13682 4114 13694
rect 4286 13746 4338 13758
rect 4286 13682 4338 13694
rect 4510 13746 4562 13758
rect 4510 13682 4562 13694
rect 4958 13746 5010 13758
rect 4958 13682 5010 13694
rect 5294 13746 5346 13758
rect 5294 13682 5346 13694
rect 5630 13746 5682 13758
rect 5630 13682 5682 13694
rect 5854 13746 5906 13758
rect 5854 13682 5906 13694
rect 9998 13746 10050 13758
rect 9998 13682 10050 13694
rect 22206 13746 22258 13758
rect 22206 13682 22258 13694
rect 3726 13634 3778 13646
rect 3726 13570 3778 13582
rect 5406 13634 5458 13646
rect 5406 13570 5458 13582
rect 5966 13634 6018 13646
rect 5966 13570 6018 13582
rect 21646 13634 21698 13646
rect 21646 13570 21698 13582
rect 1344 13354 22624 13388
rect 1344 13302 3874 13354
rect 3926 13302 3978 13354
rect 4030 13302 4082 13354
rect 4134 13302 9194 13354
rect 9246 13302 9298 13354
rect 9350 13302 9402 13354
rect 9454 13302 14514 13354
rect 14566 13302 14618 13354
rect 14670 13302 14722 13354
rect 14774 13302 19834 13354
rect 19886 13302 19938 13354
rect 19990 13302 20042 13354
rect 20094 13302 22624 13354
rect 1344 13268 22624 13302
rect 5630 13186 5682 13198
rect 5630 13122 5682 13134
rect 8430 13186 8482 13198
rect 10222 13186 10274 13198
rect 9202 13134 9214 13186
rect 9266 13183 9278 13186
rect 9266 13137 9935 13183
rect 9266 13134 9278 13137
rect 8430 13122 8482 13134
rect 3502 13074 3554 13086
rect 9889 13074 9935 13137
rect 10222 13122 10274 13134
rect 10558 13186 10610 13198
rect 10558 13122 10610 13134
rect 14590 13186 14642 13198
rect 14590 13122 14642 13134
rect 15038 13186 15090 13198
rect 15038 13122 15090 13134
rect 15598 13186 15650 13198
rect 15598 13122 15650 13134
rect 16270 13186 16322 13198
rect 16270 13122 16322 13134
rect 18846 13186 18898 13198
rect 18846 13122 18898 13134
rect 17950 13074 18002 13086
rect 9874 13022 9886 13074
rect 9938 13022 9950 13074
rect 3502 13010 3554 13022
rect 17950 13010 18002 13022
rect 4398 12962 4450 12974
rect 4162 12910 4174 12962
rect 4226 12910 4238 12962
rect 4398 12898 4450 12910
rect 5742 12962 5794 12974
rect 5742 12898 5794 12910
rect 9102 12962 9154 12974
rect 9102 12898 9154 12910
rect 10446 12962 10498 12974
rect 10446 12898 10498 12910
rect 14814 12962 14866 12974
rect 15710 12962 15762 12974
rect 15250 12910 15262 12962
rect 15314 12910 15326 12962
rect 14814 12898 14866 12910
rect 15710 12898 15762 12910
rect 15934 12962 15986 12974
rect 15934 12898 15986 12910
rect 16158 12962 16210 12974
rect 16158 12898 16210 12910
rect 18174 12962 18226 12974
rect 18174 12898 18226 12910
rect 18398 12962 18450 12974
rect 18398 12898 18450 12910
rect 14478 12850 14530 12862
rect 20750 12850 20802 12862
rect 19058 12798 19070 12850
rect 19122 12798 19134 12850
rect 14478 12786 14530 12798
rect 20750 12786 20802 12798
rect 5854 12738 5906 12750
rect 5854 12674 5906 12686
rect 8542 12738 8594 12750
rect 8542 12674 8594 12686
rect 8766 12738 8818 12750
rect 8766 12674 8818 12686
rect 9438 12738 9490 12750
rect 9438 12674 9490 12686
rect 10558 12738 10610 12750
rect 10558 12674 10610 12686
rect 19406 12738 19458 12750
rect 19406 12674 19458 12686
rect 20638 12738 20690 12750
rect 20638 12674 20690 12686
rect 1344 12570 22784 12604
rect 1344 12518 6534 12570
rect 6586 12518 6638 12570
rect 6690 12518 6742 12570
rect 6794 12518 11854 12570
rect 11906 12518 11958 12570
rect 12010 12518 12062 12570
rect 12114 12518 17174 12570
rect 17226 12518 17278 12570
rect 17330 12518 17382 12570
rect 17434 12518 22494 12570
rect 22546 12518 22598 12570
rect 22650 12518 22702 12570
rect 22754 12518 22784 12570
rect 1344 12484 22784 12518
rect 4958 12402 5010 12414
rect 10446 12402 10498 12414
rect 4610 12350 4622 12402
rect 4674 12350 4686 12402
rect 8978 12350 8990 12402
rect 9042 12350 9054 12402
rect 4958 12338 5010 12350
rect 10446 12338 10498 12350
rect 19406 12402 19458 12414
rect 21422 12402 21474 12414
rect 20738 12350 20750 12402
rect 20802 12350 20814 12402
rect 19406 12338 19458 12350
rect 21422 12338 21474 12350
rect 21534 12402 21586 12414
rect 21534 12338 21586 12350
rect 21870 12402 21922 12414
rect 21870 12338 21922 12350
rect 19294 12290 19346 12302
rect 9986 12238 9998 12290
rect 10050 12238 10062 12290
rect 19294 12226 19346 12238
rect 21646 12290 21698 12302
rect 21646 12226 21698 12238
rect 10446 12178 10498 12190
rect 9762 12126 9774 12178
rect 9826 12126 9838 12178
rect 10446 12114 10498 12126
rect 11566 12178 11618 12190
rect 11566 12114 11618 12126
rect 18062 12178 18114 12190
rect 18062 12114 18114 12126
rect 18286 12178 18338 12190
rect 18286 12114 18338 12126
rect 19182 12178 19234 12190
rect 19182 12114 19234 12126
rect 19630 12178 19682 12190
rect 19630 12114 19682 12126
rect 20302 12178 20354 12190
rect 20750 12178 20802 12190
rect 20514 12126 20526 12178
rect 20578 12126 20590 12178
rect 21074 12126 21086 12178
rect 21138 12126 21150 12178
rect 20302 12114 20354 12126
rect 20750 12114 20802 12126
rect 8430 12066 8482 12078
rect 8430 12002 8482 12014
rect 10782 12066 10834 12078
rect 10782 12002 10834 12014
rect 11342 12066 11394 12078
rect 11342 12002 11394 12014
rect 8654 11954 8706 11966
rect 8654 11890 8706 11902
rect 10558 11954 10610 11966
rect 10558 11890 10610 11902
rect 11230 11954 11282 11966
rect 11230 11890 11282 11902
rect 11678 11954 11730 11966
rect 11678 11890 11730 11902
rect 17950 11954 18002 11966
rect 17950 11890 18002 11902
rect 18398 11954 18450 11966
rect 18398 11890 18450 11902
rect 1344 11786 22624 11820
rect 1344 11734 3874 11786
rect 3926 11734 3978 11786
rect 4030 11734 4082 11786
rect 4134 11734 9194 11786
rect 9246 11734 9298 11786
rect 9350 11734 9402 11786
rect 9454 11734 14514 11786
rect 14566 11734 14618 11786
rect 14670 11734 14722 11786
rect 14774 11734 19834 11786
rect 19886 11734 19938 11786
rect 19990 11734 20042 11786
rect 20094 11734 22624 11786
rect 1344 11700 22624 11734
rect 10110 11618 10162 11630
rect 10110 11554 10162 11566
rect 12238 11618 12290 11630
rect 12238 11554 12290 11566
rect 12574 11618 12626 11630
rect 12574 11554 12626 11566
rect 13918 11618 13970 11630
rect 13918 11554 13970 11566
rect 14702 11618 14754 11630
rect 14702 11554 14754 11566
rect 15038 11618 15090 11630
rect 15038 11554 15090 11566
rect 17054 11618 17106 11630
rect 17054 11554 17106 11566
rect 17166 11618 17218 11630
rect 17166 11554 17218 11566
rect 17390 11618 17442 11630
rect 17390 11554 17442 11566
rect 20302 11618 20354 11630
rect 20302 11554 20354 11566
rect 20638 11618 20690 11630
rect 20638 11554 20690 11566
rect 3726 11506 3778 11518
rect 3726 11442 3778 11454
rect 10334 11394 10386 11406
rect 12462 11394 12514 11406
rect 14926 11394 14978 11406
rect 10546 11342 10558 11394
rect 10610 11342 10622 11394
rect 13682 11342 13694 11394
rect 13746 11342 13758 11394
rect 14242 11342 14254 11394
rect 14306 11342 14318 11394
rect 10334 11330 10386 11342
rect 12462 11330 12514 11342
rect 14926 11330 14978 11342
rect 15822 11394 15874 11406
rect 18062 11394 18114 11406
rect 17602 11342 17614 11394
rect 17666 11342 17678 11394
rect 15822 11330 15874 11342
rect 18062 11330 18114 11342
rect 9998 11282 10050 11294
rect 9998 11218 10050 11230
rect 13470 11282 13522 11294
rect 13470 11218 13522 11230
rect 14590 11282 14642 11294
rect 16494 11282 16546 11294
rect 20414 11282 20466 11294
rect 15474 11230 15486 11282
rect 15538 11230 15550 11282
rect 16146 11230 16158 11282
rect 16210 11230 16222 11282
rect 18386 11230 18398 11282
rect 18450 11230 18462 11282
rect 14590 11218 14642 11230
rect 16494 11218 16546 11230
rect 20414 11218 20466 11230
rect 3614 11170 3666 11182
rect 3614 11106 3666 11118
rect 12574 11170 12626 11182
rect 12574 11106 12626 11118
rect 13582 11170 13634 11182
rect 13582 11106 13634 11118
rect 1344 11002 22784 11036
rect 1344 10950 6534 11002
rect 6586 10950 6638 11002
rect 6690 10950 6742 11002
rect 6794 10950 11854 11002
rect 11906 10950 11958 11002
rect 12010 10950 12062 11002
rect 12114 10950 17174 11002
rect 17226 10950 17278 11002
rect 17330 10950 17382 11002
rect 17434 10950 22494 11002
rect 22546 10950 22598 11002
rect 22650 10950 22702 11002
rect 22754 10950 22784 11002
rect 1344 10916 22784 10950
rect 3278 10834 3330 10846
rect 3278 10770 3330 10782
rect 9550 10834 9602 10846
rect 19854 10834 19906 10846
rect 14242 10782 14254 10834
rect 14306 10782 14318 10834
rect 9550 10770 9602 10782
rect 19854 10770 19906 10782
rect 21870 10722 21922 10734
rect 21870 10658 21922 10670
rect 2942 10610 2994 10622
rect 2942 10546 2994 10558
rect 3054 10610 3106 10622
rect 3054 10546 3106 10558
rect 3390 10610 3442 10622
rect 15038 10610 15090 10622
rect 14466 10558 14478 10610
rect 14530 10558 14542 10610
rect 3390 10546 3442 10558
rect 15038 10546 15090 10558
rect 15262 10610 15314 10622
rect 15262 10546 15314 10558
rect 15598 10610 15650 10622
rect 15598 10546 15650 10558
rect 19966 10610 20018 10622
rect 19966 10546 20018 10558
rect 22206 10610 22258 10622
rect 22206 10546 22258 10558
rect 3166 10498 3218 10510
rect 3166 10434 3218 10446
rect 9662 10498 9714 10510
rect 9662 10434 9714 10446
rect 15374 10498 15426 10510
rect 15374 10434 15426 10446
rect 21646 10498 21698 10510
rect 21646 10434 21698 10446
rect 1344 10218 22624 10252
rect 1344 10166 3874 10218
rect 3926 10166 3978 10218
rect 4030 10166 4082 10218
rect 4134 10166 9194 10218
rect 9246 10166 9298 10218
rect 9350 10166 9402 10218
rect 9454 10166 14514 10218
rect 14566 10166 14618 10218
rect 14670 10166 14722 10218
rect 14774 10166 19834 10218
rect 19886 10166 19938 10218
rect 19990 10166 20042 10218
rect 20094 10166 22624 10218
rect 1344 10132 22624 10166
rect 5630 10050 5682 10062
rect 3602 9998 3614 10050
rect 3666 9998 3678 10050
rect 5630 9986 5682 9998
rect 9326 10050 9378 10062
rect 9326 9986 9378 9998
rect 9438 10050 9490 10062
rect 20514 9998 20526 10050
rect 20578 9998 20590 10050
rect 9438 9986 9490 9998
rect 4958 9938 5010 9950
rect 19518 9938 19570 9950
rect 5954 9886 5966 9938
rect 6018 9886 6030 9938
rect 4958 9874 5010 9886
rect 19518 9874 19570 9886
rect 2942 9826 2994 9838
rect 2942 9762 2994 9774
rect 3838 9826 3890 9838
rect 3838 9762 3890 9774
rect 4286 9826 4338 9838
rect 4286 9762 4338 9774
rect 4510 9826 4562 9838
rect 4510 9762 4562 9774
rect 9886 9826 9938 9838
rect 9886 9762 9938 9774
rect 10110 9826 10162 9838
rect 10110 9762 10162 9774
rect 19406 9826 19458 9838
rect 19406 9762 19458 9774
rect 19966 9826 20018 9838
rect 20178 9774 20190 9826
rect 20242 9774 20254 9826
rect 20738 9774 20750 9826
rect 20802 9774 20814 9826
rect 19966 9762 20018 9774
rect 3054 9714 3106 9726
rect 3054 9650 3106 9662
rect 3166 9714 3218 9726
rect 3166 9650 3218 9662
rect 5854 9714 5906 9726
rect 5854 9650 5906 9662
rect 9550 9714 9602 9726
rect 9550 9650 9602 9662
rect 19182 9714 19234 9726
rect 19182 9650 19234 9662
rect 19630 9714 19682 9726
rect 19630 9650 19682 9662
rect 20078 9714 20130 9726
rect 20078 9650 20130 9662
rect 4398 9602 4450 9614
rect 4398 9538 4450 9550
rect 5070 9602 5122 9614
rect 5070 9538 5122 9550
rect 1344 9434 22784 9468
rect 1344 9382 6534 9434
rect 6586 9382 6638 9434
rect 6690 9382 6742 9434
rect 6794 9382 11854 9434
rect 11906 9382 11958 9434
rect 12010 9382 12062 9434
rect 12114 9382 17174 9434
rect 17226 9382 17278 9434
rect 17330 9382 17382 9434
rect 17434 9382 22494 9434
rect 22546 9382 22598 9434
rect 22650 9382 22702 9434
rect 22754 9382 22784 9434
rect 1344 9348 22784 9382
rect 10558 9266 10610 9278
rect 5954 9214 5966 9266
rect 6018 9214 6030 9266
rect 10558 9202 10610 9214
rect 10782 9266 10834 9278
rect 10782 9202 10834 9214
rect 19854 9266 19906 9278
rect 19854 9202 19906 9214
rect 3726 9154 3778 9166
rect 4734 9154 4786 9166
rect 3938 9102 3950 9154
rect 4002 9102 4014 9154
rect 3726 9090 3778 9102
rect 4734 9090 4786 9102
rect 4958 9154 5010 9166
rect 4958 9090 5010 9102
rect 19966 9154 20018 9166
rect 19966 9090 20018 9102
rect 3614 9042 3666 9054
rect 5518 9042 5570 9054
rect 4162 8990 4174 9042
rect 4226 8990 4238 9042
rect 3614 8978 3666 8990
rect 5518 8978 5570 8990
rect 5966 9042 6018 9054
rect 5966 8978 6018 8990
rect 6302 9042 6354 9054
rect 6302 8978 6354 8990
rect 6526 9042 6578 9054
rect 10434 8990 10446 9042
rect 10498 8990 10510 9042
rect 19618 8990 19630 9042
rect 19682 8990 19694 9042
rect 6526 8978 6578 8990
rect 6078 8930 6130 8942
rect 5058 8878 5070 8930
rect 5122 8878 5134 8930
rect 10658 8878 10670 8930
rect 10722 8878 10734 8930
rect 6078 8866 6130 8878
rect 4510 8818 4562 8830
rect 4510 8754 4562 8766
rect 9886 8818 9938 8830
rect 9886 8754 9938 8766
rect 10110 8818 10162 8830
rect 10110 8754 10162 8766
rect 1344 8650 22624 8684
rect 1344 8598 3874 8650
rect 3926 8598 3978 8650
rect 4030 8598 4082 8650
rect 4134 8598 9194 8650
rect 9246 8598 9298 8650
rect 9350 8598 9402 8650
rect 9454 8598 14514 8650
rect 14566 8598 14618 8650
rect 14670 8598 14722 8650
rect 14774 8598 19834 8650
rect 19886 8598 19938 8650
rect 19990 8598 20042 8650
rect 20094 8598 22624 8650
rect 1344 8564 22624 8598
rect 10782 8482 10834 8494
rect 4834 8430 4846 8482
rect 4898 8430 4910 8482
rect 20290 8430 20302 8482
rect 20354 8430 20366 8482
rect 10782 8418 10834 8430
rect 9886 8370 9938 8382
rect 10446 8370 10498 8382
rect 11342 8370 11394 8382
rect 10098 8318 10110 8370
rect 10162 8318 10174 8370
rect 11106 8318 11118 8370
rect 11170 8318 11182 8370
rect 9886 8306 9938 8318
rect 10446 8306 10498 8318
rect 11342 8306 11394 8318
rect 15038 8370 15090 8382
rect 15038 8306 15090 8318
rect 4286 8258 4338 8270
rect 5742 8258 5794 8270
rect 9662 8258 9714 8270
rect 4498 8206 4510 8258
rect 4562 8206 4574 8258
rect 5058 8206 5070 8258
rect 5122 8206 5134 8258
rect 6066 8206 6078 8258
rect 6130 8206 6142 8258
rect 6402 8206 6414 8258
rect 6466 8206 6478 8258
rect 4286 8194 4338 8206
rect 5742 8194 5794 8206
rect 9662 8194 9714 8206
rect 11566 8258 11618 8270
rect 11566 8194 11618 8206
rect 15150 8258 15202 8270
rect 15150 8194 15202 8206
rect 15374 8258 15426 8270
rect 15374 8194 15426 8206
rect 15486 8258 15538 8270
rect 15486 8194 15538 8206
rect 15934 8258 15986 8270
rect 15934 8194 15986 8206
rect 16270 8258 16322 8270
rect 16270 8194 16322 8206
rect 16606 8258 16658 8270
rect 16606 8194 16658 8206
rect 19742 8258 19794 8270
rect 19742 8194 19794 8206
rect 20078 8258 20130 8270
rect 20514 8206 20526 8258
rect 20578 8206 20590 8258
rect 20078 8194 20130 8206
rect 5854 8146 5906 8158
rect 5854 8082 5906 8094
rect 10222 8146 10274 8158
rect 10222 8082 10274 8094
rect 11006 8146 11058 8158
rect 11006 8082 11058 8094
rect 19070 8146 19122 8158
rect 19070 8082 19122 8094
rect 19406 8146 19458 8158
rect 19406 8082 19458 8094
rect 21422 8146 21474 8158
rect 21422 8082 21474 8094
rect 21870 8146 21922 8158
rect 21870 8082 21922 8094
rect 22206 8146 22258 8158
rect 22206 8082 22258 8094
rect 5630 8034 5682 8046
rect 14590 8034 14642 8046
rect 4610 7982 4622 8034
rect 4674 7982 4686 8034
rect 14242 7982 14254 8034
rect 14306 7982 14318 8034
rect 5630 7970 5682 7982
rect 14590 7970 14642 7982
rect 16270 8034 16322 8046
rect 21310 8034 21362 8046
rect 20178 7982 20190 8034
rect 20242 7982 20254 8034
rect 16270 7970 16322 7982
rect 21310 7970 21362 7982
rect 1344 7866 22784 7900
rect 1344 7814 6534 7866
rect 6586 7814 6638 7866
rect 6690 7814 6742 7866
rect 6794 7814 11854 7866
rect 11906 7814 11958 7866
rect 12010 7814 12062 7866
rect 12114 7814 17174 7866
rect 17226 7814 17278 7866
rect 17330 7814 17382 7866
rect 17434 7814 22494 7866
rect 22546 7814 22598 7866
rect 22650 7814 22702 7866
rect 22754 7814 22784 7866
rect 1344 7780 22784 7814
rect 4734 7698 4786 7710
rect 11118 7698 11170 7710
rect 10770 7646 10782 7698
rect 10834 7646 10846 7698
rect 4734 7634 4786 7646
rect 11118 7634 11170 7646
rect 14926 7698 14978 7710
rect 19406 7698 19458 7710
rect 15250 7646 15262 7698
rect 15314 7646 15326 7698
rect 18050 7646 18062 7698
rect 18114 7646 18126 7698
rect 14926 7634 14978 7646
rect 19406 7634 19458 7646
rect 9550 7586 9602 7598
rect 9550 7522 9602 7534
rect 9886 7586 9938 7598
rect 9886 7522 9938 7534
rect 18958 7586 19010 7598
rect 18958 7522 19010 7534
rect 19966 7586 20018 7598
rect 19966 7522 20018 7534
rect 20190 7586 20242 7598
rect 20190 7522 20242 7534
rect 4622 7474 4674 7486
rect 4622 7410 4674 7422
rect 4958 7474 5010 7486
rect 9774 7474 9826 7486
rect 5170 7422 5182 7474
rect 5234 7422 5246 7474
rect 4958 7410 5010 7422
rect 9774 7410 9826 7422
rect 10110 7474 10162 7486
rect 19182 7474 19234 7486
rect 18274 7422 18286 7474
rect 18338 7422 18350 7474
rect 10110 7410 10162 7422
rect 19182 7410 19234 7422
rect 22206 7474 22258 7486
rect 22206 7410 22258 7422
rect 4846 7362 4898 7374
rect 4846 7298 4898 7310
rect 5630 7362 5682 7374
rect 5630 7298 5682 7310
rect 19070 7362 19122 7374
rect 19842 7310 19854 7362
rect 19906 7310 19918 7362
rect 19070 7298 19122 7310
rect 10334 7250 10386 7262
rect 10334 7186 10386 7198
rect 1344 7082 22624 7116
rect 1344 7030 3874 7082
rect 3926 7030 3978 7082
rect 4030 7030 4082 7082
rect 4134 7030 9194 7082
rect 9246 7030 9298 7082
rect 9350 7030 9402 7082
rect 9454 7030 14514 7082
rect 14566 7030 14618 7082
rect 14670 7030 14722 7082
rect 14774 7030 19834 7082
rect 19886 7030 19938 7082
rect 19990 7030 20042 7082
rect 20094 7030 22624 7082
rect 1344 6996 22624 7030
rect 5630 6914 5682 6926
rect 5630 6850 5682 6862
rect 10110 6914 10162 6926
rect 10110 6850 10162 6862
rect 10670 6914 10722 6926
rect 10670 6850 10722 6862
rect 5742 6802 5794 6814
rect 5742 6738 5794 6750
rect 9774 6690 9826 6702
rect 4834 6638 4846 6690
rect 4898 6638 4910 6690
rect 5954 6638 5966 6690
rect 6018 6638 6030 6690
rect 9774 6626 9826 6638
rect 10222 6690 10274 6702
rect 10222 6626 10274 6638
rect 10894 6690 10946 6702
rect 10894 6626 10946 6638
rect 11454 6690 11506 6702
rect 11454 6626 11506 6638
rect 17950 6690 18002 6702
rect 21522 6638 21534 6690
rect 21586 6638 21598 6690
rect 17950 6626 18002 6638
rect 5058 6526 5070 6578
rect 5122 6526 5134 6578
rect 9426 6526 9438 6578
rect 9490 6526 9502 6578
rect 11778 6526 11790 6578
rect 11842 6526 11854 6578
rect 15698 6526 15710 6578
rect 15762 6526 15774 6578
rect 21298 6526 21310 6578
rect 21362 6526 21374 6578
rect 11006 6466 11058 6478
rect 11006 6402 11058 6414
rect 16046 6466 16098 6478
rect 16046 6402 16098 6414
rect 17838 6466 17890 6478
rect 17838 6402 17890 6414
rect 22094 6466 22146 6478
rect 22094 6402 22146 6414
rect 1344 6298 22784 6332
rect 1344 6246 6534 6298
rect 6586 6246 6638 6298
rect 6690 6246 6742 6298
rect 6794 6246 11854 6298
rect 11906 6246 11958 6298
rect 12010 6246 12062 6298
rect 12114 6246 17174 6298
rect 17226 6246 17278 6298
rect 17330 6246 17382 6298
rect 17434 6246 22494 6298
rect 22546 6246 22598 6298
rect 22650 6246 22702 6298
rect 22754 6246 22784 6298
rect 1344 6212 22784 6246
rect 10222 6130 10274 6142
rect 11342 6130 11394 6142
rect 18510 6130 18562 6142
rect 10994 6078 11006 6130
rect 11058 6078 11070 6130
rect 17714 6078 17726 6130
rect 17778 6078 17790 6130
rect 10222 6066 10274 6078
rect 11342 6066 11394 6078
rect 18510 6066 18562 6078
rect 9886 6018 9938 6030
rect 9886 5954 9938 5966
rect 10334 6018 10386 6030
rect 10334 5954 10386 5966
rect 17938 5854 17950 5906
rect 18002 5854 18014 5906
rect 1344 5514 22624 5548
rect 1344 5462 3874 5514
rect 3926 5462 3978 5514
rect 4030 5462 4082 5514
rect 4134 5462 9194 5514
rect 9246 5462 9298 5514
rect 9350 5462 9402 5514
rect 9454 5462 14514 5514
rect 14566 5462 14618 5514
rect 14670 5462 14722 5514
rect 14774 5462 19834 5514
rect 19886 5462 19938 5514
rect 19990 5462 20042 5514
rect 20094 5462 22624 5514
rect 1344 5428 22624 5462
rect 21646 5122 21698 5134
rect 21646 5058 21698 5070
rect 22206 5122 22258 5134
rect 22206 5058 22258 5070
rect 21858 4958 21870 5010
rect 21922 4958 21934 5010
rect 1344 4730 22784 4764
rect 1344 4678 6534 4730
rect 6586 4678 6638 4730
rect 6690 4678 6742 4730
rect 6794 4678 11854 4730
rect 11906 4678 11958 4730
rect 12010 4678 12062 4730
rect 12114 4678 17174 4730
rect 17226 4678 17278 4730
rect 17330 4678 17382 4730
rect 17434 4678 22494 4730
rect 22546 4678 22598 4730
rect 22650 4678 22702 4730
rect 22754 4678 22784 4730
rect 1344 4644 22784 4678
rect 1344 3946 22624 3980
rect 1344 3894 3874 3946
rect 3926 3894 3978 3946
rect 4030 3894 4082 3946
rect 4134 3894 9194 3946
rect 9246 3894 9298 3946
rect 9350 3894 9402 3946
rect 9454 3894 14514 3946
rect 14566 3894 14618 3946
rect 14670 3894 14722 3946
rect 14774 3894 19834 3946
rect 19886 3894 19938 3946
rect 19990 3894 20042 3946
rect 20094 3894 22624 3946
rect 1344 3860 22624 3894
rect 1344 3162 22784 3196
rect 1344 3110 6534 3162
rect 6586 3110 6638 3162
rect 6690 3110 6742 3162
rect 6794 3110 11854 3162
rect 11906 3110 11958 3162
rect 12010 3110 12062 3162
rect 12114 3110 17174 3162
rect 17226 3110 17278 3162
rect 17330 3110 17382 3162
rect 17434 3110 22494 3162
rect 22546 3110 22598 3162
rect 22650 3110 22702 3162
rect 22754 3110 22784 3162
rect 1344 3076 22784 3110
<< via1 >>
rect 6534 20358 6586 20410
rect 6638 20358 6690 20410
rect 6742 20358 6794 20410
rect 11854 20358 11906 20410
rect 11958 20358 12010 20410
rect 12062 20358 12114 20410
rect 17174 20358 17226 20410
rect 17278 20358 17330 20410
rect 17382 20358 17434 20410
rect 22494 20358 22546 20410
rect 22598 20358 22650 20410
rect 22702 20358 22754 20410
rect 2046 20078 2098 20130
rect 4286 20078 4338 20130
rect 6526 20078 6578 20130
rect 9326 20078 9378 20130
rect 11006 20078 11058 20130
rect 13246 20078 13298 20130
rect 15486 20078 15538 20130
rect 17726 20078 17778 20130
rect 20190 20078 20242 20130
rect 20750 20078 20802 20130
rect 22206 20078 22258 20130
rect 2382 19966 2434 20018
rect 4510 19966 4562 20018
rect 6750 19966 6802 20018
rect 9550 19966 9602 20018
rect 11230 19966 11282 20018
rect 13582 19966 13634 20018
rect 15710 19966 15762 20018
rect 17950 19966 18002 20018
rect 19854 19966 19906 20018
rect 20974 19966 21026 20018
rect 21870 19966 21922 20018
rect 18846 19854 18898 19906
rect 18734 19742 18786 19794
rect 3874 19574 3926 19626
rect 3978 19574 4030 19626
rect 4082 19574 4134 19626
rect 9194 19574 9246 19626
rect 9298 19574 9350 19626
rect 9402 19574 9454 19626
rect 14514 19574 14566 19626
rect 14618 19574 14670 19626
rect 14722 19574 14774 19626
rect 19834 19574 19886 19626
rect 19938 19574 19990 19626
rect 20042 19574 20094 19626
rect 4510 19406 4562 19458
rect 5854 19294 5906 19346
rect 6190 19294 6242 19346
rect 6526 19294 6578 19346
rect 7534 19294 7586 19346
rect 11678 19294 11730 19346
rect 13806 19294 13858 19346
rect 18510 19294 18562 19346
rect 3054 19182 3106 19234
rect 3390 19182 3442 19234
rect 13470 19182 13522 19234
rect 15262 19182 15314 19234
rect 17950 19182 18002 19234
rect 18734 19182 18786 19234
rect 19294 19182 19346 19234
rect 21646 19182 21698 19234
rect 4622 19070 4674 19122
rect 6862 19070 6914 19122
rect 7198 19070 7250 19122
rect 10110 19070 10162 19122
rect 11454 19070 11506 19122
rect 15486 19070 15538 19122
rect 18062 19070 18114 19122
rect 18398 19070 18450 19122
rect 19182 19070 19234 19122
rect 19630 19070 19682 19122
rect 3166 18958 3218 19010
rect 3950 18958 4002 19010
rect 5966 18958 6018 19010
rect 6638 18958 6690 19010
rect 7422 18958 7474 19010
rect 9774 18958 9826 19010
rect 11678 18958 11730 19010
rect 13694 18958 13746 19010
rect 19406 18958 19458 19010
rect 21310 18958 21362 19010
rect 6534 18790 6586 18842
rect 6638 18790 6690 18842
rect 6742 18790 6794 18842
rect 11854 18790 11906 18842
rect 11958 18790 12010 18842
rect 12062 18790 12114 18842
rect 17174 18790 17226 18842
rect 17278 18790 17330 18842
rect 17382 18790 17434 18842
rect 22494 18790 22546 18842
rect 22598 18790 22650 18842
rect 22702 18790 22754 18842
rect 4062 18622 4114 18674
rect 5966 18622 6018 18674
rect 10894 18622 10946 18674
rect 14030 18622 14082 18674
rect 18622 18622 18674 18674
rect 3838 18510 3890 18562
rect 5854 18510 5906 18562
rect 7086 18510 7138 18562
rect 7982 18510 8034 18562
rect 11790 18510 11842 18562
rect 12798 18510 12850 18562
rect 15598 18510 15650 18562
rect 16606 18510 16658 18562
rect 21870 18510 21922 18562
rect 3950 18398 4002 18450
rect 4510 18398 4562 18450
rect 6190 18398 6242 18450
rect 6750 18398 6802 18450
rect 6974 18398 7026 18450
rect 7534 18398 7586 18450
rect 7646 18398 7698 18450
rect 10334 18398 10386 18450
rect 10670 18398 10722 18450
rect 11230 18398 11282 18450
rect 11454 18398 11506 18450
rect 12462 18398 12514 18450
rect 13246 18398 13298 18450
rect 13918 18398 13970 18450
rect 14142 18398 14194 18450
rect 14366 18398 14418 18450
rect 15934 18398 15986 18450
rect 16270 18398 16322 18450
rect 18286 18398 18338 18450
rect 21646 18398 21698 18450
rect 22206 18398 22258 18450
rect 2942 18286 2994 18338
rect 8430 18286 8482 18338
rect 10782 18286 10834 18338
rect 11678 18286 11730 18338
rect 3166 18174 3218 18226
rect 3502 18174 3554 18226
rect 6638 18174 6690 18226
rect 7870 18174 7922 18226
rect 13134 18174 13186 18226
rect 3874 18006 3926 18058
rect 3978 18006 4030 18058
rect 4082 18006 4134 18058
rect 9194 18006 9246 18058
rect 9298 18006 9350 18058
rect 9402 18006 9454 18058
rect 14514 18006 14566 18058
rect 14618 18006 14670 18058
rect 14722 18006 14774 18058
rect 19834 18006 19886 18058
rect 19938 18006 19990 18058
rect 20042 18006 20094 18058
rect 6862 17838 6914 17890
rect 11006 17838 11058 17890
rect 12014 17838 12066 17890
rect 19854 17838 19906 17890
rect 4510 17726 4562 17778
rect 5070 17726 5122 17778
rect 7086 17726 7138 17778
rect 19518 17726 19570 17778
rect 19966 17726 20018 17778
rect 2942 17614 2994 17666
rect 3166 17614 3218 17666
rect 3390 17614 3442 17666
rect 3502 17614 3554 17666
rect 3950 17614 4002 17666
rect 11230 17614 11282 17666
rect 20190 17614 20242 17666
rect 20302 17614 20354 17666
rect 10446 17502 10498 17554
rect 11454 17502 11506 17554
rect 11566 17502 11618 17554
rect 3614 17390 3666 17442
rect 4398 17390 4450 17442
rect 4622 17390 4674 17442
rect 6526 17390 6578 17442
rect 10670 17390 10722 17442
rect 10894 17390 10946 17442
rect 6534 17222 6586 17274
rect 6638 17222 6690 17274
rect 6742 17222 6794 17274
rect 11854 17222 11906 17274
rect 11958 17222 12010 17274
rect 12062 17222 12114 17274
rect 17174 17222 17226 17274
rect 17278 17222 17330 17274
rect 17382 17222 17434 17274
rect 22494 17222 22546 17274
rect 22598 17222 22650 17274
rect 22702 17222 22754 17274
rect 3950 17054 4002 17106
rect 11006 17054 11058 17106
rect 11118 17054 11170 17106
rect 11230 17054 11282 17106
rect 20302 17054 20354 17106
rect 3054 16942 3106 16994
rect 9662 16942 9714 16994
rect 11342 16942 11394 16994
rect 15038 16942 15090 16994
rect 20638 16942 20690 16994
rect 21870 16942 21922 16994
rect 3278 16830 3330 16882
rect 3614 16830 3666 16882
rect 11790 16830 11842 16882
rect 12238 16830 12290 16882
rect 15598 16830 15650 16882
rect 19406 16830 19458 16882
rect 19630 16830 19682 16882
rect 19966 16830 20018 16882
rect 20414 16830 20466 16882
rect 20974 16830 21026 16882
rect 21198 16830 21250 16882
rect 21646 16830 21698 16882
rect 22206 16830 22258 16882
rect 9550 16718 9602 16770
rect 15150 16718 15202 16770
rect 21086 16718 21138 16770
rect 3838 16606 3890 16658
rect 9886 16606 9938 16658
rect 15262 16606 15314 16658
rect 15598 16606 15650 16658
rect 15934 16606 15986 16658
rect 19742 16606 19794 16658
rect 3874 16438 3926 16490
rect 3978 16438 4030 16490
rect 4082 16438 4134 16490
rect 9194 16438 9246 16490
rect 9298 16438 9350 16490
rect 9402 16438 9454 16490
rect 14514 16438 14566 16490
rect 14618 16438 14670 16490
rect 14722 16438 14774 16490
rect 19834 16438 19886 16490
rect 19938 16438 19990 16490
rect 20042 16438 20094 16490
rect 15038 16270 15090 16322
rect 19406 16270 19458 16322
rect 19742 16270 19794 16322
rect 21310 16270 21362 16322
rect 19630 16158 19682 16210
rect 22318 16158 22370 16210
rect 4622 16046 4674 16098
rect 6190 16046 6242 16098
rect 14926 16046 14978 16098
rect 15262 16046 15314 16098
rect 15486 16046 15538 16098
rect 19182 16046 19234 16098
rect 20078 16046 20130 16098
rect 21422 16046 21474 16098
rect 4846 15934 4898 15986
rect 20414 15934 20466 15986
rect 20638 15934 20690 15986
rect 5854 15822 5906 15874
rect 20302 15822 20354 15874
rect 6534 15654 6586 15706
rect 6638 15654 6690 15706
rect 6742 15654 6794 15706
rect 11854 15654 11906 15706
rect 11958 15654 12010 15706
rect 12062 15654 12114 15706
rect 17174 15654 17226 15706
rect 17278 15654 17330 15706
rect 17382 15654 17434 15706
rect 22494 15654 22546 15706
rect 22598 15654 22650 15706
rect 22702 15654 22754 15706
rect 3390 15486 3442 15538
rect 8878 15486 8930 15538
rect 9662 15486 9714 15538
rect 9774 15486 9826 15538
rect 10446 15486 10498 15538
rect 19966 15486 20018 15538
rect 13918 15374 13970 15426
rect 14478 15374 14530 15426
rect 18174 15374 18226 15426
rect 20526 15374 20578 15426
rect 8654 15262 8706 15314
rect 8990 15262 9042 15314
rect 9550 15262 9602 15314
rect 10222 15262 10274 15314
rect 15822 15262 15874 15314
rect 19182 15262 19234 15314
rect 19518 15262 19570 15314
rect 19630 15262 19682 15314
rect 19742 15262 19794 15314
rect 20302 15262 20354 15314
rect 3502 15150 3554 15202
rect 11006 15150 11058 15202
rect 14814 15150 14866 15202
rect 17502 15150 17554 15202
rect 17614 15150 17666 15202
rect 17838 15150 17890 15202
rect 18062 15150 18114 15202
rect 20638 15150 20690 15202
rect 10782 15038 10834 15090
rect 13806 15038 13858 15090
rect 14142 15038 14194 15090
rect 14590 15038 14642 15090
rect 14926 15038 14978 15090
rect 15374 15038 15426 15090
rect 15486 15038 15538 15090
rect 15710 15038 15762 15090
rect 3874 14870 3926 14922
rect 3978 14870 4030 14922
rect 4082 14870 4134 14922
rect 9194 14870 9246 14922
rect 9298 14870 9350 14922
rect 9402 14870 9454 14922
rect 14514 14870 14566 14922
rect 14618 14870 14670 14922
rect 14722 14870 14774 14922
rect 19834 14870 19886 14922
rect 19938 14870 19990 14922
rect 20042 14870 20094 14922
rect 9214 14590 9266 14642
rect 3614 14478 3666 14530
rect 3838 14478 3890 14530
rect 4622 14478 4674 14530
rect 9326 14478 9378 14530
rect 14142 14478 14194 14530
rect 14702 14478 14754 14530
rect 8654 14366 8706 14418
rect 4174 14254 4226 14306
rect 4846 14254 4898 14306
rect 8878 14254 8930 14306
rect 9102 14254 9154 14306
rect 10334 14254 10386 14306
rect 14366 14254 14418 14306
rect 15038 14254 15090 14306
rect 6534 14086 6586 14138
rect 6638 14086 6690 14138
rect 6742 14086 6794 14138
rect 11854 14086 11906 14138
rect 11958 14086 12010 14138
rect 12062 14086 12114 14138
rect 17174 14086 17226 14138
rect 17278 14086 17330 14138
rect 17382 14086 17434 14138
rect 22494 14086 22546 14138
rect 22598 14086 22650 14138
rect 22702 14086 22754 14138
rect 4174 13918 4226 13970
rect 9662 13918 9714 13970
rect 9886 13806 9938 13858
rect 21870 13806 21922 13858
rect 3054 13694 3106 13746
rect 3502 13694 3554 13746
rect 4062 13694 4114 13746
rect 4286 13694 4338 13746
rect 4510 13694 4562 13746
rect 4958 13694 5010 13746
rect 5294 13694 5346 13746
rect 5630 13694 5682 13746
rect 5854 13694 5906 13746
rect 9998 13694 10050 13746
rect 22206 13694 22258 13746
rect 3726 13582 3778 13634
rect 5406 13582 5458 13634
rect 5966 13582 6018 13634
rect 21646 13582 21698 13634
rect 3874 13302 3926 13354
rect 3978 13302 4030 13354
rect 4082 13302 4134 13354
rect 9194 13302 9246 13354
rect 9298 13302 9350 13354
rect 9402 13302 9454 13354
rect 14514 13302 14566 13354
rect 14618 13302 14670 13354
rect 14722 13302 14774 13354
rect 19834 13302 19886 13354
rect 19938 13302 19990 13354
rect 20042 13302 20094 13354
rect 5630 13134 5682 13186
rect 8430 13134 8482 13186
rect 9214 13134 9266 13186
rect 10222 13134 10274 13186
rect 10558 13134 10610 13186
rect 14590 13134 14642 13186
rect 15038 13134 15090 13186
rect 15598 13134 15650 13186
rect 16270 13134 16322 13186
rect 18846 13134 18898 13186
rect 3502 13022 3554 13074
rect 9886 13022 9938 13074
rect 17950 13022 18002 13074
rect 4174 12910 4226 12962
rect 4398 12910 4450 12962
rect 5742 12910 5794 12962
rect 9102 12910 9154 12962
rect 10446 12910 10498 12962
rect 14814 12910 14866 12962
rect 15262 12910 15314 12962
rect 15710 12910 15762 12962
rect 15934 12910 15986 12962
rect 16158 12910 16210 12962
rect 18174 12910 18226 12962
rect 18398 12910 18450 12962
rect 14478 12798 14530 12850
rect 19070 12798 19122 12850
rect 20750 12798 20802 12850
rect 5854 12686 5906 12738
rect 8542 12686 8594 12738
rect 8766 12686 8818 12738
rect 9438 12686 9490 12738
rect 10558 12686 10610 12738
rect 19406 12686 19458 12738
rect 20638 12686 20690 12738
rect 6534 12518 6586 12570
rect 6638 12518 6690 12570
rect 6742 12518 6794 12570
rect 11854 12518 11906 12570
rect 11958 12518 12010 12570
rect 12062 12518 12114 12570
rect 17174 12518 17226 12570
rect 17278 12518 17330 12570
rect 17382 12518 17434 12570
rect 22494 12518 22546 12570
rect 22598 12518 22650 12570
rect 22702 12518 22754 12570
rect 4622 12350 4674 12402
rect 4958 12350 5010 12402
rect 8990 12350 9042 12402
rect 10446 12350 10498 12402
rect 19406 12350 19458 12402
rect 20750 12350 20802 12402
rect 21422 12350 21474 12402
rect 21534 12350 21586 12402
rect 21870 12350 21922 12402
rect 9998 12238 10050 12290
rect 19294 12238 19346 12290
rect 21646 12238 21698 12290
rect 9774 12126 9826 12178
rect 10446 12126 10498 12178
rect 11566 12126 11618 12178
rect 18062 12126 18114 12178
rect 18286 12126 18338 12178
rect 19182 12126 19234 12178
rect 19630 12126 19682 12178
rect 20302 12126 20354 12178
rect 20526 12126 20578 12178
rect 20750 12126 20802 12178
rect 21086 12126 21138 12178
rect 8430 12014 8482 12066
rect 10782 12014 10834 12066
rect 11342 12014 11394 12066
rect 8654 11902 8706 11954
rect 10558 11902 10610 11954
rect 11230 11902 11282 11954
rect 11678 11902 11730 11954
rect 17950 11902 18002 11954
rect 18398 11902 18450 11954
rect 3874 11734 3926 11786
rect 3978 11734 4030 11786
rect 4082 11734 4134 11786
rect 9194 11734 9246 11786
rect 9298 11734 9350 11786
rect 9402 11734 9454 11786
rect 14514 11734 14566 11786
rect 14618 11734 14670 11786
rect 14722 11734 14774 11786
rect 19834 11734 19886 11786
rect 19938 11734 19990 11786
rect 20042 11734 20094 11786
rect 10110 11566 10162 11618
rect 12238 11566 12290 11618
rect 12574 11566 12626 11618
rect 13918 11566 13970 11618
rect 14702 11566 14754 11618
rect 15038 11566 15090 11618
rect 17054 11566 17106 11618
rect 17166 11566 17218 11618
rect 17390 11566 17442 11618
rect 20302 11566 20354 11618
rect 20638 11566 20690 11618
rect 3726 11454 3778 11506
rect 10334 11342 10386 11394
rect 10558 11342 10610 11394
rect 12462 11342 12514 11394
rect 13694 11342 13746 11394
rect 14254 11342 14306 11394
rect 14926 11342 14978 11394
rect 15822 11342 15874 11394
rect 17614 11342 17666 11394
rect 18062 11342 18114 11394
rect 9998 11230 10050 11282
rect 13470 11230 13522 11282
rect 14590 11230 14642 11282
rect 15486 11230 15538 11282
rect 16158 11230 16210 11282
rect 16494 11230 16546 11282
rect 18398 11230 18450 11282
rect 20414 11230 20466 11282
rect 3614 11118 3666 11170
rect 12574 11118 12626 11170
rect 13582 11118 13634 11170
rect 6534 10950 6586 11002
rect 6638 10950 6690 11002
rect 6742 10950 6794 11002
rect 11854 10950 11906 11002
rect 11958 10950 12010 11002
rect 12062 10950 12114 11002
rect 17174 10950 17226 11002
rect 17278 10950 17330 11002
rect 17382 10950 17434 11002
rect 22494 10950 22546 11002
rect 22598 10950 22650 11002
rect 22702 10950 22754 11002
rect 3278 10782 3330 10834
rect 9550 10782 9602 10834
rect 14254 10782 14306 10834
rect 19854 10782 19906 10834
rect 21870 10670 21922 10722
rect 2942 10558 2994 10610
rect 3054 10558 3106 10610
rect 3390 10558 3442 10610
rect 14478 10558 14530 10610
rect 15038 10558 15090 10610
rect 15262 10558 15314 10610
rect 15598 10558 15650 10610
rect 19966 10558 20018 10610
rect 22206 10558 22258 10610
rect 3166 10446 3218 10498
rect 9662 10446 9714 10498
rect 15374 10446 15426 10498
rect 21646 10446 21698 10498
rect 3874 10166 3926 10218
rect 3978 10166 4030 10218
rect 4082 10166 4134 10218
rect 9194 10166 9246 10218
rect 9298 10166 9350 10218
rect 9402 10166 9454 10218
rect 14514 10166 14566 10218
rect 14618 10166 14670 10218
rect 14722 10166 14774 10218
rect 19834 10166 19886 10218
rect 19938 10166 19990 10218
rect 20042 10166 20094 10218
rect 3614 9998 3666 10050
rect 5630 9998 5682 10050
rect 9326 9998 9378 10050
rect 9438 9998 9490 10050
rect 20526 9998 20578 10050
rect 4958 9886 5010 9938
rect 5966 9886 6018 9938
rect 19518 9886 19570 9938
rect 2942 9774 2994 9826
rect 3838 9774 3890 9826
rect 4286 9774 4338 9826
rect 4510 9774 4562 9826
rect 9886 9774 9938 9826
rect 10110 9774 10162 9826
rect 19406 9774 19458 9826
rect 19966 9774 20018 9826
rect 20190 9774 20242 9826
rect 20750 9774 20802 9826
rect 3054 9662 3106 9714
rect 3166 9662 3218 9714
rect 5854 9662 5906 9714
rect 9550 9662 9602 9714
rect 19182 9662 19234 9714
rect 19630 9662 19682 9714
rect 20078 9662 20130 9714
rect 4398 9550 4450 9602
rect 5070 9550 5122 9602
rect 6534 9382 6586 9434
rect 6638 9382 6690 9434
rect 6742 9382 6794 9434
rect 11854 9382 11906 9434
rect 11958 9382 12010 9434
rect 12062 9382 12114 9434
rect 17174 9382 17226 9434
rect 17278 9382 17330 9434
rect 17382 9382 17434 9434
rect 22494 9382 22546 9434
rect 22598 9382 22650 9434
rect 22702 9382 22754 9434
rect 5966 9214 6018 9266
rect 10558 9214 10610 9266
rect 10782 9214 10834 9266
rect 19854 9214 19906 9266
rect 3726 9102 3778 9154
rect 3950 9102 4002 9154
rect 4734 9102 4786 9154
rect 4958 9102 5010 9154
rect 19966 9102 20018 9154
rect 3614 8990 3666 9042
rect 4174 8990 4226 9042
rect 5518 8990 5570 9042
rect 5966 8990 6018 9042
rect 6302 8990 6354 9042
rect 6526 8990 6578 9042
rect 10446 8990 10498 9042
rect 19630 8990 19682 9042
rect 5070 8878 5122 8930
rect 6078 8878 6130 8930
rect 10670 8878 10722 8930
rect 4510 8766 4562 8818
rect 9886 8766 9938 8818
rect 10110 8766 10162 8818
rect 3874 8598 3926 8650
rect 3978 8598 4030 8650
rect 4082 8598 4134 8650
rect 9194 8598 9246 8650
rect 9298 8598 9350 8650
rect 9402 8598 9454 8650
rect 14514 8598 14566 8650
rect 14618 8598 14670 8650
rect 14722 8598 14774 8650
rect 19834 8598 19886 8650
rect 19938 8598 19990 8650
rect 20042 8598 20094 8650
rect 4846 8430 4898 8482
rect 10782 8430 10834 8482
rect 20302 8430 20354 8482
rect 9886 8318 9938 8370
rect 10110 8318 10162 8370
rect 10446 8318 10498 8370
rect 11118 8318 11170 8370
rect 11342 8318 11394 8370
rect 15038 8318 15090 8370
rect 4286 8206 4338 8258
rect 4510 8206 4562 8258
rect 5070 8206 5122 8258
rect 5742 8206 5794 8258
rect 6078 8206 6130 8258
rect 6414 8206 6466 8258
rect 9662 8206 9714 8258
rect 11566 8206 11618 8258
rect 15150 8206 15202 8258
rect 15374 8206 15426 8258
rect 15486 8206 15538 8258
rect 15934 8206 15986 8258
rect 16270 8206 16322 8258
rect 16606 8206 16658 8258
rect 19742 8206 19794 8258
rect 20078 8206 20130 8258
rect 20526 8206 20578 8258
rect 5854 8094 5906 8146
rect 10222 8094 10274 8146
rect 11006 8094 11058 8146
rect 19070 8094 19122 8146
rect 19406 8094 19458 8146
rect 21422 8094 21474 8146
rect 21870 8094 21922 8146
rect 22206 8094 22258 8146
rect 4622 7982 4674 8034
rect 5630 7982 5682 8034
rect 14254 7982 14306 8034
rect 14590 7982 14642 8034
rect 16270 7982 16322 8034
rect 20190 7982 20242 8034
rect 21310 7982 21362 8034
rect 6534 7814 6586 7866
rect 6638 7814 6690 7866
rect 6742 7814 6794 7866
rect 11854 7814 11906 7866
rect 11958 7814 12010 7866
rect 12062 7814 12114 7866
rect 17174 7814 17226 7866
rect 17278 7814 17330 7866
rect 17382 7814 17434 7866
rect 22494 7814 22546 7866
rect 22598 7814 22650 7866
rect 22702 7814 22754 7866
rect 4734 7646 4786 7698
rect 10782 7646 10834 7698
rect 11118 7646 11170 7698
rect 14926 7646 14978 7698
rect 15262 7646 15314 7698
rect 18062 7646 18114 7698
rect 19406 7646 19458 7698
rect 9550 7534 9602 7586
rect 9886 7534 9938 7586
rect 18958 7534 19010 7586
rect 19966 7534 20018 7586
rect 20190 7534 20242 7586
rect 4622 7422 4674 7474
rect 4958 7422 5010 7474
rect 5182 7422 5234 7474
rect 9774 7422 9826 7474
rect 10110 7422 10162 7474
rect 18286 7422 18338 7474
rect 19182 7422 19234 7474
rect 22206 7422 22258 7474
rect 4846 7310 4898 7362
rect 5630 7310 5682 7362
rect 19070 7310 19122 7362
rect 19854 7310 19906 7362
rect 10334 7198 10386 7250
rect 3874 7030 3926 7082
rect 3978 7030 4030 7082
rect 4082 7030 4134 7082
rect 9194 7030 9246 7082
rect 9298 7030 9350 7082
rect 9402 7030 9454 7082
rect 14514 7030 14566 7082
rect 14618 7030 14670 7082
rect 14722 7030 14774 7082
rect 19834 7030 19886 7082
rect 19938 7030 19990 7082
rect 20042 7030 20094 7082
rect 5630 6862 5682 6914
rect 10110 6862 10162 6914
rect 10670 6862 10722 6914
rect 5742 6750 5794 6802
rect 4846 6638 4898 6690
rect 5966 6638 6018 6690
rect 9774 6638 9826 6690
rect 10222 6638 10274 6690
rect 10894 6638 10946 6690
rect 11454 6638 11506 6690
rect 17950 6638 18002 6690
rect 21534 6638 21586 6690
rect 5070 6526 5122 6578
rect 9438 6526 9490 6578
rect 11790 6526 11842 6578
rect 15710 6526 15762 6578
rect 21310 6526 21362 6578
rect 11006 6414 11058 6466
rect 16046 6414 16098 6466
rect 17838 6414 17890 6466
rect 22094 6414 22146 6466
rect 6534 6246 6586 6298
rect 6638 6246 6690 6298
rect 6742 6246 6794 6298
rect 11854 6246 11906 6298
rect 11958 6246 12010 6298
rect 12062 6246 12114 6298
rect 17174 6246 17226 6298
rect 17278 6246 17330 6298
rect 17382 6246 17434 6298
rect 22494 6246 22546 6298
rect 22598 6246 22650 6298
rect 22702 6246 22754 6298
rect 10222 6078 10274 6130
rect 11006 6078 11058 6130
rect 11342 6078 11394 6130
rect 17726 6078 17778 6130
rect 18510 6078 18562 6130
rect 9886 5966 9938 6018
rect 10334 5966 10386 6018
rect 17950 5854 18002 5906
rect 3874 5462 3926 5514
rect 3978 5462 4030 5514
rect 4082 5462 4134 5514
rect 9194 5462 9246 5514
rect 9298 5462 9350 5514
rect 9402 5462 9454 5514
rect 14514 5462 14566 5514
rect 14618 5462 14670 5514
rect 14722 5462 14774 5514
rect 19834 5462 19886 5514
rect 19938 5462 19990 5514
rect 20042 5462 20094 5514
rect 21646 5070 21698 5122
rect 22206 5070 22258 5122
rect 21870 4958 21922 5010
rect 6534 4678 6586 4730
rect 6638 4678 6690 4730
rect 6742 4678 6794 4730
rect 11854 4678 11906 4730
rect 11958 4678 12010 4730
rect 12062 4678 12114 4730
rect 17174 4678 17226 4730
rect 17278 4678 17330 4730
rect 17382 4678 17434 4730
rect 22494 4678 22546 4730
rect 22598 4678 22650 4730
rect 22702 4678 22754 4730
rect 3874 3894 3926 3946
rect 3978 3894 4030 3946
rect 4082 3894 4134 3946
rect 9194 3894 9246 3946
rect 9298 3894 9350 3946
rect 9402 3894 9454 3946
rect 14514 3894 14566 3946
rect 14618 3894 14670 3946
rect 14722 3894 14774 3946
rect 19834 3894 19886 3946
rect 19938 3894 19990 3946
rect 20042 3894 20094 3946
rect 6534 3110 6586 3162
rect 6638 3110 6690 3162
rect 6742 3110 6794 3162
rect 11854 3110 11906 3162
rect 11958 3110 12010 3162
rect 12062 3110 12114 3162
rect 17174 3110 17226 3162
rect 17278 3110 17330 3162
rect 17382 3110 17434 3162
rect 22494 3110 22546 3162
rect 22598 3110 22650 3162
rect 22702 3110 22754 3162
<< metal2 >>
rect 1792 23200 1904 24000
rect 4032 23200 4144 24000
rect 6272 23200 6384 24000
rect 8512 23200 8624 24000
rect 8876 23212 9380 23268
rect 1820 20188 1876 23200
rect 4060 21700 4116 23200
rect 4060 21644 4340 21700
rect 1820 20132 2100 20188
rect 2044 20130 2100 20132
rect 2044 20078 2046 20130
rect 2098 20078 2100 20130
rect 2044 20066 2100 20078
rect 4284 20130 4340 21644
rect 6300 20244 6356 23200
rect 8540 23044 8596 23200
rect 8876 23044 8932 23212
rect 8540 22988 8932 23044
rect 6532 20412 6796 20422
rect 6588 20356 6636 20412
rect 6692 20356 6740 20412
rect 6532 20346 6796 20356
rect 6300 20188 6580 20244
rect 4284 20078 4286 20130
rect 4338 20078 4340 20130
rect 4284 20066 4340 20078
rect 6524 20130 6580 20188
rect 6524 20078 6526 20130
rect 6578 20078 6580 20130
rect 6524 20066 6580 20078
rect 9324 20130 9380 23212
rect 10752 23200 10864 24000
rect 12992 23200 13104 24000
rect 15232 23200 15344 24000
rect 17472 23200 17584 24000
rect 19712 23200 19824 24000
rect 21952 23200 22064 24000
rect 10780 21700 10836 23200
rect 13020 21700 13076 23200
rect 10780 21644 11060 21700
rect 13020 21644 13300 21700
rect 9324 20078 9326 20130
rect 9378 20078 9380 20130
rect 9324 20066 9380 20078
rect 11004 20130 11060 21644
rect 11852 20412 12116 20422
rect 11908 20356 11956 20412
rect 12012 20356 12060 20412
rect 11852 20346 12116 20356
rect 11004 20078 11006 20130
rect 11058 20078 11060 20130
rect 11004 20066 11060 20078
rect 13244 20130 13300 21644
rect 15260 20188 15316 23200
rect 17172 20412 17436 20422
rect 17228 20356 17276 20412
rect 17332 20356 17380 20412
rect 17172 20346 17436 20356
rect 17500 20188 17556 23200
rect 15260 20132 15540 20188
rect 17500 20132 17780 20188
rect 13244 20078 13246 20130
rect 13298 20078 13300 20130
rect 13244 20066 13300 20078
rect 15484 20130 15540 20132
rect 15484 20078 15486 20130
rect 15538 20078 15540 20130
rect 15484 20066 15540 20078
rect 17724 20130 17780 20132
rect 17724 20078 17726 20130
rect 17778 20078 17780 20130
rect 17724 20066 17780 20078
rect 19740 20132 19796 23200
rect 20076 22036 20132 22046
rect 20076 20132 20132 21980
rect 21980 20188 22036 23200
rect 22492 20412 22756 20422
rect 22548 20356 22596 20412
rect 22652 20356 22700 20412
rect 22492 20346 22756 20356
rect 20188 20132 20244 20142
rect 20076 20130 20244 20132
rect 20076 20078 20190 20130
rect 20242 20078 20244 20130
rect 20076 20076 20244 20078
rect 19740 20066 19796 20076
rect 20188 20066 20244 20076
rect 20748 20132 20804 20142
rect 21980 20132 22260 20188
rect 20748 20038 20804 20076
rect 22204 20130 22260 20132
rect 22204 20078 22206 20130
rect 22258 20078 22260 20130
rect 22204 20066 22260 20078
rect 2380 20018 2436 20030
rect 2380 19966 2382 20018
rect 2434 19966 2436 20018
rect 2380 13748 2436 19966
rect 4508 20018 4564 20030
rect 4508 19966 4510 20018
rect 4562 19966 4564 20018
rect 3872 19628 4136 19638
rect 3928 19572 3976 19628
rect 4032 19572 4080 19628
rect 3872 19562 4136 19572
rect 4508 19458 4564 19966
rect 4508 19406 4510 19458
rect 4562 19406 4564 19458
rect 4508 19394 4564 19406
rect 6748 20018 6804 20030
rect 6748 19966 6750 20018
rect 6802 19966 6804 20018
rect 5852 19346 5908 19358
rect 5852 19294 5854 19346
rect 5906 19294 5908 19346
rect 3052 19236 3108 19246
rect 3052 19142 3108 19180
rect 3388 19234 3444 19246
rect 3388 19182 3390 19234
rect 3442 19182 3444 19234
rect 3164 19010 3220 19022
rect 3164 18958 3166 19010
rect 3218 18958 3220 19010
rect 3164 18564 3220 18958
rect 3164 18498 3220 18508
rect 3388 19012 3444 19182
rect 4172 19236 4228 19246
rect 3948 19012 4004 19022
rect 3388 19010 4004 19012
rect 3388 18958 3950 19010
rect 4002 18958 4004 19010
rect 3388 18956 4004 18958
rect 2940 18338 2996 18350
rect 2940 18286 2942 18338
rect 2994 18286 2996 18338
rect 2940 17666 2996 18286
rect 3164 18226 3220 18238
rect 3164 18174 3166 18226
rect 3218 18174 3220 18226
rect 2940 17614 2942 17666
rect 2994 17614 2996 17666
rect 2940 16100 2996 17614
rect 3052 17892 3108 17902
rect 3052 16994 3108 17836
rect 3052 16942 3054 16994
rect 3106 16942 3108 16994
rect 3052 16930 3108 16942
rect 3164 17666 3220 18174
rect 3164 17614 3166 17666
rect 3218 17614 3220 17666
rect 3164 17444 3220 17614
rect 3388 18228 3444 18956
rect 3948 18946 4004 18956
rect 3724 18732 4116 18788
rect 3388 17666 3444 18172
rect 3500 18226 3556 18238
rect 3500 18174 3502 18226
rect 3554 18174 3556 18226
rect 3500 17892 3556 18174
rect 3724 17892 3780 18732
rect 4060 18674 4116 18732
rect 4060 18622 4062 18674
rect 4114 18622 4116 18674
rect 4060 18610 4116 18622
rect 3836 18564 3892 18574
rect 3836 18470 3892 18508
rect 3948 18452 4004 18462
rect 4172 18452 4228 19180
rect 4620 19124 4676 19134
rect 4620 19030 4676 19068
rect 5852 18562 5908 19294
rect 6188 19348 6244 19358
rect 6524 19348 6580 19358
rect 6188 19346 6580 19348
rect 6188 19294 6190 19346
rect 6242 19294 6526 19346
rect 6578 19294 6580 19346
rect 6188 19292 6580 19294
rect 6188 19282 6244 19292
rect 5852 18510 5854 18562
rect 5906 18510 5908 18562
rect 5852 18498 5908 18510
rect 5964 19010 6020 19022
rect 5964 18958 5966 19010
rect 6018 18958 6020 19010
rect 5964 18674 6020 18958
rect 5964 18622 5966 18674
rect 6018 18622 6020 18674
rect 3948 18450 4340 18452
rect 3948 18398 3950 18450
rect 4002 18398 4340 18450
rect 3948 18396 4340 18398
rect 3948 18386 4004 18396
rect 3872 18060 4136 18070
rect 3928 18004 3976 18060
rect 4032 18004 4080 18060
rect 3872 17994 4136 18004
rect 3500 17836 4116 17892
rect 3388 17614 3390 17666
rect 3442 17614 3444 17666
rect 3388 17602 3444 17614
rect 3500 17668 3556 17706
rect 3500 17602 3556 17612
rect 3948 17666 4004 17678
rect 3948 17614 3950 17666
rect 4002 17614 4004 17666
rect 2940 16034 2996 16044
rect 3164 15204 3220 17388
rect 3612 17442 3668 17454
rect 3612 17390 3614 17442
rect 3666 17390 3668 17442
rect 3612 17332 3668 17390
rect 3948 17332 4004 17614
rect 3612 17276 4004 17332
rect 3948 17106 4004 17276
rect 3948 17054 3950 17106
rect 4002 17054 4004 17106
rect 3948 17042 4004 17054
rect 3276 16882 3332 16894
rect 3276 16830 3278 16882
rect 3330 16830 3332 16882
rect 3276 15540 3332 16830
rect 3612 16884 3668 16894
rect 4060 16884 4116 17836
rect 3612 16882 4116 16884
rect 3612 16830 3614 16882
rect 3666 16830 4116 16882
rect 3612 16828 4116 16830
rect 3612 16818 3668 16828
rect 3836 16660 3892 16670
rect 3724 16658 3892 16660
rect 3724 16606 3838 16658
rect 3890 16606 3892 16658
rect 3724 16604 3892 16606
rect 3388 15540 3444 15550
rect 3276 15538 3444 15540
rect 3276 15486 3390 15538
rect 3442 15486 3444 15538
rect 3276 15484 3444 15486
rect 3388 15474 3444 15484
rect 3164 15148 3444 15204
rect 2380 13682 2436 13692
rect 3052 14196 3108 14206
rect 3052 13748 3108 14140
rect 3052 13654 3108 13692
rect 3388 11060 3444 15148
rect 3500 15202 3556 15214
rect 3500 15150 3502 15202
rect 3554 15150 3556 15202
rect 3500 14084 3556 15150
rect 3612 14532 3668 14542
rect 3612 14438 3668 14476
rect 3724 14084 3780 16604
rect 3836 16594 3892 16604
rect 3872 16492 4136 16502
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 3872 16426 4136 16436
rect 3872 14924 4136 14934
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 3872 14858 4136 14868
rect 3836 14530 3892 14542
rect 3836 14478 3838 14530
rect 3890 14478 3892 14530
rect 3836 14308 3892 14478
rect 3836 14242 3892 14252
rect 4172 14308 4228 14346
rect 4172 14242 4228 14252
rect 3500 14028 3668 14084
rect 3724 14028 4228 14084
rect 3500 13860 3556 13870
rect 3500 13746 3556 13804
rect 3500 13694 3502 13746
rect 3554 13694 3556 13746
rect 3500 13074 3556 13694
rect 3500 13022 3502 13074
rect 3554 13022 3556 13074
rect 3500 13010 3556 13022
rect 3612 11396 3668 14028
rect 4172 13970 4228 14028
rect 4172 13918 4174 13970
rect 4226 13918 4228 13970
rect 4172 13906 4228 13918
rect 4060 13746 4116 13758
rect 4060 13694 4062 13746
rect 4114 13694 4116 13746
rect 3724 13636 3780 13646
rect 4060 13636 4116 13694
rect 4284 13748 4340 18396
rect 4508 18450 4564 18462
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 4508 17778 4564 18398
rect 5964 18452 6020 18622
rect 5964 18386 6020 18396
rect 6188 18450 6244 18462
rect 6188 18398 6190 18450
rect 6242 18398 6244 18450
rect 4508 17726 4510 17778
rect 4562 17726 4564 17778
rect 4508 17714 4564 17726
rect 5068 18228 5124 18238
rect 6188 18228 6244 18398
rect 6412 18452 6468 19292
rect 6524 19282 6580 19292
rect 6748 19236 6804 19966
rect 9548 20018 9604 20030
rect 11228 20020 11284 20030
rect 9548 19966 9550 20018
rect 9602 19966 9604 20018
rect 9192 19628 9456 19638
rect 9248 19572 9296 19628
rect 9352 19572 9400 19628
rect 9192 19562 9456 19572
rect 6748 19170 6804 19180
rect 7532 19346 7588 19358
rect 7532 19294 7534 19346
rect 7586 19294 7588 19346
rect 6860 19122 6916 19134
rect 6860 19070 6862 19122
rect 6914 19070 6916 19122
rect 6636 19012 6692 19050
rect 6636 18946 6692 18956
rect 6532 18844 6796 18854
rect 6588 18788 6636 18844
rect 6692 18788 6740 18844
rect 6532 18778 6796 18788
rect 6748 18452 6804 18462
rect 6412 18450 6804 18452
rect 6412 18398 6750 18450
rect 6802 18398 6804 18450
rect 6412 18396 6804 18398
rect 6748 18386 6804 18396
rect 6860 18340 6916 19070
rect 7196 19122 7252 19134
rect 7196 19070 7198 19122
rect 7250 19070 7252 19122
rect 7084 19012 7140 19022
rect 7196 19012 7252 19070
rect 7420 19012 7476 19022
rect 7140 18956 7252 19012
rect 7308 18956 7420 19012
rect 7084 18562 7140 18956
rect 7084 18510 7086 18562
rect 7138 18510 7140 18562
rect 7084 18498 7140 18510
rect 6972 18452 7028 18462
rect 6972 18358 7028 18396
rect 6636 18228 6692 18238
rect 6188 18226 6692 18228
rect 6188 18174 6638 18226
rect 6690 18174 6692 18226
rect 6188 18172 6692 18174
rect 5068 17778 5124 18172
rect 5068 17726 5070 17778
rect 5122 17726 5124 17778
rect 5068 17714 5124 17726
rect 4396 17442 4452 17454
rect 4396 17390 4398 17442
rect 4450 17390 4452 17442
rect 4396 16324 4452 17390
rect 4620 17444 4676 17454
rect 6524 17444 6580 17454
rect 4620 17350 4676 17388
rect 6188 17442 6580 17444
rect 6188 17390 6526 17442
rect 6578 17390 6580 17442
rect 6188 17388 6580 17390
rect 4396 16258 4452 16268
rect 4844 16324 4900 16334
rect 4620 16100 4676 16110
rect 4620 16006 4676 16044
rect 4844 15986 4900 16268
rect 4844 15934 4846 15986
rect 4898 15934 4900 15986
rect 4844 15922 4900 15934
rect 5292 16324 5348 16334
rect 4620 14530 4676 14542
rect 4620 14478 4622 14530
rect 4674 14478 4676 14530
rect 4620 14420 4676 14478
rect 4620 14354 4676 14364
rect 4844 14532 4900 14542
rect 4844 14306 4900 14476
rect 4844 14254 4846 14306
rect 4898 14254 4900 14306
rect 4284 13654 4340 13692
rect 4508 14196 4564 14206
rect 4508 13746 4564 14140
rect 4508 13694 4510 13746
rect 4562 13694 4564 13746
rect 4508 13682 4564 13694
rect 4844 13748 4900 14254
rect 4956 13748 5012 13758
rect 4844 13746 5012 13748
rect 4844 13694 4958 13746
rect 5010 13694 5012 13746
rect 4844 13692 5012 13694
rect 3724 13634 4116 13636
rect 3724 13582 3726 13634
rect 3778 13582 4116 13634
rect 3724 13580 4116 13582
rect 3724 13570 3780 13580
rect 4060 13524 4116 13580
rect 4732 13524 4788 13534
rect 4060 13468 4340 13524
rect 3872 13356 4136 13366
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 3872 13290 4136 13300
rect 4172 13188 4228 13198
rect 4172 12962 4228 13132
rect 4172 12910 4174 12962
rect 4226 12910 4228 12962
rect 4172 12898 4228 12910
rect 4284 12180 4340 13468
rect 4396 12962 4452 12974
rect 4396 12910 4398 12962
rect 4450 12910 4452 12962
rect 4396 12628 4452 12910
rect 4396 12562 4452 12572
rect 4284 12114 4340 12124
rect 4396 12404 4452 12414
rect 3872 11788 4136 11798
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 3872 11722 4136 11732
rect 4396 11620 4452 12348
rect 4620 12404 4676 12442
rect 4620 12338 4676 12348
rect 3724 11564 4452 11620
rect 4508 12292 4564 12302
rect 3724 11506 3780 11564
rect 3724 11454 3726 11506
rect 3778 11454 3780 11506
rect 3724 11442 3780 11454
rect 3612 11330 3668 11340
rect 3612 11172 3668 11182
rect 3612 11170 3780 11172
rect 3612 11118 3614 11170
rect 3666 11118 3780 11170
rect 3612 11116 3780 11118
rect 3612 11106 3668 11116
rect 3388 10994 3444 11004
rect 3612 10948 3668 10958
rect 3276 10836 3332 10874
rect 3276 10770 3332 10780
rect 2940 10724 2996 10734
rect 2940 10610 2996 10668
rect 2940 10558 2942 10610
rect 2994 10558 2996 10610
rect 2940 9826 2996 10558
rect 2940 9774 2942 9826
rect 2994 9774 2996 9826
rect 2940 9762 2996 9774
rect 3052 10610 3108 10622
rect 3052 10558 3054 10610
rect 3106 10558 3108 10610
rect 3052 9714 3108 10558
rect 3388 10610 3444 10622
rect 3388 10558 3390 10610
rect 3442 10558 3444 10610
rect 3164 10498 3220 10510
rect 3164 10446 3166 10498
rect 3218 10446 3220 10498
rect 3164 10052 3220 10446
rect 3164 9986 3220 9996
rect 3388 9828 3444 10558
rect 3612 10050 3668 10892
rect 3612 9998 3614 10050
rect 3666 9998 3668 10050
rect 3612 9986 3668 9998
rect 3724 10724 3780 11116
rect 3388 9762 3444 9772
rect 3052 9662 3054 9714
rect 3106 9662 3108 9714
rect 3052 8820 3108 9662
rect 3052 8754 3108 8764
rect 3164 9716 3220 9726
rect 3164 8148 3220 9660
rect 3724 9154 3780 10668
rect 4284 10836 4340 10846
rect 4508 10836 4564 12236
rect 4340 10780 4564 10836
rect 4620 12180 4676 12190
rect 3872 10220 4136 10230
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 3872 10154 4136 10164
rect 3836 10052 3892 10062
rect 3836 9826 3892 9996
rect 3836 9774 3838 9826
rect 3890 9774 3892 9826
rect 3836 9762 3892 9774
rect 4284 9826 4340 10780
rect 4284 9774 4286 9826
rect 4338 9774 4340 9826
rect 4284 9762 4340 9774
rect 4508 9828 4564 9838
rect 4620 9828 4676 12124
rect 4732 11508 4788 13468
rect 4844 11732 4900 13692
rect 4956 13682 5012 13692
rect 5292 13746 5348 16268
rect 6188 16098 6244 17388
rect 6524 17378 6580 17388
rect 6636 17444 6692 18172
rect 6860 17890 6916 18284
rect 6860 17838 6862 17890
rect 6914 17838 6916 17890
rect 6860 17826 6916 17838
rect 7084 17780 7140 17790
rect 7308 17780 7364 18956
rect 7420 18918 7476 18956
rect 7532 18450 7588 19294
rect 7980 19012 8036 19022
rect 7980 18562 8036 18956
rect 9548 19012 9604 19966
rect 11116 20018 11284 20020
rect 11116 19966 11230 20018
rect 11282 19966 11284 20018
rect 11116 19964 11284 19966
rect 11116 19460 11172 19964
rect 11228 19954 11284 19964
rect 13580 20020 13636 20030
rect 15708 20020 15764 20030
rect 13580 19926 13636 19964
rect 15596 20018 15764 20020
rect 15596 19966 15710 20018
rect 15762 19966 15764 20018
rect 15596 19964 15764 19966
rect 10108 19404 11172 19460
rect 11340 19908 11396 19918
rect 10108 19122 10164 19404
rect 11340 19348 11396 19852
rect 13692 19796 13748 19806
rect 10108 19070 10110 19122
rect 10162 19070 10164 19122
rect 10108 19058 10164 19070
rect 10780 19292 11396 19348
rect 11676 19346 11732 19358
rect 11676 19294 11678 19346
rect 11730 19294 11732 19346
rect 10780 19124 10836 19292
rect 11676 19236 11732 19294
rect 11564 19180 11676 19236
rect 11452 19124 11508 19134
rect 9548 18946 9604 18956
rect 9772 19010 9828 19022
rect 9772 18958 9774 19010
rect 9826 18958 9828 19010
rect 7980 18510 7982 18562
rect 8034 18510 8036 18562
rect 7980 18498 8036 18510
rect 7532 18398 7534 18450
rect 7586 18398 7588 18450
rect 7532 18386 7588 18398
rect 7644 18452 7700 18462
rect 7644 18358 7700 18396
rect 8428 18338 8484 18350
rect 8428 18286 8430 18338
rect 8482 18286 8484 18338
rect 7868 18228 7924 18238
rect 7868 18134 7924 18172
rect 8428 18228 8484 18286
rect 8428 18162 8484 18172
rect 9192 18060 9456 18070
rect 9248 18004 9296 18060
rect 9352 18004 9400 18060
rect 9192 17994 9456 18004
rect 7084 17778 7364 17780
rect 7084 17726 7086 17778
rect 7138 17726 7364 17778
rect 7084 17724 7364 17726
rect 7084 17714 7140 17724
rect 6636 17378 6692 17388
rect 8428 17444 8484 17454
rect 6532 17276 6796 17286
rect 6588 17220 6636 17276
rect 6692 17220 6740 17276
rect 6532 17210 6796 17220
rect 6188 16046 6190 16098
rect 6242 16046 6244 16098
rect 6188 16034 6244 16046
rect 5852 15874 5908 15886
rect 5852 15822 5854 15874
rect 5906 15822 5908 15874
rect 5852 15148 5908 15822
rect 6532 15708 6796 15718
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6532 15642 6796 15652
rect 5292 13694 5294 13746
rect 5346 13694 5348 13746
rect 5292 13682 5348 13694
rect 5516 15092 5908 15148
rect 5404 13636 5460 13646
rect 5404 13542 5460 13580
rect 5516 13524 5572 15092
rect 6076 14420 6132 14430
rect 5628 13748 5684 13758
rect 5852 13748 5908 13758
rect 5628 13746 5908 13748
rect 5628 13694 5630 13746
rect 5682 13694 5854 13746
rect 5906 13694 5908 13746
rect 5628 13692 5908 13694
rect 5628 13682 5684 13692
rect 5852 13682 5908 13692
rect 5516 13458 5572 13468
rect 5964 13634 6020 13646
rect 5964 13582 5966 13634
rect 6018 13582 6020 13634
rect 5628 13188 5684 13198
rect 5964 13188 6020 13582
rect 5628 13186 6020 13188
rect 5628 13134 5630 13186
rect 5682 13134 6020 13186
rect 5628 13132 6020 13134
rect 4956 12852 5012 12862
rect 4956 12402 5012 12796
rect 4956 12350 4958 12402
rect 5010 12350 5012 12402
rect 4956 12338 5012 12350
rect 4844 11676 5124 11732
rect 4732 11452 5012 11508
rect 4564 9772 4676 9828
rect 4956 9938 5012 11452
rect 5068 10052 5124 11676
rect 5628 10276 5684 13132
rect 6076 13076 6132 14364
rect 6532 14140 6796 14150
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6532 14074 6796 14084
rect 5740 13020 6132 13076
rect 6188 13636 6244 13646
rect 5740 12962 5796 13020
rect 5740 12910 5742 12962
rect 5794 12910 5796 12962
rect 5740 12898 5796 12910
rect 5404 10220 5684 10276
rect 5852 12740 5908 12750
rect 6188 12740 6244 13580
rect 8428 13186 8484 17388
rect 9548 17444 9604 17454
rect 8876 16772 8932 16782
rect 8876 16100 8932 16716
rect 9548 16770 9604 17388
rect 9660 16996 9716 17006
rect 9660 16902 9716 16940
rect 9772 16772 9828 18958
rect 10332 18450 10388 18462
rect 10332 18398 10334 18450
rect 10386 18398 10388 18450
rect 10332 17444 10388 18398
rect 10668 18450 10724 18462
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 10668 17668 10724 18398
rect 10780 18338 10836 19068
rect 11004 19122 11508 19124
rect 11004 19070 11454 19122
rect 11506 19070 11508 19122
rect 11004 19068 11508 19070
rect 10892 18676 10948 18686
rect 10892 18582 10948 18620
rect 10780 18286 10782 18338
rect 10834 18286 10836 18338
rect 10780 18274 10836 18286
rect 10892 18340 10948 18350
rect 10556 17612 10724 17668
rect 10892 17668 10948 18284
rect 11004 17890 11060 19068
rect 11452 19058 11508 19068
rect 11228 18450 11284 18462
rect 11452 18452 11508 18462
rect 11564 18452 11620 19180
rect 11676 19170 11732 19180
rect 13468 19236 13524 19246
rect 13468 19142 13524 19180
rect 11676 19010 11732 19022
rect 11676 18958 11678 19010
rect 11730 18958 11732 19010
rect 11676 18564 11732 18958
rect 13692 19010 13748 19740
rect 14512 19628 14776 19638
rect 14568 19572 14616 19628
rect 14672 19572 14720 19628
rect 14512 19562 14776 19572
rect 13804 19348 13860 19358
rect 13804 19346 13972 19348
rect 13804 19294 13806 19346
rect 13858 19294 13972 19346
rect 13804 19292 13972 19294
rect 13804 19282 13860 19292
rect 13692 18958 13694 19010
rect 13746 18958 13748 19010
rect 11852 18844 12116 18854
rect 11908 18788 11956 18844
rect 12012 18788 12060 18844
rect 11852 18778 12116 18788
rect 13692 18676 13748 18958
rect 13692 18610 13748 18620
rect 11788 18564 11844 18574
rect 11676 18562 11844 18564
rect 11676 18510 11790 18562
rect 11842 18510 11844 18562
rect 11676 18508 11844 18510
rect 11788 18498 11844 18508
rect 12796 18562 12852 18574
rect 12796 18510 12798 18562
rect 12850 18510 12852 18562
rect 12460 18452 12516 18462
rect 11228 18398 11230 18450
rect 11282 18398 11284 18450
rect 11228 18340 11284 18398
rect 11228 18274 11284 18284
rect 11340 18450 11620 18452
rect 11340 18398 11454 18450
rect 11506 18398 11620 18450
rect 11340 18396 11620 18398
rect 12012 18450 12516 18452
rect 12012 18398 12462 18450
rect 12514 18398 12516 18450
rect 12012 18396 12516 18398
rect 12796 18452 12852 18510
rect 13244 18452 13300 18462
rect 12796 18396 13244 18452
rect 11004 17838 11006 17890
rect 11058 17838 11060 17890
rect 11004 17826 11060 17838
rect 10892 17612 11060 17668
rect 10332 17378 10388 17388
rect 10444 17554 10500 17566
rect 10444 17502 10446 17554
rect 10498 17502 10500 17554
rect 9548 16718 9550 16770
rect 9602 16718 9604 16770
rect 9548 16706 9604 16718
rect 9660 16716 9828 16772
rect 10444 16772 10500 17502
rect 9192 16492 9456 16502
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9192 16426 9456 16436
rect 8876 15538 8932 16044
rect 9660 15988 9716 16716
rect 10444 16706 10500 16716
rect 9884 16658 9940 16670
rect 9884 16606 9886 16658
rect 9938 16606 9940 16658
rect 8876 15486 8878 15538
rect 8930 15486 8932 15538
rect 8876 15474 8932 15486
rect 9100 15932 9716 15988
rect 9772 16548 9828 16558
rect 8652 15316 8708 15326
rect 8988 15316 9044 15326
rect 8652 15314 9044 15316
rect 8652 15262 8654 15314
rect 8706 15262 8990 15314
rect 9042 15262 9044 15314
rect 8652 15260 9044 15262
rect 8652 15148 8708 15260
rect 8988 15250 9044 15260
rect 9100 15148 9156 15932
rect 9772 15876 9828 16492
rect 9660 15820 9828 15876
rect 9660 15538 9716 15820
rect 9660 15486 9662 15538
rect 9714 15486 9716 15538
rect 9660 15474 9716 15486
rect 9772 15540 9828 15550
rect 9884 15540 9940 16606
rect 9772 15538 9940 15540
rect 9772 15486 9774 15538
rect 9826 15486 9940 15538
rect 9772 15484 9940 15486
rect 10444 15540 10500 15550
rect 10556 15540 10612 17612
rect 10668 17444 10724 17454
rect 10668 17350 10724 17388
rect 10892 17442 10948 17454
rect 10892 17390 10894 17442
rect 10946 17390 10948 17442
rect 10892 16996 10948 17390
rect 10892 16930 10948 16940
rect 11004 17106 11060 17612
rect 11228 17666 11284 17678
rect 11228 17614 11230 17666
rect 11282 17614 11284 17666
rect 11004 17054 11006 17106
rect 11058 17054 11060 17106
rect 11004 16884 11060 17054
rect 11116 17556 11172 17566
rect 11116 17106 11172 17500
rect 11228 17444 11284 17614
rect 11228 17378 11284 17388
rect 11340 17220 11396 18396
rect 11452 18386 11508 18396
rect 11676 18340 11732 18350
rect 11676 18246 11732 18284
rect 12012 17890 12068 18396
rect 12460 18386 12516 18396
rect 13244 18358 13300 18396
rect 13916 18450 13972 19292
rect 15260 19234 15316 19246
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 14028 18676 14084 18686
rect 14028 18582 14084 18620
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13916 18386 13972 18398
rect 14140 18452 14196 18462
rect 14140 18358 14196 18396
rect 14364 18452 14420 18462
rect 14364 18358 14420 18396
rect 12012 17838 12014 17890
rect 12066 17838 12068 17890
rect 12012 17826 12068 17838
rect 13132 18226 13188 18238
rect 13132 18174 13134 18226
rect 13186 18174 13188 18226
rect 11116 17054 11118 17106
rect 11170 17054 11172 17106
rect 11116 17042 11172 17054
rect 11228 17164 11396 17220
rect 11452 17554 11508 17566
rect 11452 17502 11454 17554
rect 11506 17502 11508 17554
rect 11228 17106 11284 17164
rect 11228 17054 11230 17106
rect 11282 17054 11284 17106
rect 11228 17042 11284 17054
rect 11004 16818 11060 16828
rect 11340 16994 11396 17006
rect 11340 16942 11342 16994
rect 11394 16942 11396 16994
rect 11340 16884 11396 16942
rect 10444 15538 10612 15540
rect 10444 15486 10446 15538
rect 10498 15486 10612 15538
rect 10444 15484 10612 15486
rect 8428 13134 8430 13186
rect 8482 13134 8484 13186
rect 8428 13122 8484 13134
rect 8540 15092 8708 15148
rect 8764 15092 9156 15148
rect 9548 15314 9604 15326
rect 9548 15262 9550 15314
rect 9602 15262 9604 15314
rect 5852 12738 6244 12740
rect 5852 12686 5854 12738
rect 5906 12686 6244 12738
rect 5852 12684 6244 12686
rect 8540 12740 8596 15092
rect 8652 14420 8708 14430
rect 8652 14326 8708 14364
rect 8764 12964 8820 15092
rect 9192 14924 9456 14934
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9192 14858 9456 14868
rect 9548 14756 9604 15262
rect 9212 14700 9604 14756
rect 9212 14642 9268 14700
rect 9212 14590 9214 14642
rect 9266 14590 9268 14642
rect 9212 14578 9268 14590
rect 9100 14532 9156 14542
rect 8988 14476 9100 14532
rect 8876 14308 8932 14318
rect 8876 14214 8932 14252
rect 8764 12908 8932 12964
rect 5068 9996 5236 10052
rect 4956 9886 4958 9938
rect 5010 9886 5012 9938
rect 4508 9734 4564 9772
rect 4956 9716 5012 9886
rect 4732 9660 5012 9716
rect 4396 9602 4452 9614
rect 4396 9550 4398 9602
rect 4450 9550 4452 9602
rect 3724 9102 3726 9154
rect 3778 9102 3780 9154
rect 3724 9090 3780 9102
rect 3948 9156 4004 9166
rect 3948 9062 4004 9100
rect 3612 9044 3668 9054
rect 3612 8950 3668 8988
rect 4172 9042 4228 9054
rect 4172 8990 4174 9042
rect 4226 8990 4228 9042
rect 4172 8820 4228 8990
rect 4396 9044 4452 9550
rect 4732 9154 4788 9660
rect 5068 9604 5124 9614
rect 5068 9510 5124 9548
rect 4732 9102 4734 9154
rect 4786 9102 4788 9154
rect 4732 9090 4788 9102
rect 4844 9268 4900 9278
rect 4396 8988 4676 9044
rect 4508 8820 4564 8830
rect 4172 8754 4228 8764
rect 4284 8818 4564 8820
rect 4284 8766 4510 8818
rect 4562 8766 4564 8818
rect 4284 8764 4564 8766
rect 3872 8652 4136 8662
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 3872 8586 4136 8596
rect 4284 8258 4340 8764
rect 4508 8754 4564 8764
rect 4284 8206 4286 8258
rect 4338 8206 4340 8258
rect 4284 8194 4340 8206
rect 4508 8596 4564 8606
rect 4508 8258 4564 8540
rect 4620 8484 4676 8988
rect 4620 8428 4788 8484
rect 4508 8206 4510 8258
rect 4562 8206 4564 8258
rect 4508 8194 4564 8206
rect 3164 8082 3220 8092
rect 4620 8034 4676 8046
rect 4620 7982 4622 8034
rect 4674 7982 4676 8034
rect 4620 7474 4676 7982
rect 4732 7698 4788 8428
rect 4844 8482 4900 9212
rect 4956 9156 5012 9166
rect 5180 9156 5236 9996
rect 4956 9154 5236 9156
rect 4956 9102 4958 9154
rect 5010 9102 5236 9154
rect 4956 9100 5236 9102
rect 4956 9044 5012 9100
rect 4956 8978 5012 8988
rect 5068 8932 5124 8942
rect 5068 8838 5124 8876
rect 4844 8430 4846 8482
rect 4898 8430 4900 8482
rect 4844 8418 4900 8430
rect 5068 8260 5124 8270
rect 5068 8166 5124 8204
rect 4732 7646 4734 7698
rect 4786 7646 4788 7698
rect 4732 7634 4788 7646
rect 4620 7422 4622 7474
rect 4674 7422 4676 7474
rect 4620 7410 4676 7422
rect 4956 7474 5012 7486
rect 5180 7476 5236 7486
rect 5404 7476 5460 10220
rect 5628 10052 5684 10062
rect 5852 10052 5908 12684
rect 6532 12572 6796 12582
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6532 12506 6796 12516
rect 8540 12292 8596 12684
rect 8316 12236 8596 12292
rect 8764 12738 8820 12750
rect 8764 12686 8766 12738
rect 8818 12686 8820 12738
rect 6532 11004 6796 11014
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6532 10938 6796 10948
rect 8316 10724 8372 12236
rect 8764 12180 8820 12686
rect 8876 12404 8932 12908
rect 8988 12628 9044 14476
rect 9100 14466 9156 14476
rect 9324 14530 9380 14542
rect 9324 14478 9326 14530
rect 9378 14478 9380 14530
rect 9100 14306 9156 14318
rect 9100 14254 9102 14306
rect 9154 14254 9156 14306
rect 9100 13636 9156 14254
rect 9100 13570 9156 13580
rect 9324 13524 9380 14478
rect 9772 14532 9828 15484
rect 10444 15474 10500 15484
rect 10220 15314 10276 15326
rect 10220 15262 10222 15314
rect 10274 15262 10276 15314
rect 9772 14466 9828 14476
rect 9996 15204 10052 15214
rect 9996 14084 10052 15148
rect 10220 15148 10276 15262
rect 11004 15204 11060 15242
rect 10220 15092 10388 15148
rect 11004 15138 11060 15148
rect 9772 14028 10052 14084
rect 10332 14306 10388 15092
rect 10780 15092 10836 15102
rect 10780 15090 10948 15092
rect 10780 15038 10782 15090
rect 10834 15038 10948 15090
rect 10780 15036 10948 15038
rect 10780 15026 10836 15036
rect 10332 14254 10334 14306
rect 10386 14254 10388 14306
rect 9660 13972 9716 13982
rect 9660 13878 9716 13916
rect 9772 13524 9828 14028
rect 9884 13858 9940 13870
rect 9884 13806 9886 13858
rect 9938 13806 9940 13858
rect 9884 13636 9940 13806
rect 9884 13570 9940 13580
rect 9996 13746 10052 13758
rect 9996 13694 9998 13746
rect 10050 13694 10052 13746
rect 9324 13468 9828 13524
rect 9192 13356 9456 13366
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9192 13290 9456 13300
rect 9212 13188 9268 13198
rect 9100 13186 9268 13188
rect 9100 13134 9214 13186
rect 9266 13134 9268 13186
rect 9100 13132 9268 13134
rect 9100 12962 9156 13132
rect 9212 13122 9268 13132
rect 9100 12910 9102 12962
rect 9154 12910 9156 12962
rect 9100 12898 9156 12910
rect 9212 12740 9268 12750
rect 9436 12740 9492 12750
rect 9268 12738 9492 12740
rect 9268 12686 9438 12738
rect 9490 12686 9492 12738
rect 9268 12684 9492 12686
rect 9212 12674 9268 12684
rect 9436 12674 9492 12684
rect 8988 12572 9156 12628
rect 8988 12404 9044 12414
rect 8876 12402 9044 12404
rect 8876 12350 8990 12402
rect 9042 12350 9044 12402
rect 8876 12348 9044 12350
rect 8988 12338 9044 12348
rect 8540 12124 8820 12180
rect 8428 12068 8484 12078
rect 8540 12068 8596 12124
rect 8428 12066 8596 12068
rect 8428 12014 8430 12066
rect 8482 12014 8596 12066
rect 8428 12012 8596 12014
rect 8428 12002 8484 12012
rect 8540 10836 8596 12012
rect 8652 11956 8708 11966
rect 9100 11956 9156 12572
rect 8652 11862 8708 11900
rect 8988 11900 9156 11956
rect 8540 10770 8596 10780
rect 8316 10668 8484 10724
rect 5628 10050 5908 10052
rect 5628 9998 5630 10050
rect 5682 9998 5908 10050
rect 5628 9996 5908 9998
rect 5628 9986 5684 9996
rect 5964 9940 6020 9950
rect 5964 9938 6356 9940
rect 5964 9886 5966 9938
rect 6018 9886 6356 9938
rect 5964 9884 6356 9886
rect 5964 9874 6020 9884
rect 5852 9716 5908 9726
rect 5740 9714 5908 9716
rect 5740 9662 5854 9714
rect 5906 9662 5908 9714
rect 5740 9660 5908 9662
rect 5740 9604 5796 9660
rect 5740 9538 5796 9548
rect 5516 9042 5572 9054
rect 5516 8990 5518 9042
rect 5570 8990 5572 9042
rect 5516 8932 5572 8990
rect 5516 8866 5572 8876
rect 5740 8260 5796 8270
rect 5740 8166 5796 8204
rect 5852 8146 5908 9660
rect 5964 9268 6020 9278
rect 5964 9174 6020 9212
rect 5964 9042 6020 9054
rect 5964 8990 5966 9042
rect 6018 8990 6020 9042
rect 5964 8484 6020 8990
rect 6300 9042 6356 9884
rect 6532 9436 6796 9446
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6532 9370 6796 9380
rect 6300 8990 6302 9042
rect 6354 8990 6356 9042
rect 6300 8978 6356 8990
rect 6524 9044 6580 9054
rect 6524 8950 6580 8988
rect 6076 8932 6132 8942
rect 6076 8596 6132 8876
rect 6076 8530 6132 8540
rect 6188 8820 6244 8830
rect 5964 8418 6020 8428
rect 5852 8094 5854 8146
rect 5906 8094 5908 8146
rect 5852 8082 5908 8094
rect 6076 8258 6132 8270
rect 6076 8206 6078 8258
rect 6130 8206 6132 8258
rect 6076 8148 6132 8206
rect 6076 8082 6132 8092
rect 5628 8034 5684 8046
rect 5628 7982 5630 8034
rect 5682 7982 5684 8034
rect 5628 7924 5684 7982
rect 6188 7924 6244 8764
rect 5628 7868 6244 7924
rect 6412 8258 6468 8270
rect 6412 8206 6414 8258
rect 6466 8206 6468 8258
rect 4956 7422 4958 7474
rect 5010 7422 5012 7474
rect 4844 7362 4900 7374
rect 4844 7310 4846 7362
rect 4898 7310 4900 7362
rect 3872 7084 4136 7094
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 3872 7018 4136 7028
rect 4844 7028 4900 7310
rect 4956 7364 5012 7422
rect 4956 7298 5012 7308
rect 5068 7474 5460 7476
rect 5068 7422 5182 7474
rect 5234 7422 5460 7474
rect 5068 7420 5460 7422
rect 4844 6962 4900 6972
rect 4844 6804 4900 6814
rect 4844 6690 4900 6748
rect 4844 6638 4846 6690
rect 4898 6638 4900 6690
rect 4844 6626 4900 6638
rect 5068 6578 5124 7420
rect 5180 7410 5236 7420
rect 5628 7364 5684 7374
rect 5628 7270 5684 7308
rect 5628 7028 5684 7038
rect 5628 6914 5684 6972
rect 5628 6862 5630 6914
rect 5682 6862 5684 6914
rect 5628 6850 5684 6862
rect 5740 6804 5796 6814
rect 5740 6710 5796 6748
rect 5068 6526 5070 6578
rect 5122 6526 5124 6578
rect 5068 6514 5124 6526
rect 5964 6690 6020 6702
rect 5964 6638 5966 6690
rect 6018 6638 6020 6690
rect 5964 6580 6020 6638
rect 5964 6514 6020 6524
rect 6412 6580 6468 8206
rect 6532 7868 6796 7878
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6532 7802 6796 7812
rect 6412 6514 6468 6524
rect 6532 6300 6796 6310
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6532 6234 6796 6244
rect 8428 6132 8484 10668
rect 8988 8372 9044 11900
rect 9192 11788 9456 11798
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9192 11722 9456 11732
rect 9660 11620 9716 13468
rect 9884 13074 9940 13086
rect 9884 13022 9886 13074
rect 9938 13022 9940 13074
rect 9772 12178 9828 12190
rect 9772 12126 9774 12178
rect 9826 12126 9828 12178
rect 9772 11844 9828 12126
rect 9772 11778 9828 11788
rect 9660 11564 9828 11620
rect 9548 10836 9604 10846
rect 9548 10742 9604 10780
rect 9660 10498 9716 10510
rect 9660 10446 9662 10498
rect 9714 10446 9716 10498
rect 9192 10220 9456 10230
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9192 10154 9456 10164
rect 9324 10052 9380 10062
rect 9324 9958 9380 9996
rect 9436 10050 9492 10062
rect 9436 9998 9438 10050
rect 9490 9998 9492 10050
rect 9436 8820 9492 9998
rect 9660 9828 9716 10446
rect 9772 10164 9828 11564
rect 9884 11284 9940 13022
rect 9996 12516 10052 13694
rect 10220 13524 10276 13534
rect 10220 13188 10276 13468
rect 10332 13412 10388 14254
rect 10892 14308 10948 15036
rect 10556 13412 10612 13422
rect 10332 13356 10556 13412
rect 10556 13346 10612 13356
rect 10556 13188 10612 13198
rect 9996 12450 10052 12460
rect 10108 13186 10276 13188
rect 10108 13134 10222 13186
rect 10274 13134 10276 13186
rect 10108 13132 10276 13134
rect 9996 12290 10052 12302
rect 9996 12238 9998 12290
rect 10050 12238 10052 12290
rect 9996 12180 10052 12238
rect 9996 12114 10052 12124
rect 10108 11618 10164 13132
rect 10220 13122 10276 13132
rect 10332 13186 10612 13188
rect 10332 13134 10558 13186
rect 10610 13134 10612 13186
rect 10332 13132 10612 13134
rect 10332 12180 10388 13132
rect 10556 13122 10612 13132
rect 10444 12964 10500 12974
rect 10444 12870 10500 12908
rect 10556 12740 10612 12750
rect 10892 12740 10948 14252
rect 10556 12738 10948 12740
rect 10556 12686 10558 12738
rect 10610 12686 10948 12738
rect 10556 12684 10948 12686
rect 11116 13412 11172 13422
rect 10556 12674 10612 12684
rect 10444 12516 10500 12526
rect 10444 12404 10500 12460
rect 10444 12402 10724 12404
rect 10444 12350 10446 12402
rect 10498 12350 10724 12402
rect 10444 12348 10724 12350
rect 10444 12338 10500 12348
rect 10444 12180 10500 12190
rect 10332 12124 10444 12180
rect 10444 12086 10500 12124
rect 10556 11956 10612 11966
rect 10108 11566 10110 11618
rect 10162 11566 10164 11618
rect 10108 11554 10164 11566
rect 10444 11954 10612 11956
rect 10444 11902 10558 11954
rect 10610 11902 10612 11954
rect 10444 11900 10612 11902
rect 10332 11396 10388 11406
rect 10444 11396 10500 11900
rect 10556 11890 10612 11900
rect 10332 11394 10500 11396
rect 10332 11342 10334 11394
rect 10386 11342 10500 11394
rect 10332 11340 10500 11342
rect 10556 11620 10612 11630
rect 10556 11394 10612 11564
rect 10556 11342 10558 11394
rect 10610 11342 10612 11394
rect 9996 11284 10052 11294
rect 9884 11282 10052 11284
rect 9884 11230 9998 11282
rect 10050 11230 10052 11282
rect 9884 11228 10052 11230
rect 9772 10098 9828 10108
rect 9884 9828 9940 9838
rect 9660 9772 9884 9828
rect 9884 9734 9940 9772
rect 9548 9716 9604 9726
rect 9548 9622 9604 9660
rect 9996 9604 10052 11228
rect 10332 11284 10388 11340
rect 10556 11330 10612 11342
rect 10332 11218 10388 11228
rect 9660 9548 10052 9604
rect 10108 9826 10164 9838
rect 10108 9774 10110 9826
rect 10162 9774 10164 9826
rect 9660 9492 9716 9548
rect 9436 8754 9492 8764
rect 9548 9436 9716 9492
rect 10108 9492 10164 9774
rect 10332 9828 10388 9838
rect 10108 9436 10276 9492
rect 9192 8652 9456 8662
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9192 8586 9456 8596
rect 8988 8306 9044 8316
rect 9548 7586 9604 9436
rect 9996 9156 10052 9166
rect 9884 8820 9940 8830
rect 9772 8818 9940 8820
rect 9772 8766 9886 8818
rect 9938 8766 9940 8818
rect 9772 8764 9940 8766
rect 9660 8260 9716 8270
rect 9772 8260 9828 8764
rect 9884 8754 9940 8764
rect 9884 8372 9940 8382
rect 9884 8278 9940 8316
rect 9716 8204 9828 8260
rect 9660 8166 9716 8204
rect 9548 7534 9550 7586
rect 9602 7534 9604 7586
rect 9548 7522 9604 7534
rect 9884 7588 9940 7598
rect 9996 7588 10052 9100
rect 10108 8820 10164 8830
rect 10108 8726 10164 8764
rect 10220 8596 10276 9436
rect 10332 8820 10388 9772
rect 10332 8754 10388 8764
rect 10444 9716 10500 9726
rect 10444 9042 10500 9660
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 10444 8708 10500 8990
rect 10556 9268 10612 9278
rect 10668 9268 10724 12348
rect 10780 12068 10836 12078
rect 10780 11974 10836 12012
rect 10892 11956 10948 11966
rect 10556 9266 10724 9268
rect 10556 9214 10558 9266
rect 10610 9214 10724 9266
rect 10556 9212 10724 9214
rect 10780 11172 10836 11182
rect 10780 9266 10836 11116
rect 10780 9214 10782 9266
rect 10834 9214 10836 9266
rect 10556 8708 10612 9212
rect 10780 9202 10836 9214
rect 10668 8932 10724 8942
rect 10668 8838 10724 8876
rect 10556 8652 10836 8708
rect 10444 8642 10500 8652
rect 10220 8540 10388 8596
rect 10108 8484 10164 8494
rect 10108 8370 10164 8428
rect 10108 8318 10110 8370
rect 10162 8318 10164 8370
rect 10108 8306 10164 8318
rect 10332 8260 10388 8540
rect 10444 8484 10500 8494
rect 10444 8370 10500 8428
rect 10780 8482 10836 8652
rect 10780 8430 10782 8482
rect 10834 8430 10836 8482
rect 10780 8418 10836 8430
rect 10444 8318 10446 8370
rect 10498 8318 10500 8370
rect 10444 8306 10500 8318
rect 10668 8372 10724 8382
rect 10668 8260 10724 8316
rect 10668 8204 10836 8260
rect 10220 8148 10276 8158
rect 9884 7586 10052 7588
rect 9884 7534 9886 7586
rect 9938 7534 10052 7586
rect 9884 7532 10052 7534
rect 10108 8036 10164 8046
rect 9884 7522 9940 7532
rect 9772 7474 9828 7486
rect 9772 7422 9774 7474
rect 9826 7422 9828 7474
rect 9660 7364 9716 7374
rect 9192 7084 9456 7094
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9192 7018 9456 7028
rect 9436 6916 9492 6926
rect 9436 6578 9492 6860
rect 9436 6526 9438 6578
rect 9490 6526 9492 6578
rect 9436 6514 9492 6526
rect 8540 6132 8596 6142
rect 8428 6076 8540 6132
rect 8540 6066 8596 6076
rect 9660 6020 9716 7308
rect 9772 6692 9828 7422
rect 10108 7474 10164 7980
rect 10108 7422 10110 7474
rect 10162 7422 10164 7474
rect 10108 7410 10164 7422
rect 10220 7252 10276 8092
rect 9996 7196 10276 7252
rect 10332 7252 10388 8204
rect 10668 8036 10724 8046
rect 10332 7250 10500 7252
rect 10332 7198 10334 7250
rect 10386 7198 10500 7250
rect 10332 7196 10500 7198
rect 9996 6916 10052 7196
rect 10332 7186 10388 7196
rect 9996 6850 10052 6860
rect 10108 6916 10164 6926
rect 10332 6916 10388 6926
rect 10108 6914 10332 6916
rect 10108 6862 10110 6914
rect 10162 6862 10332 6914
rect 10108 6860 10332 6862
rect 10108 6850 10164 6860
rect 10332 6850 10388 6860
rect 10220 6692 10276 6702
rect 9772 6690 10220 6692
rect 9772 6638 9774 6690
rect 9826 6638 10220 6690
rect 9772 6636 10220 6638
rect 9772 6626 9828 6636
rect 10220 6130 10276 6636
rect 10220 6078 10222 6130
rect 10274 6078 10276 6130
rect 10220 6066 10276 6078
rect 10444 6132 10500 7196
rect 10668 6914 10724 7980
rect 10780 7698 10836 8204
rect 10780 7646 10782 7698
rect 10834 7646 10836 7698
rect 10780 7634 10836 7646
rect 10668 6862 10670 6914
rect 10722 6862 10724 6914
rect 10668 6850 10724 6862
rect 10892 6916 10948 11900
rect 11116 11732 11172 13356
rect 11340 12292 11396 16828
rect 11452 16772 11508 17502
rect 11564 17556 11620 17566
rect 11564 17462 11620 17500
rect 11852 17276 12116 17286
rect 11908 17220 11956 17276
rect 12012 17220 12060 17276
rect 11852 17210 12116 17220
rect 11788 16996 11844 17006
rect 11788 16882 11844 16940
rect 13132 16996 13188 18174
rect 14512 18060 14776 18070
rect 14568 18004 14616 18060
rect 14672 18004 14720 18060
rect 14512 17994 14776 18004
rect 15260 17108 15316 19182
rect 15484 19124 15540 19134
rect 15596 19124 15652 19964
rect 15708 19954 15764 19964
rect 17948 20018 18004 20030
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17948 19796 18004 19966
rect 17948 19730 18004 19740
rect 18508 20020 18564 20030
rect 18508 19346 18564 19964
rect 19852 20018 19908 20030
rect 20972 20020 21028 20030
rect 21868 20020 21924 20030
rect 19852 19966 19854 20018
rect 19906 19966 19908 20018
rect 18844 19906 18900 19918
rect 18844 19854 18846 19906
rect 18898 19854 18900 19906
rect 18508 19294 18510 19346
rect 18562 19294 18564 19346
rect 18508 19282 18564 19294
rect 18732 19794 18788 19806
rect 18732 19742 18734 19794
rect 18786 19742 18788 19794
rect 17948 19236 18004 19246
rect 17948 19142 18004 19180
rect 18732 19234 18788 19742
rect 18732 19182 18734 19234
rect 18786 19182 18788 19234
rect 18732 19170 18788 19182
rect 18844 19460 18900 19854
rect 19852 19908 19908 19966
rect 19852 19842 19908 19852
rect 20860 20018 21028 20020
rect 20860 19966 20974 20018
rect 21026 19966 21028 20018
rect 20860 19964 21028 19966
rect 19832 19628 20096 19638
rect 19888 19572 19936 19628
rect 19992 19572 20040 19628
rect 19832 19562 20096 19572
rect 18844 19404 19684 19460
rect 15484 19122 15652 19124
rect 15484 19070 15486 19122
rect 15538 19070 15652 19122
rect 15484 19068 15652 19070
rect 18060 19124 18116 19134
rect 18396 19124 18452 19134
rect 18060 19122 18396 19124
rect 18060 19070 18062 19122
rect 18114 19070 18396 19122
rect 18060 19068 18396 19070
rect 15484 19058 15540 19068
rect 18060 19058 18116 19068
rect 18396 19030 18452 19068
rect 18844 19012 18900 19404
rect 19292 19236 19348 19246
rect 19292 19142 19348 19180
rect 19180 19124 19236 19134
rect 19180 19030 19236 19068
rect 19628 19122 19684 19404
rect 19628 19070 19630 19122
rect 19682 19070 19684 19122
rect 19628 19058 19684 19070
rect 20636 19236 20692 19246
rect 18620 18956 18900 19012
rect 19404 19012 19460 19022
rect 17172 18844 17436 18854
rect 17228 18788 17276 18844
rect 17332 18788 17380 18844
rect 17172 18778 17436 18788
rect 18620 18674 18676 18956
rect 19404 18918 19460 18956
rect 18620 18622 18622 18674
rect 18674 18622 18676 18674
rect 18620 18610 18676 18622
rect 15596 18562 15652 18574
rect 15596 18510 15598 18562
rect 15650 18510 15652 18562
rect 15596 18452 15652 18510
rect 16604 18562 16660 18574
rect 16604 18510 16606 18562
rect 16658 18510 16660 18562
rect 15596 18386 15652 18396
rect 15932 18450 15988 18462
rect 15932 18398 15934 18450
rect 15986 18398 15988 18450
rect 15932 18340 15988 18398
rect 15932 18274 15988 18284
rect 16044 18452 16100 18462
rect 15260 17052 15764 17108
rect 13132 16930 13188 16940
rect 15036 16994 15092 17006
rect 15036 16942 15038 16994
rect 15090 16942 15092 16994
rect 11788 16830 11790 16882
rect 11842 16830 11844 16882
rect 11788 16818 11844 16830
rect 12236 16884 12292 16894
rect 12236 16790 12292 16828
rect 11452 15428 11508 16716
rect 14512 16492 14776 16502
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14512 16426 14776 16436
rect 15036 16324 15092 16942
rect 15596 16884 15652 16894
rect 15036 16230 15092 16268
rect 15148 16882 15652 16884
rect 15148 16830 15598 16882
rect 15650 16830 15652 16882
rect 15148 16828 15652 16830
rect 15148 16770 15204 16828
rect 15596 16818 15652 16828
rect 15148 16718 15150 16770
rect 15202 16718 15204 16770
rect 14140 16100 14196 16110
rect 11852 15708 12116 15718
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 11852 15642 12116 15652
rect 11452 15362 11508 15372
rect 13916 15426 13972 15438
rect 13916 15374 13918 15426
rect 13970 15374 13972 15426
rect 13804 15090 13860 15102
rect 13804 15038 13806 15090
rect 13858 15038 13860 15090
rect 13804 14532 13860 15038
rect 13916 14868 13972 15374
rect 14140 15090 14196 16044
rect 14924 16100 14980 16110
rect 15148 16100 15204 16718
rect 15260 16660 15316 16670
rect 15596 16660 15652 16670
rect 15260 16658 15652 16660
rect 15260 16606 15262 16658
rect 15314 16606 15598 16658
rect 15650 16606 15652 16658
rect 15260 16604 15652 16606
rect 15260 16594 15316 16604
rect 15596 16594 15652 16604
rect 15484 16324 15540 16334
rect 15260 16100 15316 16110
rect 15148 16098 15316 16100
rect 15148 16046 15262 16098
rect 15314 16046 15316 16098
rect 15148 16044 15316 16046
rect 14924 16006 14980 16044
rect 14476 15428 14532 15438
rect 14476 15334 14532 15372
rect 15260 15316 15316 16044
rect 15484 16098 15540 16268
rect 15484 16046 15486 16098
rect 15538 16046 15540 16098
rect 15484 16034 15540 16046
rect 15708 16100 15764 17052
rect 15932 16658 15988 16670
rect 15932 16606 15934 16658
rect 15986 16606 15988 16658
rect 15932 16324 15988 16606
rect 15932 16258 15988 16268
rect 15708 16044 15988 16100
rect 15820 15316 15876 15326
rect 14812 15260 15092 15316
rect 15260 15314 15876 15316
rect 15260 15262 15822 15314
rect 15874 15262 15876 15314
rect 15260 15260 15876 15262
rect 14812 15202 14868 15260
rect 14812 15150 14814 15202
rect 14866 15150 14868 15202
rect 14812 15138 14868 15150
rect 15036 15204 15092 15260
rect 15820 15250 15876 15260
rect 14588 15092 14644 15102
rect 14140 15038 14142 15090
rect 14194 15038 14196 15090
rect 14140 15026 14196 15038
rect 14364 15090 14644 15092
rect 14364 15038 14590 15090
rect 14642 15038 14644 15090
rect 14364 15036 14644 15038
rect 14364 14868 14420 15036
rect 14588 15026 14644 15036
rect 14924 15090 14980 15102
rect 14924 15038 14926 15090
rect 14978 15038 14980 15090
rect 13916 14812 14420 14868
rect 14512 14924 14776 14934
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14512 14858 14776 14868
rect 11852 14140 12116 14150
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 11852 14074 12116 14084
rect 12236 13524 12292 13534
rect 11452 12964 11508 12974
rect 11508 12908 11620 12964
rect 11452 12898 11508 12908
rect 11340 12236 11508 12292
rect 11340 12068 11396 12078
rect 11340 11974 11396 12012
rect 11228 11956 11284 11966
rect 11228 11862 11284 11900
rect 11116 11676 11284 11732
rect 11116 9044 11172 9054
rect 11004 8708 11060 8718
rect 11004 8148 11060 8652
rect 11116 8370 11172 8988
rect 11116 8318 11118 8370
rect 11170 8318 11172 8370
rect 11116 8306 11172 8318
rect 11004 8082 11060 8092
rect 11116 8036 11172 8046
rect 10892 6850 10948 6860
rect 11004 7924 11060 7934
rect 10892 6690 10948 6702
rect 10892 6638 10894 6690
rect 10946 6638 10948 6690
rect 10892 6468 10948 6638
rect 10892 6402 10948 6412
rect 11004 6466 11060 7868
rect 11116 7698 11172 7980
rect 11116 7646 11118 7698
rect 11170 7646 11172 7698
rect 11116 7634 11172 7646
rect 11228 7588 11284 11676
rect 11340 8372 11396 8382
rect 11340 8278 11396 8316
rect 11340 7588 11396 7598
rect 11228 7532 11340 7588
rect 11340 7522 11396 7532
rect 11452 7252 11508 12236
rect 11564 12178 11620 12908
rect 11852 12572 12116 12582
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 11852 12506 12116 12516
rect 11564 12126 11566 12178
rect 11618 12126 11620 12178
rect 11564 11732 11620 12126
rect 11564 11666 11620 11676
rect 11676 11954 11732 11966
rect 11676 11902 11678 11954
rect 11730 11902 11732 11954
rect 11676 11620 11732 11902
rect 11676 11554 11732 11564
rect 12236 11618 12292 13468
rect 13804 12068 13860 14476
rect 14140 14530 14196 14542
rect 14140 14478 14142 14530
rect 14194 14478 14196 14530
rect 14140 14420 14196 14478
rect 14140 13524 14196 14364
rect 14364 14308 14420 14812
rect 14700 14532 14756 14542
rect 14700 14438 14756 14476
rect 14140 13458 14196 13468
rect 14252 14306 14420 14308
rect 14252 14254 14366 14306
rect 14418 14254 14420 14306
rect 14252 14252 14420 14254
rect 14252 13188 14308 14252
rect 14364 14242 14420 14252
rect 14476 14308 14532 14318
rect 14476 14084 14532 14252
rect 14252 13122 14308 13132
rect 14364 14028 14532 14084
rect 12236 11566 12238 11618
rect 12290 11566 12292 11618
rect 12236 11554 12292 11566
rect 12572 11732 12628 11742
rect 12572 11618 12628 11676
rect 12572 11566 12574 11618
rect 12626 11566 12628 11618
rect 12572 11554 12628 11566
rect 13692 11732 13748 11742
rect 13692 11508 13748 11676
rect 13804 11620 13860 12012
rect 13916 11620 13972 11630
rect 13804 11618 13972 11620
rect 13804 11566 13918 11618
rect 13970 11566 13972 11618
rect 13804 11564 13972 11566
rect 14364 11620 14420 14028
rect 14924 13412 14980 15038
rect 15036 14532 15092 15148
rect 15372 15090 15428 15102
rect 15372 15038 15374 15090
rect 15426 15038 15428 15090
rect 15372 14532 15428 15038
rect 15484 15090 15540 15102
rect 15484 15038 15486 15090
rect 15538 15038 15540 15090
rect 15484 14980 15540 15038
rect 15484 14914 15540 14924
rect 15708 15092 15876 15148
rect 15708 15090 15764 15092
rect 15708 15038 15710 15090
rect 15762 15038 15764 15090
rect 15036 14476 15204 14532
rect 15036 14308 15092 14318
rect 15036 14214 15092 14252
rect 14512 13356 14776 13366
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14512 13290 14776 13300
rect 14588 13188 14644 13198
rect 14924 13188 14980 13356
rect 15036 13188 15092 13198
rect 14924 13186 15092 13188
rect 14924 13134 15038 13186
rect 15090 13134 15092 13186
rect 14924 13132 15092 13134
rect 14588 13094 14644 13132
rect 15036 13122 15092 13132
rect 14812 12964 14868 12974
rect 15148 12964 15204 14476
rect 15372 14466 15428 14476
rect 15708 14308 15764 15038
rect 15820 15026 15876 15036
rect 15708 14242 15764 14252
rect 15372 13188 15428 13198
rect 15596 13188 15652 13198
rect 15932 13188 15988 16044
rect 16044 14980 16100 18396
rect 16268 18450 16324 18462
rect 16268 18398 16270 18450
rect 16322 18398 16324 18450
rect 16268 18340 16324 18398
rect 16268 15148 16324 18284
rect 16604 18228 16660 18510
rect 16604 18162 16660 18172
rect 18284 18450 18340 18462
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 17172 17276 17436 17286
rect 17228 17220 17276 17276
rect 17332 17220 17380 17276
rect 17172 17210 17436 17220
rect 17172 15708 17436 15718
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17172 15642 17436 15652
rect 18172 15428 18228 15438
rect 18284 15428 18340 18398
rect 19516 18228 19572 18238
rect 19516 17780 19572 18172
rect 19832 18060 20096 18070
rect 19888 18004 19936 18060
rect 19992 18004 20040 18060
rect 19832 17994 20096 18004
rect 19852 17892 19908 17902
rect 19516 17686 19572 17724
rect 19628 17836 19852 17892
rect 19628 17108 19684 17836
rect 19852 17798 19908 17836
rect 20636 17892 20692 19180
rect 19964 17780 20020 17790
rect 19964 17686 20020 17724
rect 19516 17052 19684 17108
rect 20188 17666 20244 17678
rect 20188 17614 20190 17666
rect 20242 17614 20244 17666
rect 19404 16884 19460 16922
rect 19404 16818 19460 16828
rect 19404 16324 19460 16334
rect 19516 16324 19572 17052
rect 19628 16884 19684 16894
rect 19964 16884 20020 16894
rect 19628 16882 20020 16884
rect 19628 16830 19630 16882
rect 19682 16830 19966 16882
rect 20018 16830 20020 16882
rect 19628 16828 20020 16830
rect 19628 16818 19684 16828
rect 19740 16660 19796 16698
rect 19964 16660 20020 16828
rect 20188 16884 20244 17614
rect 20300 17666 20356 17678
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20300 17106 20356 17614
rect 20300 17054 20302 17106
rect 20354 17054 20356 17106
rect 20300 17042 20356 17054
rect 20524 16996 20580 17006
rect 20188 16818 20244 16828
rect 20412 16940 20524 16996
rect 20412 16882 20468 16940
rect 20524 16930 20580 16940
rect 20636 16994 20692 17836
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16930 20692 16942
rect 20412 16830 20414 16882
rect 20466 16830 20468 16882
rect 20412 16818 20468 16830
rect 20300 16660 20356 16670
rect 19964 16604 20244 16660
rect 19740 16594 19796 16604
rect 19832 16492 20096 16502
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 19832 16426 20096 16436
rect 19404 16322 19572 16324
rect 19404 16270 19406 16322
rect 19458 16270 19572 16322
rect 19404 16268 19572 16270
rect 19404 16258 19460 16268
rect 19180 16100 19236 16110
rect 19180 16006 19236 16044
rect 19516 15876 19572 16268
rect 19740 16324 19796 16334
rect 20188 16324 20244 16604
rect 19740 16230 19796 16268
rect 20076 16268 20244 16324
rect 19628 16212 19684 16222
rect 19628 16118 19684 16156
rect 20076 16098 20132 16268
rect 20076 16046 20078 16098
rect 20130 16046 20132 16098
rect 20076 16034 20132 16046
rect 19516 15820 19684 15876
rect 18172 15426 18340 15428
rect 18172 15374 18174 15426
rect 18226 15374 18340 15426
rect 18172 15372 18340 15374
rect 18172 15362 18228 15372
rect 18844 15316 18900 15326
rect 17500 15202 17556 15214
rect 17500 15150 17502 15202
rect 17554 15150 17556 15202
rect 16268 15092 16436 15148
rect 16044 14914 16100 14924
rect 16268 13188 16324 13198
rect 15428 13132 15540 13188
rect 15372 13122 15428 13132
rect 14812 12962 15204 12964
rect 14812 12910 14814 12962
rect 14866 12910 15204 12962
rect 14812 12908 15204 12910
rect 15260 12962 15316 12974
rect 15260 12910 15262 12962
rect 15314 12910 15316 12962
rect 14812 12898 14868 12908
rect 14476 12852 14532 12862
rect 14476 12758 14532 12796
rect 14512 11788 14776 11798
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14512 11722 14776 11732
rect 14924 11732 14980 12908
rect 15148 12740 15204 12750
rect 15260 12740 15316 12910
rect 15484 12964 15540 13132
rect 15596 13186 15988 13188
rect 15596 13134 15598 13186
rect 15650 13134 15988 13186
rect 15596 13132 15988 13134
rect 16044 13186 16324 13188
rect 16044 13134 16270 13186
rect 16322 13134 16324 13186
rect 16044 13132 16324 13134
rect 15596 13122 15652 13132
rect 15708 12964 15764 12974
rect 15484 12962 15764 12964
rect 15484 12910 15710 12962
rect 15762 12910 15764 12962
rect 15484 12908 15764 12910
rect 15708 12898 15764 12908
rect 15932 12964 15988 12974
rect 15932 12870 15988 12908
rect 16044 12740 16100 13132
rect 16268 13122 16324 13132
rect 15260 12684 16100 12740
rect 16156 12962 16212 12974
rect 16156 12910 16158 12962
rect 16210 12910 16212 12962
rect 15148 11844 15204 12684
rect 15372 12292 15428 12302
rect 14924 11666 14980 11676
rect 15036 11788 15204 11844
rect 15260 12180 15316 12190
rect 14700 11620 14756 11630
rect 14364 11618 14756 11620
rect 14364 11566 14702 11618
rect 14754 11566 14756 11618
rect 14364 11564 14756 11566
rect 13916 11554 13972 11564
rect 14700 11554 14756 11564
rect 15036 11618 15092 11788
rect 15036 11566 15038 11618
rect 15090 11566 15092 11618
rect 15036 11554 15092 11566
rect 12460 11394 12516 11406
rect 12460 11342 12462 11394
rect 12514 11342 12516 11394
rect 11852 11004 12116 11014
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 11852 10938 12116 10948
rect 12460 10836 12516 11342
rect 13692 11394 13748 11452
rect 13692 11342 13694 11394
rect 13746 11342 13748 11394
rect 13692 11330 13748 11342
rect 14252 11394 14308 11406
rect 14252 11342 14254 11394
rect 14306 11342 14308 11394
rect 13468 11284 13524 11294
rect 13468 11190 13524 11228
rect 14252 11284 14308 11342
rect 14924 11394 14980 11406
rect 14924 11342 14926 11394
rect 14978 11342 14980 11394
rect 14588 11284 14644 11294
rect 12460 10770 12516 10780
rect 12572 11170 12628 11182
rect 12572 11118 12574 11170
rect 12626 11118 12628 11170
rect 12572 10164 12628 11118
rect 13580 11172 13636 11182
rect 13580 11078 13636 11116
rect 14252 10834 14308 11228
rect 14252 10782 14254 10834
rect 14306 10782 14308 10834
rect 14252 10770 14308 10782
rect 14364 11282 14644 11284
rect 14364 11230 14590 11282
rect 14642 11230 14644 11282
rect 14364 11228 14644 11230
rect 12572 10098 12628 10108
rect 11852 9436 12116 9446
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 11852 9370 12116 9380
rect 14252 8820 14308 8830
rect 11564 8260 11620 8270
rect 11564 8166 11620 8204
rect 14252 8034 14308 8764
rect 14364 8484 14420 11228
rect 14588 11218 14644 11228
rect 14924 11284 14980 11342
rect 14924 11218 14980 11228
rect 15036 11060 15092 11070
rect 14476 10836 14532 10846
rect 14476 10610 14532 10780
rect 14476 10558 14478 10610
rect 14530 10558 14532 10610
rect 14476 10546 14532 10558
rect 15036 10610 15092 11004
rect 15260 11060 15316 12124
rect 15260 10994 15316 11004
rect 15372 10836 15428 12236
rect 15484 11508 15540 11518
rect 15484 11282 15540 11452
rect 15820 11508 15876 11518
rect 15820 11394 15876 11452
rect 15820 11342 15822 11394
rect 15874 11342 15876 11394
rect 15820 11330 15876 11342
rect 15484 11230 15486 11282
rect 15538 11230 15540 11282
rect 15484 11218 15540 11230
rect 15036 10558 15038 10610
rect 15090 10558 15092 10610
rect 15036 10546 15092 10558
rect 15260 10780 15428 10836
rect 15260 10610 15316 10780
rect 15260 10558 15262 10610
rect 15314 10558 15316 10610
rect 15260 10546 15316 10558
rect 15596 10610 15652 10622
rect 15596 10558 15598 10610
rect 15650 10558 15652 10610
rect 15372 10498 15428 10510
rect 15372 10446 15374 10498
rect 15426 10446 15428 10498
rect 15260 10388 15316 10398
rect 15372 10388 15428 10446
rect 15316 10332 15428 10388
rect 15260 10322 15316 10332
rect 14512 10220 14776 10230
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14512 10154 14776 10164
rect 15596 9828 15652 10558
rect 15596 9762 15652 9772
rect 14512 8652 14776 8662
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14512 8586 14776 8596
rect 15932 8428 15988 12684
rect 16156 12180 16212 12910
rect 16156 12114 16212 12124
rect 16268 12292 16324 12302
rect 16156 11732 16212 11742
rect 16156 11282 16212 11676
rect 16156 11230 16158 11282
rect 16210 11230 16212 11282
rect 16156 11218 16212 11230
rect 14364 8418 14420 8428
rect 15036 8372 15988 8428
rect 15036 8370 15092 8372
rect 15036 8318 15038 8370
rect 15090 8318 15092 8370
rect 15036 8306 15092 8318
rect 15148 8258 15204 8270
rect 15372 8260 15428 8270
rect 15148 8206 15150 8258
rect 15202 8206 15204 8258
rect 14252 7982 14254 8034
rect 14306 7982 14308 8034
rect 11852 7868 12116 7878
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 11852 7802 12116 7812
rect 11004 6414 11006 6466
rect 11058 6414 11060 6466
rect 11004 6402 11060 6414
rect 11228 7196 11508 7252
rect 11788 7700 11844 7710
rect 14252 7700 14308 7982
rect 14588 8036 14644 8046
rect 14588 7942 14644 7980
rect 15148 7924 15204 8206
rect 15148 7858 15204 7868
rect 15260 8204 15372 8260
rect 14924 7700 14980 7710
rect 14252 7698 14980 7700
rect 14252 7646 14926 7698
rect 14978 7646 14980 7698
rect 14252 7644 14980 7646
rect 11004 6132 11060 6142
rect 10444 6130 11060 6132
rect 10444 6078 11006 6130
rect 11058 6078 11060 6130
rect 10444 6076 11060 6078
rect 11004 6066 11060 6076
rect 9884 6020 9940 6030
rect 9660 5964 9884 6020
rect 9884 5926 9940 5964
rect 10332 6020 10388 6030
rect 10332 5926 10388 5964
rect 11228 6020 11284 7196
rect 11452 6692 11508 6702
rect 11452 6598 11508 6636
rect 11788 6578 11844 7644
rect 14924 7634 14980 7644
rect 15260 7698 15316 8204
rect 15372 8166 15428 8204
rect 15484 8258 15540 8270
rect 15484 8206 15486 8258
rect 15538 8206 15540 8258
rect 15484 8148 15540 8206
rect 15932 8258 15988 8372
rect 15932 8206 15934 8258
rect 15986 8206 15988 8258
rect 15932 8194 15988 8206
rect 16268 8260 16324 12236
rect 16268 8194 16324 8204
rect 15540 8092 15764 8148
rect 15484 8082 15540 8092
rect 15260 7646 15262 7698
rect 15314 7646 15316 7698
rect 15260 7634 15316 7646
rect 15708 7476 15764 8092
rect 16268 8036 16324 8046
rect 16268 7942 16324 7980
rect 16380 7924 16436 15092
rect 16940 14980 16996 14990
rect 16996 14924 17108 14980
rect 16940 14914 16996 14924
rect 17052 12404 17108 14924
rect 17172 14140 17436 14150
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17172 14074 17436 14084
rect 17500 13412 17556 15150
rect 17612 15204 17668 15214
rect 17612 15110 17668 15148
rect 17836 15204 17892 15214
rect 18060 15204 18116 15214
rect 17500 13346 17556 13356
rect 17172 12572 17436 12582
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17172 12506 17436 12516
rect 17052 12348 17220 12404
rect 17164 12180 17220 12348
rect 17052 11620 17108 11630
rect 17052 11526 17108 11564
rect 17164 11618 17220 12124
rect 17164 11566 17166 11618
rect 17218 11566 17220 11618
rect 17164 11554 17220 11566
rect 17388 11732 17444 11742
rect 17388 11618 17444 11676
rect 17388 11566 17390 11618
rect 17442 11566 17444 11618
rect 17388 11554 17444 11566
rect 17612 11396 17668 11406
rect 17612 11302 17668 11340
rect 16492 11284 16548 11294
rect 16492 11190 16548 11228
rect 17172 11004 17436 11014
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17172 10938 17436 10948
rect 17172 9436 17436 9446
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17172 9370 17436 9380
rect 17836 8372 17892 15148
rect 17948 15202 18116 15204
rect 17948 15150 18062 15202
rect 18114 15150 18116 15202
rect 17948 15148 18116 15150
rect 17948 15092 18004 15148
rect 18060 15138 18116 15148
rect 17948 13074 18004 15036
rect 17948 13022 17950 13074
rect 18002 13022 18004 13074
rect 17948 13010 18004 13022
rect 18284 13412 18340 13422
rect 18172 12962 18228 12974
rect 18172 12910 18174 12962
rect 18226 12910 18228 12962
rect 18060 12180 18116 12190
rect 18060 12086 18116 12124
rect 17948 11954 18004 11966
rect 17948 11902 17950 11954
rect 18002 11902 18004 11954
rect 17948 11508 18004 11902
rect 17948 11396 18004 11452
rect 18060 11396 18116 11406
rect 17948 11394 18116 11396
rect 17948 11342 18062 11394
rect 18114 11342 18116 11394
rect 17948 11340 18116 11342
rect 18060 11330 18116 11340
rect 18172 11284 18228 12910
rect 18284 12852 18340 13356
rect 18844 13186 18900 15260
rect 19180 15314 19236 15326
rect 19180 15262 19182 15314
rect 19234 15262 19236 15314
rect 19180 13972 19236 15262
rect 19516 15316 19572 15326
rect 19516 15222 19572 15260
rect 19628 15314 19684 15820
rect 20300 15874 20356 16604
rect 20300 15822 20302 15874
rect 20354 15822 20356 15874
rect 20300 15810 20356 15822
rect 20412 15986 20468 15998
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 19964 15540 20020 15550
rect 19964 15446 20020 15484
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19628 15250 19684 15262
rect 19740 15428 19796 15438
rect 19740 15314 19796 15372
rect 19740 15262 19742 15314
rect 19794 15262 19796 15314
rect 19740 15204 19796 15262
rect 20300 15316 20356 15326
rect 20300 15222 20356 15260
rect 19740 15138 19796 15148
rect 19832 14924 20096 14934
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 19832 14858 20096 14868
rect 19180 13906 19236 13916
rect 19832 13356 20096 13366
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 19832 13290 20096 13300
rect 18844 13134 18846 13186
rect 18898 13134 18900 13186
rect 18844 13122 18900 13134
rect 18396 12964 18452 12974
rect 19404 12964 19460 12974
rect 18452 12908 18564 12964
rect 18396 12870 18452 12908
rect 18284 12178 18340 12796
rect 18284 12126 18286 12178
rect 18338 12126 18340 12178
rect 18284 12114 18340 12126
rect 18508 12180 18564 12908
rect 19292 12908 19404 12964
rect 19068 12852 19124 12862
rect 19068 12758 19124 12796
rect 19292 12292 19348 12908
rect 19404 12898 19460 12908
rect 20412 12964 20468 15934
rect 20636 15986 20692 15998
rect 20636 15934 20638 15986
rect 20690 15934 20692 15986
rect 20636 15540 20692 15934
rect 20860 15652 20916 19964
rect 20972 19954 21028 19964
rect 21644 20018 21924 20020
rect 21644 19966 21870 20018
rect 21922 19966 21924 20018
rect 21644 19964 21924 19966
rect 21644 19236 21700 19964
rect 21868 19954 21924 19964
rect 21644 19142 21700 19180
rect 22204 19124 22260 19134
rect 21308 19012 21364 19022
rect 21364 18956 21588 19012
rect 21308 18918 21364 18956
rect 20972 16882 21028 16894
rect 20972 16830 20974 16882
rect 21026 16830 21028 16882
rect 20972 16660 21028 16830
rect 21196 16884 21252 16894
rect 20972 16594 21028 16604
rect 21084 16770 21140 16782
rect 21084 16718 21086 16770
rect 21138 16718 21140 16770
rect 21084 16100 21140 16718
rect 21196 16324 21252 16828
rect 21308 16324 21364 16334
rect 21196 16322 21364 16324
rect 21196 16270 21310 16322
rect 21362 16270 21364 16322
rect 21196 16268 21364 16270
rect 21308 16258 21364 16268
rect 21420 16100 21476 16110
rect 21084 16098 21476 16100
rect 21084 16046 21422 16098
rect 21474 16046 21476 16098
rect 21084 16044 21476 16046
rect 21420 16034 21476 16044
rect 20860 15586 20916 15596
rect 20636 15474 20692 15484
rect 20524 15428 20580 15438
rect 20524 15334 20580 15372
rect 20636 15316 20692 15326
rect 20636 15202 20692 15260
rect 20636 15150 20638 15202
rect 20690 15150 20692 15202
rect 20636 15138 20692 15150
rect 20412 12898 20468 12908
rect 20748 12852 20804 12862
rect 20748 12758 20804 12796
rect 21420 12852 21476 12862
rect 19292 12198 19348 12236
rect 19404 12738 19460 12750
rect 19404 12686 19406 12738
rect 19458 12686 19460 12738
rect 19404 12402 19460 12686
rect 20636 12738 20692 12750
rect 20636 12686 20638 12738
rect 20690 12686 20692 12738
rect 20636 12516 20692 12686
rect 21420 12628 21476 12796
rect 21532 12740 21588 18956
rect 21868 18562 21924 18574
rect 21868 18510 21870 18562
rect 21922 18510 21924 18562
rect 21644 18452 21700 18462
rect 21644 18358 21700 18396
rect 21868 17444 21924 18510
rect 22204 18452 22260 19068
rect 22492 18844 22756 18854
rect 22548 18788 22596 18844
rect 22652 18788 22700 18844
rect 22492 18778 22756 18788
rect 22204 18358 22260 18396
rect 21868 17388 22932 17444
rect 22492 17276 22756 17286
rect 22548 17220 22596 17276
rect 22652 17220 22700 17276
rect 22492 17210 22756 17220
rect 21644 16996 21700 17006
rect 21644 16884 21700 16940
rect 21868 16994 21924 17006
rect 21868 16942 21870 16994
rect 21922 16942 21924 16994
rect 21644 16882 21812 16884
rect 21644 16830 21646 16882
rect 21698 16830 21812 16882
rect 21644 16828 21812 16830
rect 21644 16818 21700 16828
rect 21644 13636 21700 13646
rect 21644 13542 21700 13580
rect 21756 13076 21812 16828
rect 21868 16212 21924 16942
rect 22204 16882 22260 16894
rect 22204 16830 22206 16882
rect 22258 16830 22260 16882
rect 22204 16212 22260 16830
rect 22316 16212 22372 16222
rect 22204 16156 22316 16212
rect 21868 16146 21924 16156
rect 22316 16118 22372 16156
rect 22492 15708 22756 15718
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22492 15642 22756 15652
rect 22492 14140 22756 14150
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22492 14074 22756 14084
rect 21868 13860 21924 13870
rect 21868 13858 22036 13860
rect 21868 13806 21870 13858
rect 21922 13806 22036 13858
rect 21868 13804 22036 13806
rect 21868 13794 21924 13804
rect 21756 13020 21924 13076
rect 21532 12684 21700 12740
rect 21420 12572 21588 12628
rect 19404 12350 19406 12402
rect 19458 12350 19460 12402
rect 18396 11956 18452 11966
rect 18396 11862 18452 11900
rect 18508 11732 18564 12124
rect 19180 12180 19236 12190
rect 19180 12086 19236 12124
rect 18172 11218 18228 11228
rect 18396 11676 18564 11732
rect 18396 11282 18452 11676
rect 18396 11230 18398 11282
rect 18450 11230 18452 11282
rect 18396 11218 18452 11230
rect 19404 11172 19460 12350
rect 20412 12460 20692 12516
rect 21084 12516 21140 12526
rect 20412 12292 20468 12460
rect 20748 12404 20804 12414
rect 21084 12404 21140 12460
rect 19628 12180 19684 12190
rect 19628 12086 19684 12124
rect 20300 12180 20356 12190
rect 19832 11788 20096 11798
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 19832 11722 20096 11732
rect 20300 11618 20356 12124
rect 20300 11566 20302 11618
rect 20354 11566 20356 11618
rect 20300 11554 20356 11566
rect 20412 11956 20468 12236
rect 20636 12348 20748 12404
rect 19404 11106 19460 11116
rect 19852 11396 19908 11406
rect 19852 10836 19908 11340
rect 20412 11282 20468 11900
rect 20412 11230 20414 11282
rect 20466 11230 20468 11282
rect 20412 11218 20468 11230
rect 20524 12178 20580 12190
rect 20524 12126 20526 12178
rect 20578 12126 20580 12178
rect 19404 10834 19908 10836
rect 19404 10782 19854 10834
rect 19906 10782 19908 10834
rect 19404 10780 19908 10782
rect 19180 9940 19236 9950
rect 19180 9716 19236 9884
rect 19404 9826 19460 10780
rect 19852 10770 19908 10780
rect 19964 10612 20020 10622
rect 19516 10610 20020 10612
rect 19516 10558 19966 10610
rect 20018 10558 20020 10610
rect 19516 10556 20020 10558
rect 19516 9938 19572 10556
rect 19964 10546 20020 10556
rect 20524 10276 20580 12126
rect 20636 11618 20692 12348
rect 20748 12310 20804 12348
rect 20972 12348 21140 12404
rect 21196 12404 21252 12414
rect 21420 12404 21476 12414
rect 21252 12402 21476 12404
rect 21252 12350 21422 12402
rect 21474 12350 21476 12402
rect 21252 12348 21476 12350
rect 20636 11566 20638 11618
rect 20690 11566 20692 11618
rect 20636 11554 20692 11566
rect 20748 12180 20804 12190
rect 20972 12180 21028 12348
rect 21196 12338 21252 12348
rect 21420 12338 21476 12348
rect 21532 12402 21588 12572
rect 21644 12516 21700 12684
rect 21644 12450 21700 12460
rect 21532 12350 21534 12402
rect 21586 12350 21588 12402
rect 21532 12338 21588 12350
rect 21868 12402 21924 13020
rect 21868 12350 21870 12402
rect 21922 12350 21924 12402
rect 21644 12292 21700 12302
rect 21644 12198 21700 12236
rect 20748 12178 21028 12180
rect 20748 12126 20750 12178
rect 20802 12126 21028 12178
rect 20748 12124 21028 12126
rect 21084 12180 21140 12190
rect 19832 10220 20096 10230
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 19832 10154 20096 10164
rect 20188 10220 20580 10276
rect 19516 9886 19518 9938
rect 19570 9886 19572 9938
rect 19516 9874 19572 9886
rect 20188 9940 20244 10220
rect 20748 10164 20804 12124
rect 21084 12086 21140 12124
rect 21868 11844 21924 12350
rect 21980 12180 22036 13804
rect 22204 13746 22260 13758
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 22204 13636 22260 13694
rect 22204 13300 22260 13580
rect 22204 13234 22260 13244
rect 22492 12572 22756 12582
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22492 12506 22756 12516
rect 21980 12114 22036 12124
rect 21532 11788 21924 11844
rect 20972 10724 21028 10734
rect 20524 10108 20804 10164
rect 20860 10668 20972 10724
rect 20524 10052 20580 10108
rect 19964 9828 20020 9838
rect 19404 9774 19406 9826
rect 19458 9774 19460 9826
rect 19180 9714 19348 9716
rect 19180 9662 19182 9714
rect 19234 9662 19348 9714
rect 19180 9660 19348 9662
rect 19180 9650 19236 9660
rect 17836 8306 17892 8316
rect 16604 8260 16660 8270
rect 16604 8166 16660 8204
rect 18060 8148 18116 8158
rect 16380 7858 16436 7868
rect 17172 7868 17436 7878
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17172 7802 17436 7812
rect 18060 7698 18116 8092
rect 18060 7646 18062 7698
rect 18114 7646 18116 7698
rect 18060 7634 18116 7646
rect 18284 8148 18340 8158
rect 14512 7084 14776 7094
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14512 7018 14776 7028
rect 11788 6526 11790 6578
rect 11842 6526 11844 6578
rect 11788 6514 11844 6526
rect 15708 6578 15764 7420
rect 18284 7474 18340 8092
rect 19068 8148 19124 8158
rect 19292 8148 19348 9660
rect 19404 9044 19460 9774
rect 19852 9772 19964 9828
rect 19628 9716 19684 9726
rect 19628 9622 19684 9660
rect 19852 9266 19908 9772
rect 19964 9734 20020 9772
rect 20188 9826 20244 9884
rect 20188 9774 20190 9826
rect 20242 9774 20244 9826
rect 19852 9214 19854 9266
rect 19906 9214 19908 9266
rect 19852 9202 19908 9214
rect 20076 9716 20132 9726
rect 19964 9156 20020 9166
rect 20076 9156 20132 9660
rect 19964 9154 20132 9156
rect 19964 9102 19966 9154
rect 20018 9102 20132 9154
rect 19964 9100 20132 9102
rect 19964 9090 20020 9100
rect 19628 9044 19684 9054
rect 19404 9042 19684 9044
rect 19404 8990 19630 9042
rect 19682 8990 19684 9042
rect 19404 8988 19684 8990
rect 19628 8978 19684 8988
rect 19832 8652 20096 8662
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 19832 8586 20096 8596
rect 20188 8484 20244 9774
rect 20076 8428 20244 8484
rect 20300 10050 20580 10052
rect 20300 9998 20526 10050
rect 20578 9998 20580 10050
rect 20300 9996 20580 9998
rect 20300 8482 20356 9996
rect 20524 9986 20580 9996
rect 20748 9828 20804 9838
rect 20860 9828 20916 10668
rect 20972 10658 21028 10668
rect 20748 9826 20916 9828
rect 20748 9774 20750 9826
rect 20802 9774 20916 9826
rect 20748 9772 20916 9774
rect 20748 9762 20804 9772
rect 20300 8430 20302 8482
rect 20354 8430 20356 8482
rect 19740 8260 19796 8270
rect 19404 8148 19460 8158
rect 19292 8146 19460 8148
rect 19292 8094 19406 8146
rect 19458 8094 19460 8146
rect 19292 8092 19460 8094
rect 19068 8054 19124 8092
rect 19404 8082 19460 8092
rect 19404 7700 19460 7710
rect 19404 7606 19460 7644
rect 18956 7588 19012 7598
rect 18956 7494 19012 7532
rect 18284 7422 18286 7474
rect 18338 7422 18340 7474
rect 17948 7364 18004 7374
rect 17948 6690 18004 7308
rect 17948 6638 17950 6690
rect 18002 6638 18004 6690
rect 17948 6626 18004 6638
rect 15708 6526 15710 6578
rect 15762 6526 15764 6578
rect 15708 6514 15764 6526
rect 17724 6580 17780 6590
rect 11340 6468 11396 6478
rect 11340 6130 11396 6412
rect 16044 6468 16100 6478
rect 16044 6374 16100 6412
rect 11852 6300 12116 6310
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 11852 6234 12116 6244
rect 17172 6300 17436 6310
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17172 6234 17436 6244
rect 11340 6078 11342 6130
rect 11394 6078 11396 6130
rect 11340 6066 11396 6078
rect 17724 6130 17780 6524
rect 18284 6580 18340 7422
rect 19180 7476 19236 7486
rect 19180 7382 19236 7420
rect 19068 7364 19124 7374
rect 19740 7364 19796 8204
rect 20076 8258 20132 8428
rect 20300 8418 20356 8430
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 20076 8194 20132 8206
rect 20524 8260 20580 8270
rect 20524 8166 20580 8204
rect 21420 8148 21476 8158
rect 21420 8054 21476 8092
rect 20188 8034 20244 8046
rect 20188 7982 20190 8034
rect 20242 7982 20244 8034
rect 19964 7586 20020 7598
rect 19964 7534 19966 7586
rect 20018 7534 20020 7586
rect 19964 7476 20020 7534
rect 20188 7588 20244 7982
rect 21308 8036 21364 8046
rect 21308 7942 21364 7980
rect 21532 7812 21588 11788
rect 22492 11004 22756 11014
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22492 10938 22756 10948
rect 21868 10724 21924 10734
rect 21868 10630 21924 10668
rect 22204 10610 22260 10622
rect 22204 10558 22206 10610
rect 22258 10558 22260 10610
rect 21644 10498 21700 10510
rect 21644 10446 21646 10498
rect 21698 10446 21700 10498
rect 21644 10388 21700 10446
rect 21644 10322 21700 10332
rect 22204 10388 22260 10558
rect 22204 10322 22260 10332
rect 22492 9436 22756 9446
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22492 9370 22756 9380
rect 22876 8260 22932 17388
rect 22876 8194 22932 8204
rect 21868 8148 21924 8158
rect 21868 8054 21924 8092
rect 22204 8146 22260 8158
rect 22204 8094 22206 8146
rect 22258 8094 22260 8146
rect 20188 7494 20244 7532
rect 21308 7756 21588 7812
rect 21308 7700 21364 7756
rect 19964 7410 20020 7420
rect 19852 7364 19908 7374
rect 19740 7362 19908 7364
rect 19740 7310 19854 7362
rect 19906 7310 19908 7362
rect 19740 7308 19908 7310
rect 19068 7270 19124 7308
rect 19852 7298 19908 7308
rect 19832 7084 20096 7094
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 19832 7018 20096 7028
rect 18284 6514 18340 6524
rect 21308 6578 21364 7644
rect 22204 7476 22260 8094
rect 22492 7868 22756 7878
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22492 7802 22756 7812
rect 22204 7382 22260 7420
rect 21308 6526 21310 6578
rect 21362 6526 21364 6578
rect 21308 6514 21364 6526
rect 21532 6690 21588 6702
rect 21532 6638 21534 6690
rect 21586 6638 21588 6690
rect 17836 6468 17892 6478
rect 17836 6374 17892 6412
rect 21532 6468 21588 6638
rect 22092 6468 22148 6478
rect 21532 6466 22148 6468
rect 21532 6414 22094 6466
rect 22146 6414 22148 6466
rect 21532 6412 22148 6414
rect 17724 6078 17726 6130
rect 17778 6078 17780 6130
rect 17724 6066 17780 6078
rect 17948 6132 18004 6142
rect 11228 5954 11284 5964
rect 17948 5906 18004 6076
rect 18508 6132 18564 6142
rect 18508 6038 18564 6076
rect 21532 6132 21588 6412
rect 21532 6066 21588 6076
rect 17948 5854 17950 5906
rect 18002 5854 18004 5906
rect 17948 5842 18004 5854
rect 21868 6020 21924 6030
rect 3872 5516 4136 5526
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 3872 5450 4136 5460
rect 9192 5516 9456 5526
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9192 5450 9456 5460
rect 14512 5516 14776 5526
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14512 5450 14776 5460
rect 19832 5516 20096 5526
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 19832 5450 20096 5460
rect 21644 5124 21700 5134
rect 21644 5030 21700 5068
rect 21868 5010 21924 5964
rect 21868 4958 21870 5010
rect 21922 4958 21924 5010
rect 21868 4946 21924 4958
rect 6532 4732 6796 4742
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6532 4666 6796 4676
rect 11852 4732 12116 4742
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 11852 4666 12116 4676
rect 17172 4732 17436 4742
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17172 4666 17436 4676
rect 3872 3948 4136 3958
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 3872 3882 4136 3892
rect 9192 3948 9456 3958
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9192 3882 9456 3892
rect 14512 3948 14776 3958
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14512 3882 14776 3892
rect 19832 3948 20096 3958
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 19832 3882 20096 3892
rect 6532 3164 6796 3174
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6532 3098 6796 3108
rect 11852 3164 12116 3174
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 11852 3098 12116 3108
rect 17172 3164 17436 3174
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17172 3098 17436 3108
rect 22092 1652 22148 6412
rect 22492 6300 22756 6310
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22492 6234 22756 6244
rect 22204 5124 22260 5134
rect 22204 4564 22260 5068
rect 22492 4732 22756 4742
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22492 4666 22756 4676
rect 22204 4498 22260 4508
rect 22492 3164 22756 3174
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22492 3098 22756 3108
rect 22092 1586 22148 1596
<< via2 >>
rect 6532 20410 6588 20412
rect 6532 20358 6534 20410
rect 6534 20358 6586 20410
rect 6586 20358 6588 20410
rect 6532 20356 6588 20358
rect 6636 20410 6692 20412
rect 6636 20358 6638 20410
rect 6638 20358 6690 20410
rect 6690 20358 6692 20410
rect 6636 20356 6692 20358
rect 6740 20410 6796 20412
rect 6740 20358 6742 20410
rect 6742 20358 6794 20410
rect 6794 20358 6796 20410
rect 6740 20356 6796 20358
rect 11852 20410 11908 20412
rect 11852 20358 11854 20410
rect 11854 20358 11906 20410
rect 11906 20358 11908 20410
rect 11852 20356 11908 20358
rect 11956 20410 12012 20412
rect 11956 20358 11958 20410
rect 11958 20358 12010 20410
rect 12010 20358 12012 20410
rect 11956 20356 12012 20358
rect 12060 20410 12116 20412
rect 12060 20358 12062 20410
rect 12062 20358 12114 20410
rect 12114 20358 12116 20410
rect 12060 20356 12116 20358
rect 17172 20410 17228 20412
rect 17172 20358 17174 20410
rect 17174 20358 17226 20410
rect 17226 20358 17228 20410
rect 17172 20356 17228 20358
rect 17276 20410 17332 20412
rect 17276 20358 17278 20410
rect 17278 20358 17330 20410
rect 17330 20358 17332 20410
rect 17276 20356 17332 20358
rect 17380 20410 17436 20412
rect 17380 20358 17382 20410
rect 17382 20358 17434 20410
rect 17434 20358 17436 20410
rect 17380 20356 17436 20358
rect 19740 20076 19796 20132
rect 20076 21980 20132 22036
rect 22492 20410 22548 20412
rect 22492 20358 22494 20410
rect 22494 20358 22546 20410
rect 22546 20358 22548 20410
rect 22492 20356 22548 20358
rect 22596 20410 22652 20412
rect 22596 20358 22598 20410
rect 22598 20358 22650 20410
rect 22650 20358 22652 20410
rect 22596 20356 22652 20358
rect 22700 20410 22756 20412
rect 22700 20358 22702 20410
rect 22702 20358 22754 20410
rect 22754 20358 22756 20410
rect 22700 20356 22756 20358
rect 20748 20130 20804 20132
rect 20748 20078 20750 20130
rect 20750 20078 20802 20130
rect 20802 20078 20804 20130
rect 20748 20076 20804 20078
rect 3872 19626 3928 19628
rect 3872 19574 3874 19626
rect 3874 19574 3926 19626
rect 3926 19574 3928 19626
rect 3872 19572 3928 19574
rect 3976 19626 4032 19628
rect 3976 19574 3978 19626
rect 3978 19574 4030 19626
rect 4030 19574 4032 19626
rect 3976 19572 4032 19574
rect 4080 19626 4136 19628
rect 4080 19574 4082 19626
rect 4082 19574 4134 19626
rect 4134 19574 4136 19626
rect 4080 19572 4136 19574
rect 3052 19234 3108 19236
rect 3052 19182 3054 19234
rect 3054 19182 3106 19234
rect 3106 19182 3108 19234
rect 3052 19180 3108 19182
rect 3164 18508 3220 18564
rect 4172 19180 4228 19236
rect 3052 17836 3108 17892
rect 3388 18172 3444 18228
rect 3836 18562 3892 18564
rect 3836 18510 3838 18562
rect 3838 18510 3890 18562
rect 3890 18510 3892 18562
rect 3836 18508 3892 18510
rect 4620 19122 4676 19124
rect 4620 19070 4622 19122
rect 4622 19070 4674 19122
rect 4674 19070 4676 19122
rect 4620 19068 4676 19070
rect 3872 18058 3928 18060
rect 3872 18006 3874 18058
rect 3874 18006 3926 18058
rect 3926 18006 3928 18058
rect 3872 18004 3928 18006
rect 3976 18058 4032 18060
rect 3976 18006 3978 18058
rect 3978 18006 4030 18058
rect 4030 18006 4032 18058
rect 3976 18004 4032 18006
rect 4080 18058 4136 18060
rect 4080 18006 4082 18058
rect 4082 18006 4134 18058
rect 4134 18006 4136 18058
rect 4080 18004 4136 18006
rect 3500 17666 3556 17668
rect 3500 17614 3502 17666
rect 3502 17614 3554 17666
rect 3554 17614 3556 17666
rect 3500 17612 3556 17614
rect 3164 17388 3220 17444
rect 2940 16044 2996 16100
rect 2380 13692 2436 13748
rect 3052 14140 3108 14196
rect 3052 13746 3108 13748
rect 3052 13694 3054 13746
rect 3054 13694 3106 13746
rect 3106 13694 3108 13746
rect 3052 13692 3108 13694
rect 3612 14530 3668 14532
rect 3612 14478 3614 14530
rect 3614 14478 3666 14530
rect 3666 14478 3668 14530
rect 3612 14476 3668 14478
rect 3872 16490 3928 16492
rect 3872 16438 3874 16490
rect 3874 16438 3926 16490
rect 3926 16438 3928 16490
rect 3872 16436 3928 16438
rect 3976 16490 4032 16492
rect 3976 16438 3978 16490
rect 3978 16438 4030 16490
rect 4030 16438 4032 16490
rect 3976 16436 4032 16438
rect 4080 16490 4136 16492
rect 4080 16438 4082 16490
rect 4082 16438 4134 16490
rect 4134 16438 4136 16490
rect 4080 16436 4136 16438
rect 3872 14922 3928 14924
rect 3872 14870 3874 14922
rect 3874 14870 3926 14922
rect 3926 14870 3928 14922
rect 3872 14868 3928 14870
rect 3976 14922 4032 14924
rect 3976 14870 3978 14922
rect 3978 14870 4030 14922
rect 4030 14870 4032 14922
rect 3976 14868 4032 14870
rect 4080 14922 4136 14924
rect 4080 14870 4082 14922
rect 4082 14870 4134 14922
rect 4134 14870 4136 14922
rect 4080 14868 4136 14870
rect 3836 14252 3892 14308
rect 4172 14306 4228 14308
rect 4172 14254 4174 14306
rect 4174 14254 4226 14306
rect 4226 14254 4228 14306
rect 4172 14252 4228 14254
rect 3500 13804 3556 13860
rect 5964 18396 6020 18452
rect 5068 18172 5124 18228
rect 9192 19626 9248 19628
rect 9192 19574 9194 19626
rect 9194 19574 9246 19626
rect 9246 19574 9248 19626
rect 9192 19572 9248 19574
rect 9296 19626 9352 19628
rect 9296 19574 9298 19626
rect 9298 19574 9350 19626
rect 9350 19574 9352 19626
rect 9296 19572 9352 19574
rect 9400 19626 9456 19628
rect 9400 19574 9402 19626
rect 9402 19574 9454 19626
rect 9454 19574 9456 19626
rect 9400 19572 9456 19574
rect 6748 19180 6804 19236
rect 6636 19010 6692 19012
rect 6636 18958 6638 19010
rect 6638 18958 6690 19010
rect 6690 18958 6692 19010
rect 6636 18956 6692 18958
rect 6532 18842 6588 18844
rect 6532 18790 6534 18842
rect 6534 18790 6586 18842
rect 6586 18790 6588 18842
rect 6532 18788 6588 18790
rect 6636 18842 6692 18844
rect 6636 18790 6638 18842
rect 6638 18790 6690 18842
rect 6690 18790 6692 18842
rect 6636 18788 6692 18790
rect 6740 18842 6796 18844
rect 6740 18790 6742 18842
rect 6742 18790 6794 18842
rect 6794 18790 6796 18842
rect 6740 18788 6796 18790
rect 7084 18956 7140 19012
rect 7420 19010 7476 19012
rect 7420 18958 7422 19010
rect 7422 18958 7474 19010
rect 7474 18958 7476 19010
rect 7420 18956 7476 18958
rect 6972 18450 7028 18452
rect 6972 18398 6974 18450
rect 6974 18398 7026 18450
rect 7026 18398 7028 18450
rect 6972 18396 7028 18398
rect 6860 18284 6916 18340
rect 4620 17442 4676 17444
rect 4620 17390 4622 17442
rect 4622 17390 4674 17442
rect 4674 17390 4676 17442
rect 4620 17388 4676 17390
rect 4396 16268 4452 16324
rect 4844 16268 4900 16324
rect 4620 16098 4676 16100
rect 4620 16046 4622 16098
rect 4622 16046 4674 16098
rect 4674 16046 4676 16098
rect 4620 16044 4676 16046
rect 5292 16268 5348 16324
rect 4620 14364 4676 14420
rect 4844 14476 4900 14532
rect 4284 13746 4340 13748
rect 4284 13694 4286 13746
rect 4286 13694 4338 13746
rect 4338 13694 4340 13746
rect 4284 13692 4340 13694
rect 4508 14140 4564 14196
rect 3872 13354 3928 13356
rect 3872 13302 3874 13354
rect 3874 13302 3926 13354
rect 3926 13302 3928 13354
rect 3872 13300 3928 13302
rect 3976 13354 4032 13356
rect 3976 13302 3978 13354
rect 3978 13302 4030 13354
rect 4030 13302 4032 13354
rect 3976 13300 4032 13302
rect 4080 13354 4136 13356
rect 4080 13302 4082 13354
rect 4082 13302 4134 13354
rect 4134 13302 4136 13354
rect 4080 13300 4136 13302
rect 4172 13132 4228 13188
rect 4732 13468 4788 13524
rect 4396 12572 4452 12628
rect 4284 12124 4340 12180
rect 4396 12348 4452 12404
rect 3872 11786 3928 11788
rect 3872 11734 3874 11786
rect 3874 11734 3926 11786
rect 3926 11734 3928 11786
rect 3872 11732 3928 11734
rect 3976 11786 4032 11788
rect 3976 11734 3978 11786
rect 3978 11734 4030 11786
rect 4030 11734 4032 11786
rect 3976 11732 4032 11734
rect 4080 11786 4136 11788
rect 4080 11734 4082 11786
rect 4082 11734 4134 11786
rect 4134 11734 4136 11786
rect 4080 11732 4136 11734
rect 4620 12402 4676 12404
rect 4620 12350 4622 12402
rect 4622 12350 4674 12402
rect 4674 12350 4676 12402
rect 4620 12348 4676 12350
rect 4508 12236 4564 12292
rect 3612 11340 3668 11396
rect 3388 11004 3444 11060
rect 3612 10892 3668 10948
rect 3276 10834 3332 10836
rect 3276 10782 3278 10834
rect 3278 10782 3330 10834
rect 3330 10782 3332 10834
rect 3276 10780 3332 10782
rect 2940 10668 2996 10724
rect 3164 9996 3220 10052
rect 3724 10668 3780 10724
rect 3388 9772 3444 9828
rect 3052 8764 3108 8820
rect 3164 9714 3220 9716
rect 3164 9662 3166 9714
rect 3166 9662 3218 9714
rect 3218 9662 3220 9714
rect 3164 9660 3220 9662
rect 4284 10780 4340 10836
rect 4620 12124 4676 12180
rect 3872 10218 3928 10220
rect 3872 10166 3874 10218
rect 3874 10166 3926 10218
rect 3926 10166 3928 10218
rect 3872 10164 3928 10166
rect 3976 10218 4032 10220
rect 3976 10166 3978 10218
rect 3978 10166 4030 10218
rect 4030 10166 4032 10218
rect 3976 10164 4032 10166
rect 4080 10218 4136 10220
rect 4080 10166 4082 10218
rect 4082 10166 4134 10218
rect 4134 10166 4136 10218
rect 4080 10164 4136 10166
rect 3836 9996 3892 10052
rect 7980 18956 8036 19012
rect 13580 20018 13636 20020
rect 13580 19966 13582 20018
rect 13582 19966 13634 20018
rect 13634 19966 13636 20018
rect 13580 19964 13636 19966
rect 11340 19852 11396 19908
rect 13692 19740 13748 19796
rect 11676 19180 11732 19236
rect 10780 19068 10836 19124
rect 9548 18956 9604 19012
rect 7644 18450 7700 18452
rect 7644 18398 7646 18450
rect 7646 18398 7698 18450
rect 7698 18398 7700 18450
rect 7644 18396 7700 18398
rect 7868 18226 7924 18228
rect 7868 18174 7870 18226
rect 7870 18174 7922 18226
rect 7922 18174 7924 18226
rect 7868 18172 7924 18174
rect 8428 18172 8484 18228
rect 9192 18058 9248 18060
rect 9192 18006 9194 18058
rect 9194 18006 9246 18058
rect 9246 18006 9248 18058
rect 9192 18004 9248 18006
rect 9296 18058 9352 18060
rect 9296 18006 9298 18058
rect 9298 18006 9350 18058
rect 9350 18006 9352 18058
rect 9296 18004 9352 18006
rect 9400 18058 9456 18060
rect 9400 18006 9402 18058
rect 9402 18006 9454 18058
rect 9454 18006 9456 18058
rect 9400 18004 9456 18006
rect 6636 17388 6692 17444
rect 8428 17388 8484 17444
rect 6532 17274 6588 17276
rect 6532 17222 6534 17274
rect 6534 17222 6586 17274
rect 6586 17222 6588 17274
rect 6532 17220 6588 17222
rect 6636 17274 6692 17276
rect 6636 17222 6638 17274
rect 6638 17222 6690 17274
rect 6690 17222 6692 17274
rect 6636 17220 6692 17222
rect 6740 17274 6796 17276
rect 6740 17222 6742 17274
rect 6742 17222 6794 17274
rect 6794 17222 6796 17274
rect 6740 17220 6796 17222
rect 6532 15706 6588 15708
rect 6532 15654 6534 15706
rect 6534 15654 6586 15706
rect 6586 15654 6588 15706
rect 6532 15652 6588 15654
rect 6636 15706 6692 15708
rect 6636 15654 6638 15706
rect 6638 15654 6690 15706
rect 6690 15654 6692 15706
rect 6636 15652 6692 15654
rect 6740 15706 6796 15708
rect 6740 15654 6742 15706
rect 6742 15654 6794 15706
rect 6794 15654 6796 15706
rect 6740 15652 6796 15654
rect 5404 13634 5460 13636
rect 5404 13582 5406 13634
rect 5406 13582 5458 13634
rect 5458 13582 5460 13634
rect 5404 13580 5460 13582
rect 6076 14364 6132 14420
rect 5516 13468 5572 13524
rect 4956 12796 5012 12852
rect 4508 9826 4564 9828
rect 4508 9774 4510 9826
rect 4510 9774 4562 9826
rect 4562 9774 4564 9826
rect 4508 9772 4564 9774
rect 6532 14138 6588 14140
rect 6532 14086 6534 14138
rect 6534 14086 6586 14138
rect 6586 14086 6588 14138
rect 6532 14084 6588 14086
rect 6636 14138 6692 14140
rect 6636 14086 6638 14138
rect 6638 14086 6690 14138
rect 6690 14086 6692 14138
rect 6636 14084 6692 14086
rect 6740 14138 6796 14140
rect 6740 14086 6742 14138
rect 6742 14086 6794 14138
rect 6794 14086 6796 14138
rect 6740 14084 6796 14086
rect 6188 13580 6244 13636
rect 9548 17388 9604 17444
rect 8876 16716 8932 16772
rect 9660 16994 9716 16996
rect 9660 16942 9662 16994
rect 9662 16942 9714 16994
rect 9714 16942 9716 16994
rect 9660 16940 9716 16942
rect 10892 18674 10948 18676
rect 10892 18622 10894 18674
rect 10894 18622 10946 18674
rect 10946 18622 10948 18674
rect 10892 18620 10948 18622
rect 10892 18284 10948 18340
rect 13468 19234 13524 19236
rect 13468 19182 13470 19234
rect 13470 19182 13522 19234
rect 13522 19182 13524 19234
rect 13468 19180 13524 19182
rect 14512 19626 14568 19628
rect 14512 19574 14514 19626
rect 14514 19574 14566 19626
rect 14566 19574 14568 19626
rect 14512 19572 14568 19574
rect 14616 19626 14672 19628
rect 14616 19574 14618 19626
rect 14618 19574 14670 19626
rect 14670 19574 14672 19626
rect 14616 19572 14672 19574
rect 14720 19626 14776 19628
rect 14720 19574 14722 19626
rect 14722 19574 14774 19626
rect 14774 19574 14776 19626
rect 14720 19572 14776 19574
rect 11852 18842 11908 18844
rect 11852 18790 11854 18842
rect 11854 18790 11906 18842
rect 11906 18790 11908 18842
rect 11852 18788 11908 18790
rect 11956 18842 12012 18844
rect 11956 18790 11958 18842
rect 11958 18790 12010 18842
rect 12010 18790 12012 18842
rect 11956 18788 12012 18790
rect 12060 18842 12116 18844
rect 12060 18790 12062 18842
rect 12062 18790 12114 18842
rect 12114 18790 12116 18842
rect 12060 18788 12116 18790
rect 13692 18620 13748 18676
rect 11228 18284 11284 18340
rect 13244 18450 13300 18452
rect 13244 18398 13246 18450
rect 13246 18398 13298 18450
rect 13298 18398 13300 18450
rect 13244 18396 13300 18398
rect 10332 17388 10388 17444
rect 10444 16716 10500 16772
rect 9192 16490 9248 16492
rect 9192 16438 9194 16490
rect 9194 16438 9246 16490
rect 9246 16438 9248 16490
rect 9192 16436 9248 16438
rect 9296 16490 9352 16492
rect 9296 16438 9298 16490
rect 9298 16438 9350 16490
rect 9350 16438 9352 16490
rect 9296 16436 9352 16438
rect 9400 16490 9456 16492
rect 9400 16438 9402 16490
rect 9402 16438 9454 16490
rect 9454 16438 9456 16490
rect 9400 16436 9456 16438
rect 8876 16044 8932 16100
rect 9772 16492 9828 16548
rect 10668 17442 10724 17444
rect 10668 17390 10670 17442
rect 10670 17390 10722 17442
rect 10722 17390 10724 17442
rect 10668 17388 10724 17390
rect 10892 16940 10948 16996
rect 11116 17500 11172 17556
rect 11228 17388 11284 17444
rect 11676 18338 11732 18340
rect 11676 18286 11678 18338
rect 11678 18286 11730 18338
rect 11730 18286 11732 18338
rect 11676 18284 11732 18286
rect 14028 18674 14084 18676
rect 14028 18622 14030 18674
rect 14030 18622 14082 18674
rect 14082 18622 14084 18674
rect 14028 18620 14084 18622
rect 14140 18450 14196 18452
rect 14140 18398 14142 18450
rect 14142 18398 14194 18450
rect 14194 18398 14196 18450
rect 14140 18396 14196 18398
rect 14364 18450 14420 18452
rect 14364 18398 14366 18450
rect 14366 18398 14418 18450
rect 14418 18398 14420 18450
rect 14364 18396 14420 18398
rect 11004 16828 11060 16884
rect 11340 16828 11396 16884
rect 8652 14418 8708 14420
rect 8652 14366 8654 14418
rect 8654 14366 8706 14418
rect 8706 14366 8708 14418
rect 8652 14364 8708 14366
rect 9192 14922 9248 14924
rect 9192 14870 9194 14922
rect 9194 14870 9246 14922
rect 9246 14870 9248 14922
rect 9192 14868 9248 14870
rect 9296 14922 9352 14924
rect 9296 14870 9298 14922
rect 9298 14870 9350 14922
rect 9350 14870 9352 14922
rect 9296 14868 9352 14870
rect 9400 14922 9456 14924
rect 9400 14870 9402 14922
rect 9402 14870 9454 14922
rect 9454 14870 9456 14922
rect 9400 14868 9456 14870
rect 9100 14476 9156 14532
rect 8876 14306 8932 14308
rect 8876 14254 8878 14306
rect 8878 14254 8930 14306
rect 8930 14254 8932 14306
rect 8876 14252 8932 14254
rect 8540 12738 8596 12740
rect 8540 12686 8542 12738
rect 8542 12686 8594 12738
rect 8594 12686 8596 12738
rect 8540 12684 8596 12686
rect 3948 9154 4004 9156
rect 3948 9102 3950 9154
rect 3950 9102 4002 9154
rect 4002 9102 4004 9154
rect 3948 9100 4004 9102
rect 3612 9042 3668 9044
rect 3612 8990 3614 9042
rect 3614 8990 3666 9042
rect 3666 8990 3668 9042
rect 3612 8988 3668 8990
rect 5068 9602 5124 9604
rect 5068 9550 5070 9602
rect 5070 9550 5122 9602
rect 5122 9550 5124 9602
rect 5068 9548 5124 9550
rect 4844 9212 4900 9268
rect 4172 8764 4228 8820
rect 3872 8650 3928 8652
rect 3872 8598 3874 8650
rect 3874 8598 3926 8650
rect 3926 8598 3928 8650
rect 3872 8596 3928 8598
rect 3976 8650 4032 8652
rect 3976 8598 3978 8650
rect 3978 8598 4030 8650
rect 4030 8598 4032 8650
rect 3976 8596 4032 8598
rect 4080 8650 4136 8652
rect 4080 8598 4082 8650
rect 4082 8598 4134 8650
rect 4134 8598 4136 8650
rect 4080 8596 4136 8598
rect 4508 8540 4564 8596
rect 3164 8092 3220 8148
rect 4956 8988 5012 9044
rect 5068 8930 5124 8932
rect 5068 8878 5070 8930
rect 5070 8878 5122 8930
rect 5122 8878 5124 8930
rect 5068 8876 5124 8878
rect 5068 8258 5124 8260
rect 5068 8206 5070 8258
rect 5070 8206 5122 8258
rect 5122 8206 5124 8258
rect 5068 8204 5124 8206
rect 6532 12570 6588 12572
rect 6532 12518 6534 12570
rect 6534 12518 6586 12570
rect 6586 12518 6588 12570
rect 6532 12516 6588 12518
rect 6636 12570 6692 12572
rect 6636 12518 6638 12570
rect 6638 12518 6690 12570
rect 6690 12518 6692 12570
rect 6636 12516 6692 12518
rect 6740 12570 6796 12572
rect 6740 12518 6742 12570
rect 6742 12518 6794 12570
rect 6794 12518 6796 12570
rect 6740 12516 6796 12518
rect 6532 11002 6588 11004
rect 6532 10950 6534 11002
rect 6534 10950 6586 11002
rect 6586 10950 6588 11002
rect 6532 10948 6588 10950
rect 6636 11002 6692 11004
rect 6636 10950 6638 11002
rect 6638 10950 6690 11002
rect 6690 10950 6692 11002
rect 6636 10948 6692 10950
rect 6740 11002 6796 11004
rect 6740 10950 6742 11002
rect 6742 10950 6794 11002
rect 6794 10950 6796 11002
rect 6740 10948 6796 10950
rect 9100 13580 9156 13636
rect 9772 14476 9828 14532
rect 9996 15148 10052 15204
rect 11004 15202 11060 15204
rect 11004 15150 11006 15202
rect 11006 15150 11058 15202
rect 11058 15150 11060 15202
rect 11004 15148 11060 15150
rect 9660 13970 9716 13972
rect 9660 13918 9662 13970
rect 9662 13918 9714 13970
rect 9714 13918 9716 13970
rect 9660 13916 9716 13918
rect 9884 13580 9940 13636
rect 9192 13354 9248 13356
rect 9192 13302 9194 13354
rect 9194 13302 9246 13354
rect 9246 13302 9248 13354
rect 9192 13300 9248 13302
rect 9296 13354 9352 13356
rect 9296 13302 9298 13354
rect 9298 13302 9350 13354
rect 9350 13302 9352 13354
rect 9296 13300 9352 13302
rect 9400 13354 9456 13356
rect 9400 13302 9402 13354
rect 9402 13302 9454 13354
rect 9454 13302 9456 13354
rect 9400 13300 9456 13302
rect 9212 12684 9268 12740
rect 8652 11954 8708 11956
rect 8652 11902 8654 11954
rect 8654 11902 8706 11954
rect 8706 11902 8708 11954
rect 8652 11900 8708 11902
rect 8540 10780 8596 10836
rect 5740 9548 5796 9604
rect 5516 8876 5572 8932
rect 5740 8258 5796 8260
rect 5740 8206 5742 8258
rect 5742 8206 5794 8258
rect 5794 8206 5796 8258
rect 5740 8204 5796 8206
rect 5964 9266 6020 9268
rect 5964 9214 5966 9266
rect 5966 9214 6018 9266
rect 6018 9214 6020 9266
rect 5964 9212 6020 9214
rect 6532 9434 6588 9436
rect 6532 9382 6534 9434
rect 6534 9382 6586 9434
rect 6586 9382 6588 9434
rect 6532 9380 6588 9382
rect 6636 9434 6692 9436
rect 6636 9382 6638 9434
rect 6638 9382 6690 9434
rect 6690 9382 6692 9434
rect 6636 9380 6692 9382
rect 6740 9434 6796 9436
rect 6740 9382 6742 9434
rect 6742 9382 6794 9434
rect 6794 9382 6796 9434
rect 6740 9380 6796 9382
rect 6524 9042 6580 9044
rect 6524 8990 6526 9042
rect 6526 8990 6578 9042
rect 6578 8990 6580 9042
rect 6524 8988 6580 8990
rect 6076 8930 6132 8932
rect 6076 8878 6078 8930
rect 6078 8878 6130 8930
rect 6130 8878 6132 8930
rect 6076 8876 6132 8878
rect 6076 8540 6132 8596
rect 6188 8764 6244 8820
rect 5964 8428 6020 8484
rect 6076 8092 6132 8148
rect 3872 7082 3928 7084
rect 3872 7030 3874 7082
rect 3874 7030 3926 7082
rect 3926 7030 3928 7082
rect 3872 7028 3928 7030
rect 3976 7082 4032 7084
rect 3976 7030 3978 7082
rect 3978 7030 4030 7082
rect 4030 7030 4032 7082
rect 3976 7028 4032 7030
rect 4080 7082 4136 7084
rect 4080 7030 4082 7082
rect 4082 7030 4134 7082
rect 4134 7030 4136 7082
rect 4080 7028 4136 7030
rect 4956 7308 5012 7364
rect 4844 6972 4900 7028
rect 4844 6748 4900 6804
rect 5628 7362 5684 7364
rect 5628 7310 5630 7362
rect 5630 7310 5682 7362
rect 5682 7310 5684 7362
rect 5628 7308 5684 7310
rect 5628 6972 5684 7028
rect 5740 6802 5796 6804
rect 5740 6750 5742 6802
rect 5742 6750 5794 6802
rect 5794 6750 5796 6802
rect 5740 6748 5796 6750
rect 5964 6524 6020 6580
rect 6532 7866 6588 7868
rect 6532 7814 6534 7866
rect 6534 7814 6586 7866
rect 6586 7814 6588 7866
rect 6532 7812 6588 7814
rect 6636 7866 6692 7868
rect 6636 7814 6638 7866
rect 6638 7814 6690 7866
rect 6690 7814 6692 7866
rect 6636 7812 6692 7814
rect 6740 7866 6796 7868
rect 6740 7814 6742 7866
rect 6742 7814 6794 7866
rect 6794 7814 6796 7866
rect 6740 7812 6796 7814
rect 6412 6524 6468 6580
rect 6532 6298 6588 6300
rect 6532 6246 6534 6298
rect 6534 6246 6586 6298
rect 6586 6246 6588 6298
rect 6532 6244 6588 6246
rect 6636 6298 6692 6300
rect 6636 6246 6638 6298
rect 6638 6246 6690 6298
rect 6690 6246 6692 6298
rect 6636 6244 6692 6246
rect 6740 6298 6796 6300
rect 6740 6246 6742 6298
rect 6742 6246 6794 6298
rect 6794 6246 6796 6298
rect 6740 6244 6796 6246
rect 9192 11786 9248 11788
rect 9192 11734 9194 11786
rect 9194 11734 9246 11786
rect 9246 11734 9248 11786
rect 9192 11732 9248 11734
rect 9296 11786 9352 11788
rect 9296 11734 9298 11786
rect 9298 11734 9350 11786
rect 9350 11734 9352 11786
rect 9296 11732 9352 11734
rect 9400 11786 9456 11788
rect 9400 11734 9402 11786
rect 9402 11734 9454 11786
rect 9454 11734 9456 11786
rect 9400 11732 9456 11734
rect 9772 11788 9828 11844
rect 9548 10834 9604 10836
rect 9548 10782 9550 10834
rect 9550 10782 9602 10834
rect 9602 10782 9604 10834
rect 9548 10780 9604 10782
rect 9192 10218 9248 10220
rect 9192 10166 9194 10218
rect 9194 10166 9246 10218
rect 9246 10166 9248 10218
rect 9192 10164 9248 10166
rect 9296 10218 9352 10220
rect 9296 10166 9298 10218
rect 9298 10166 9350 10218
rect 9350 10166 9352 10218
rect 9296 10164 9352 10166
rect 9400 10218 9456 10220
rect 9400 10166 9402 10218
rect 9402 10166 9454 10218
rect 9454 10166 9456 10218
rect 9400 10164 9456 10166
rect 9324 10050 9380 10052
rect 9324 9998 9326 10050
rect 9326 9998 9378 10050
rect 9378 9998 9380 10050
rect 9324 9996 9380 9998
rect 10220 13468 10276 13524
rect 10892 14252 10948 14308
rect 10556 13356 10612 13412
rect 9996 12460 10052 12516
rect 9996 12124 10052 12180
rect 10444 12962 10500 12964
rect 10444 12910 10446 12962
rect 10446 12910 10498 12962
rect 10498 12910 10500 12962
rect 10444 12908 10500 12910
rect 11116 13356 11172 13412
rect 10444 12460 10500 12516
rect 10444 12178 10500 12180
rect 10444 12126 10446 12178
rect 10446 12126 10498 12178
rect 10498 12126 10500 12178
rect 10444 12124 10500 12126
rect 10556 11564 10612 11620
rect 9772 10108 9828 10164
rect 9884 9826 9940 9828
rect 9884 9774 9886 9826
rect 9886 9774 9938 9826
rect 9938 9774 9940 9826
rect 9884 9772 9940 9774
rect 9548 9714 9604 9716
rect 9548 9662 9550 9714
rect 9550 9662 9602 9714
rect 9602 9662 9604 9714
rect 9548 9660 9604 9662
rect 10332 11228 10388 11284
rect 9436 8764 9492 8820
rect 10332 9772 10388 9828
rect 9192 8650 9248 8652
rect 9192 8598 9194 8650
rect 9194 8598 9246 8650
rect 9246 8598 9248 8650
rect 9192 8596 9248 8598
rect 9296 8650 9352 8652
rect 9296 8598 9298 8650
rect 9298 8598 9350 8650
rect 9350 8598 9352 8650
rect 9296 8596 9352 8598
rect 9400 8650 9456 8652
rect 9400 8598 9402 8650
rect 9402 8598 9454 8650
rect 9454 8598 9456 8650
rect 9400 8596 9456 8598
rect 8988 8316 9044 8372
rect 9996 9100 10052 9156
rect 9884 8370 9940 8372
rect 9884 8318 9886 8370
rect 9886 8318 9938 8370
rect 9938 8318 9940 8370
rect 9884 8316 9940 8318
rect 9660 8258 9716 8260
rect 9660 8206 9662 8258
rect 9662 8206 9714 8258
rect 9714 8206 9716 8258
rect 9660 8204 9716 8206
rect 10108 8818 10164 8820
rect 10108 8766 10110 8818
rect 10110 8766 10162 8818
rect 10162 8766 10164 8818
rect 10108 8764 10164 8766
rect 10332 8764 10388 8820
rect 10444 9660 10500 9716
rect 10444 8652 10500 8708
rect 10780 12066 10836 12068
rect 10780 12014 10782 12066
rect 10782 12014 10834 12066
rect 10834 12014 10836 12066
rect 10780 12012 10836 12014
rect 10892 11900 10948 11956
rect 10780 11116 10836 11172
rect 10668 8930 10724 8932
rect 10668 8878 10670 8930
rect 10670 8878 10722 8930
rect 10722 8878 10724 8930
rect 10668 8876 10724 8878
rect 10108 8428 10164 8484
rect 10444 8428 10500 8484
rect 10668 8316 10724 8372
rect 10332 8204 10388 8260
rect 10220 8146 10276 8148
rect 10220 8094 10222 8146
rect 10222 8094 10274 8146
rect 10274 8094 10276 8146
rect 10220 8092 10276 8094
rect 10108 7980 10164 8036
rect 9660 7308 9716 7364
rect 9192 7082 9248 7084
rect 9192 7030 9194 7082
rect 9194 7030 9246 7082
rect 9246 7030 9248 7082
rect 9192 7028 9248 7030
rect 9296 7082 9352 7084
rect 9296 7030 9298 7082
rect 9298 7030 9350 7082
rect 9350 7030 9352 7082
rect 9296 7028 9352 7030
rect 9400 7082 9456 7084
rect 9400 7030 9402 7082
rect 9402 7030 9454 7082
rect 9454 7030 9456 7082
rect 9400 7028 9456 7030
rect 9436 6860 9492 6916
rect 8540 6076 8596 6132
rect 10668 7980 10724 8036
rect 9996 6860 10052 6916
rect 10332 6860 10388 6916
rect 10220 6690 10276 6692
rect 10220 6638 10222 6690
rect 10222 6638 10274 6690
rect 10274 6638 10276 6690
rect 10220 6636 10276 6638
rect 11564 17554 11620 17556
rect 11564 17502 11566 17554
rect 11566 17502 11618 17554
rect 11618 17502 11620 17554
rect 11564 17500 11620 17502
rect 11852 17274 11908 17276
rect 11852 17222 11854 17274
rect 11854 17222 11906 17274
rect 11906 17222 11908 17274
rect 11852 17220 11908 17222
rect 11956 17274 12012 17276
rect 11956 17222 11958 17274
rect 11958 17222 12010 17274
rect 12010 17222 12012 17274
rect 11956 17220 12012 17222
rect 12060 17274 12116 17276
rect 12060 17222 12062 17274
rect 12062 17222 12114 17274
rect 12114 17222 12116 17274
rect 12060 17220 12116 17222
rect 11788 16940 11844 16996
rect 14512 18058 14568 18060
rect 14512 18006 14514 18058
rect 14514 18006 14566 18058
rect 14566 18006 14568 18058
rect 14512 18004 14568 18006
rect 14616 18058 14672 18060
rect 14616 18006 14618 18058
rect 14618 18006 14670 18058
rect 14670 18006 14672 18058
rect 14616 18004 14672 18006
rect 14720 18058 14776 18060
rect 14720 18006 14722 18058
rect 14722 18006 14774 18058
rect 14774 18006 14776 18058
rect 14720 18004 14776 18006
rect 17948 19740 18004 19796
rect 18508 19964 18564 20020
rect 17948 19234 18004 19236
rect 17948 19182 17950 19234
rect 17950 19182 18002 19234
rect 18002 19182 18004 19234
rect 17948 19180 18004 19182
rect 19852 19852 19908 19908
rect 19832 19626 19888 19628
rect 19832 19574 19834 19626
rect 19834 19574 19886 19626
rect 19886 19574 19888 19626
rect 19832 19572 19888 19574
rect 19936 19626 19992 19628
rect 19936 19574 19938 19626
rect 19938 19574 19990 19626
rect 19990 19574 19992 19626
rect 19936 19572 19992 19574
rect 20040 19626 20096 19628
rect 20040 19574 20042 19626
rect 20042 19574 20094 19626
rect 20094 19574 20096 19626
rect 20040 19572 20096 19574
rect 18396 19122 18452 19124
rect 18396 19070 18398 19122
rect 18398 19070 18450 19122
rect 18450 19070 18452 19122
rect 18396 19068 18452 19070
rect 19292 19234 19348 19236
rect 19292 19182 19294 19234
rect 19294 19182 19346 19234
rect 19346 19182 19348 19234
rect 19292 19180 19348 19182
rect 19180 19122 19236 19124
rect 19180 19070 19182 19122
rect 19182 19070 19234 19122
rect 19234 19070 19236 19122
rect 19180 19068 19236 19070
rect 20636 19180 20692 19236
rect 19404 19010 19460 19012
rect 19404 18958 19406 19010
rect 19406 18958 19458 19010
rect 19458 18958 19460 19010
rect 19404 18956 19460 18958
rect 17172 18842 17228 18844
rect 17172 18790 17174 18842
rect 17174 18790 17226 18842
rect 17226 18790 17228 18842
rect 17172 18788 17228 18790
rect 17276 18842 17332 18844
rect 17276 18790 17278 18842
rect 17278 18790 17330 18842
rect 17330 18790 17332 18842
rect 17276 18788 17332 18790
rect 17380 18842 17436 18844
rect 17380 18790 17382 18842
rect 17382 18790 17434 18842
rect 17434 18790 17436 18842
rect 17380 18788 17436 18790
rect 15596 18396 15652 18452
rect 15932 18284 15988 18340
rect 16044 18396 16100 18452
rect 13132 16940 13188 16996
rect 12236 16882 12292 16884
rect 12236 16830 12238 16882
rect 12238 16830 12290 16882
rect 12290 16830 12292 16882
rect 12236 16828 12292 16830
rect 11452 16716 11508 16772
rect 14512 16490 14568 16492
rect 14512 16438 14514 16490
rect 14514 16438 14566 16490
rect 14566 16438 14568 16490
rect 14512 16436 14568 16438
rect 14616 16490 14672 16492
rect 14616 16438 14618 16490
rect 14618 16438 14670 16490
rect 14670 16438 14672 16490
rect 14616 16436 14672 16438
rect 14720 16490 14776 16492
rect 14720 16438 14722 16490
rect 14722 16438 14774 16490
rect 14774 16438 14776 16490
rect 14720 16436 14776 16438
rect 15036 16322 15092 16324
rect 15036 16270 15038 16322
rect 15038 16270 15090 16322
rect 15090 16270 15092 16322
rect 15036 16268 15092 16270
rect 14140 16044 14196 16100
rect 11852 15706 11908 15708
rect 11852 15654 11854 15706
rect 11854 15654 11906 15706
rect 11906 15654 11908 15706
rect 11852 15652 11908 15654
rect 11956 15706 12012 15708
rect 11956 15654 11958 15706
rect 11958 15654 12010 15706
rect 12010 15654 12012 15706
rect 11956 15652 12012 15654
rect 12060 15706 12116 15708
rect 12060 15654 12062 15706
rect 12062 15654 12114 15706
rect 12114 15654 12116 15706
rect 12060 15652 12116 15654
rect 11452 15372 11508 15428
rect 14924 16098 14980 16100
rect 14924 16046 14926 16098
rect 14926 16046 14978 16098
rect 14978 16046 14980 16098
rect 14924 16044 14980 16046
rect 15484 16268 15540 16324
rect 14476 15426 14532 15428
rect 14476 15374 14478 15426
rect 14478 15374 14530 15426
rect 14530 15374 14532 15426
rect 14476 15372 14532 15374
rect 15932 16268 15988 16324
rect 15036 15148 15092 15204
rect 14512 14922 14568 14924
rect 14512 14870 14514 14922
rect 14514 14870 14566 14922
rect 14566 14870 14568 14922
rect 14512 14868 14568 14870
rect 14616 14922 14672 14924
rect 14616 14870 14618 14922
rect 14618 14870 14670 14922
rect 14670 14870 14672 14922
rect 14616 14868 14672 14870
rect 14720 14922 14776 14924
rect 14720 14870 14722 14922
rect 14722 14870 14774 14922
rect 14774 14870 14776 14922
rect 14720 14868 14776 14870
rect 13804 14476 13860 14532
rect 11852 14138 11908 14140
rect 11852 14086 11854 14138
rect 11854 14086 11906 14138
rect 11906 14086 11908 14138
rect 11852 14084 11908 14086
rect 11956 14138 12012 14140
rect 11956 14086 11958 14138
rect 11958 14086 12010 14138
rect 12010 14086 12012 14138
rect 11956 14084 12012 14086
rect 12060 14138 12116 14140
rect 12060 14086 12062 14138
rect 12062 14086 12114 14138
rect 12114 14086 12116 14138
rect 12060 14084 12116 14086
rect 12236 13468 12292 13524
rect 11452 12908 11508 12964
rect 11340 12066 11396 12068
rect 11340 12014 11342 12066
rect 11342 12014 11394 12066
rect 11394 12014 11396 12066
rect 11340 12012 11396 12014
rect 11228 11954 11284 11956
rect 11228 11902 11230 11954
rect 11230 11902 11282 11954
rect 11282 11902 11284 11954
rect 11228 11900 11284 11902
rect 11116 8988 11172 9044
rect 11004 8652 11060 8708
rect 11004 8146 11060 8148
rect 11004 8094 11006 8146
rect 11006 8094 11058 8146
rect 11058 8094 11060 8146
rect 11004 8092 11060 8094
rect 11116 7980 11172 8036
rect 10892 6860 10948 6916
rect 11004 7868 11060 7924
rect 10892 6412 10948 6468
rect 11340 8370 11396 8372
rect 11340 8318 11342 8370
rect 11342 8318 11394 8370
rect 11394 8318 11396 8370
rect 11340 8316 11396 8318
rect 11340 7532 11396 7588
rect 11852 12570 11908 12572
rect 11852 12518 11854 12570
rect 11854 12518 11906 12570
rect 11906 12518 11908 12570
rect 11852 12516 11908 12518
rect 11956 12570 12012 12572
rect 11956 12518 11958 12570
rect 11958 12518 12010 12570
rect 12010 12518 12012 12570
rect 11956 12516 12012 12518
rect 12060 12570 12116 12572
rect 12060 12518 12062 12570
rect 12062 12518 12114 12570
rect 12114 12518 12116 12570
rect 12060 12516 12116 12518
rect 11564 11676 11620 11732
rect 11676 11564 11732 11620
rect 14140 14364 14196 14420
rect 14700 14530 14756 14532
rect 14700 14478 14702 14530
rect 14702 14478 14754 14530
rect 14754 14478 14756 14530
rect 14700 14476 14756 14478
rect 14140 13468 14196 13524
rect 14476 14252 14532 14308
rect 14252 13132 14308 13188
rect 13804 12012 13860 12068
rect 12572 11676 12628 11732
rect 13692 11676 13748 11732
rect 15484 14924 15540 14980
rect 15036 14306 15092 14308
rect 15036 14254 15038 14306
rect 15038 14254 15090 14306
rect 15090 14254 15092 14306
rect 15036 14252 15092 14254
rect 14512 13354 14568 13356
rect 14512 13302 14514 13354
rect 14514 13302 14566 13354
rect 14566 13302 14568 13354
rect 14512 13300 14568 13302
rect 14616 13354 14672 13356
rect 14616 13302 14618 13354
rect 14618 13302 14670 13354
rect 14670 13302 14672 13354
rect 14616 13300 14672 13302
rect 14720 13354 14776 13356
rect 14720 13302 14722 13354
rect 14722 13302 14774 13354
rect 14774 13302 14776 13354
rect 14720 13300 14776 13302
rect 14924 13356 14980 13412
rect 14588 13186 14644 13188
rect 14588 13134 14590 13186
rect 14590 13134 14642 13186
rect 14642 13134 14644 13186
rect 14588 13132 14644 13134
rect 15372 14476 15428 14532
rect 15820 15036 15876 15092
rect 15708 14252 15764 14308
rect 16268 18284 16324 18340
rect 16604 18172 16660 18228
rect 17172 17274 17228 17276
rect 17172 17222 17174 17274
rect 17174 17222 17226 17274
rect 17226 17222 17228 17274
rect 17172 17220 17228 17222
rect 17276 17274 17332 17276
rect 17276 17222 17278 17274
rect 17278 17222 17330 17274
rect 17330 17222 17332 17274
rect 17276 17220 17332 17222
rect 17380 17274 17436 17276
rect 17380 17222 17382 17274
rect 17382 17222 17434 17274
rect 17434 17222 17436 17274
rect 17380 17220 17436 17222
rect 17172 15706 17228 15708
rect 17172 15654 17174 15706
rect 17174 15654 17226 15706
rect 17226 15654 17228 15706
rect 17172 15652 17228 15654
rect 17276 15706 17332 15708
rect 17276 15654 17278 15706
rect 17278 15654 17330 15706
rect 17330 15654 17332 15706
rect 17276 15652 17332 15654
rect 17380 15706 17436 15708
rect 17380 15654 17382 15706
rect 17382 15654 17434 15706
rect 17434 15654 17436 15706
rect 17380 15652 17436 15654
rect 19516 18172 19572 18228
rect 19832 18058 19888 18060
rect 19832 18006 19834 18058
rect 19834 18006 19886 18058
rect 19886 18006 19888 18058
rect 19832 18004 19888 18006
rect 19936 18058 19992 18060
rect 19936 18006 19938 18058
rect 19938 18006 19990 18058
rect 19990 18006 19992 18058
rect 19936 18004 19992 18006
rect 20040 18058 20096 18060
rect 20040 18006 20042 18058
rect 20042 18006 20094 18058
rect 20094 18006 20096 18058
rect 20040 18004 20096 18006
rect 19516 17778 19572 17780
rect 19516 17726 19518 17778
rect 19518 17726 19570 17778
rect 19570 17726 19572 17778
rect 19516 17724 19572 17726
rect 19852 17890 19908 17892
rect 19852 17838 19854 17890
rect 19854 17838 19906 17890
rect 19906 17838 19908 17890
rect 19852 17836 19908 17838
rect 20636 17836 20692 17892
rect 19964 17778 20020 17780
rect 19964 17726 19966 17778
rect 19966 17726 20018 17778
rect 20018 17726 20020 17778
rect 19964 17724 20020 17726
rect 19404 16882 19460 16884
rect 19404 16830 19406 16882
rect 19406 16830 19458 16882
rect 19458 16830 19460 16882
rect 19404 16828 19460 16830
rect 19740 16658 19796 16660
rect 19740 16606 19742 16658
rect 19742 16606 19794 16658
rect 19794 16606 19796 16658
rect 19740 16604 19796 16606
rect 20188 16828 20244 16884
rect 20524 16940 20580 16996
rect 19832 16490 19888 16492
rect 19832 16438 19834 16490
rect 19834 16438 19886 16490
rect 19886 16438 19888 16490
rect 19832 16436 19888 16438
rect 19936 16490 19992 16492
rect 19936 16438 19938 16490
rect 19938 16438 19990 16490
rect 19990 16438 19992 16490
rect 19936 16436 19992 16438
rect 20040 16490 20096 16492
rect 20040 16438 20042 16490
rect 20042 16438 20094 16490
rect 20094 16438 20096 16490
rect 20040 16436 20096 16438
rect 19180 16098 19236 16100
rect 19180 16046 19182 16098
rect 19182 16046 19234 16098
rect 19234 16046 19236 16098
rect 19180 16044 19236 16046
rect 19740 16322 19796 16324
rect 19740 16270 19742 16322
rect 19742 16270 19794 16322
rect 19794 16270 19796 16322
rect 19740 16268 19796 16270
rect 20300 16604 20356 16660
rect 19628 16210 19684 16212
rect 19628 16158 19630 16210
rect 19630 16158 19682 16210
rect 19682 16158 19684 16210
rect 19628 16156 19684 16158
rect 18844 15260 18900 15316
rect 16044 14924 16100 14980
rect 15372 13132 15428 13188
rect 14476 12850 14532 12852
rect 14476 12798 14478 12850
rect 14478 12798 14530 12850
rect 14530 12798 14532 12850
rect 14476 12796 14532 12798
rect 14512 11786 14568 11788
rect 14512 11734 14514 11786
rect 14514 11734 14566 11786
rect 14566 11734 14568 11786
rect 14512 11732 14568 11734
rect 14616 11786 14672 11788
rect 14616 11734 14618 11786
rect 14618 11734 14670 11786
rect 14670 11734 14672 11786
rect 14616 11732 14672 11734
rect 14720 11786 14776 11788
rect 14720 11734 14722 11786
rect 14722 11734 14774 11786
rect 14774 11734 14776 11786
rect 14720 11732 14776 11734
rect 15148 12684 15204 12740
rect 15932 12962 15988 12964
rect 15932 12910 15934 12962
rect 15934 12910 15986 12962
rect 15986 12910 15988 12962
rect 15932 12908 15988 12910
rect 15372 12236 15428 12292
rect 14924 11676 14980 11732
rect 15260 12124 15316 12180
rect 13692 11452 13748 11508
rect 11852 11002 11908 11004
rect 11852 10950 11854 11002
rect 11854 10950 11906 11002
rect 11906 10950 11908 11002
rect 11852 10948 11908 10950
rect 11956 11002 12012 11004
rect 11956 10950 11958 11002
rect 11958 10950 12010 11002
rect 12010 10950 12012 11002
rect 11956 10948 12012 10950
rect 12060 11002 12116 11004
rect 12060 10950 12062 11002
rect 12062 10950 12114 11002
rect 12114 10950 12116 11002
rect 12060 10948 12116 10950
rect 13468 11282 13524 11284
rect 13468 11230 13470 11282
rect 13470 11230 13522 11282
rect 13522 11230 13524 11282
rect 13468 11228 13524 11230
rect 14252 11228 14308 11284
rect 12460 10780 12516 10836
rect 13580 11170 13636 11172
rect 13580 11118 13582 11170
rect 13582 11118 13634 11170
rect 13634 11118 13636 11170
rect 13580 11116 13636 11118
rect 12572 10108 12628 10164
rect 11852 9434 11908 9436
rect 11852 9382 11854 9434
rect 11854 9382 11906 9434
rect 11906 9382 11908 9434
rect 11852 9380 11908 9382
rect 11956 9434 12012 9436
rect 11956 9382 11958 9434
rect 11958 9382 12010 9434
rect 12010 9382 12012 9434
rect 11956 9380 12012 9382
rect 12060 9434 12116 9436
rect 12060 9382 12062 9434
rect 12062 9382 12114 9434
rect 12114 9382 12116 9434
rect 12060 9380 12116 9382
rect 14252 8764 14308 8820
rect 11564 8258 11620 8260
rect 11564 8206 11566 8258
rect 11566 8206 11618 8258
rect 11618 8206 11620 8258
rect 11564 8204 11620 8206
rect 14924 11228 14980 11284
rect 15036 11004 15092 11060
rect 14476 10780 14532 10836
rect 15260 11004 15316 11060
rect 15484 11452 15540 11508
rect 15820 11452 15876 11508
rect 15260 10332 15316 10388
rect 14512 10218 14568 10220
rect 14512 10166 14514 10218
rect 14514 10166 14566 10218
rect 14566 10166 14568 10218
rect 14512 10164 14568 10166
rect 14616 10218 14672 10220
rect 14616 10166 14618 10218
rect 14618 10166 14670 10218
rect 14670 10166 14672 10218
rect 14616 10164 14672 10166
rect 14720 10218 14776 10220
rect 14720 10166 14722 10218
rect 14722 10166 14774 10218
rect 14774 10166 14776 10218
rect 14720 10164 14776 10166
rect 15596 9772 15652 9828
rect 14512 8650 14568 8652
rect 14512 8598 14514 8650
rect 14514 8598 14566 8650
rect 14566 8598 14568 8650
rect 14512 8596 14568 8598
rect 14616 8650 14672 8652
rect 14616 8598 14618 8650
rect 14618 8598 14670 8650
rect 14670 8598 14672 8650
rect 14616 8596 14672 8598
rect 14720 8650 14776 8652
rect 14720 8598 14722 8650
rect 14722 8598 14774 8650
rect 14774 8598 14776 8650
rect 14720 8596 14776 8598
rect 14364 8428 14420 8484
rect 16156 12124 16212 12180
rect 16268 12236 16324 12292
rect 16156 11676 16212 11732
rect 11852 7866 11908 7868
rect 11852 7814 11854 7866
rect 11854 7814 11906 7866
rect 11906 7814 11908 7866
rect 11852 7812 11908 7814
rect 11956 7866 12012 7868
rect 11956 7814 11958 7866
rect 11958 7814 12010 7866
rect 12010 7814 12012 7866
rect 11956 7812 12012 7814
rect 12060 7866 12116 7868
rect 12060 7814 12062 7866
rect 12062 7814 12114 7866
rect 12114 7814 12116 7866
rect 12060 7812 12116 7814
rect 11788 7644 11844 7700
rect 14588 8034 14644 8036
rect 14588 7982 14590 8034
rect 14590 7982 14642 8034
rect 14642 7982 14644 8034
rect 14588 7980 14644 7982
rect 15148 7868 15204 7924
rect 15372 8258 15428 8260
rect 15372 8206 15374 8258
rect 15374 8206 15426 8258
rect 15426 8206 15428 8258
rect 15372 8204 15428 8206
rect 9884 6018 9940 6020
rect 9884 5966 9886 6018
rect 9886 5966 9938 6018
rect 9938 5966 9940 6018
rect 9884 5964 9940 5966
rect 10332 6018 10388 6020
rect 10332 5966 10334 6018
rect 10334 5966 10386 6018
rect 10386 5966 10388 6018
rect 10332 5964 10388 5966
rect 11452 6690 11508 6692
rect 11452 6638 11454 6690
rect 11454 6638 11506 6690
rect 11506 6638 11508 6690
rect 11452 6636 11508 6638
rect 16268 8258 16324 8260
rect 16268 8206 16270 8258
rect 16270 8206 16322 8258
rect 16322 8206 16324 8258
rect 16268 8204 16324 8206
rect 15484 8092 15540 8148
rect 16268 8034 16324 8036
rect 16268 7982 16270 8034
rect 16270 7982 16322 8034
rect 16322 7982 16324 8034
rect 16268 7980 16324 7982
rect 16940 14924 16996 14980
rect 17172 14138 17228 14140
rect 17172 14086 17174 14138
rect 17174 14086 17226 14138
rect 17226 14086 17228 14138
rect 17172 14084 17228 14086
rect 17276 14138 17332 14140
rect 17276 14086 17278 14138
rect 17278 14086 17330 14138
rect 17330 14086 17332 14138
rect 17276 14084 17332 14086
rect 17380 14138 17436 14140
rect 17380 14086 17382 14138
rect 17382 14086 17434 14138
rect 17434 14086 17436 14138
rect 17380 14084 17436 14086
rect 17612 15202 17668 15204
rect 17612 15150 17614 15202
rect 17614 15150 17666 15202
rect 17666 15150 17668 15202
rect 17612 15148 17668 15150
rect 17836 15202 17892 15204
rect 17836 15150 17838 15202
rect 17838 15150 17890 15202
rect 17890 15150 17892 15202
rect 17836 15148 17892 15150
rect 17500 13356 17556 13412
rect 17172 12570 17228 12572
rect 17172 12518 17174 12570
rect 17174 12518 17226 12570
rect 17226 12518 17228 12570
rect 17172 12516 17228 12518
rect 17276 12570 17332 12572
rect 17276 12518 17278 12570
rect 17278 12518 17330 12570
rect 17330 12518 17332 12570
rect 17276 12516 17332 12518
rect 17380 12570 17436 12572
rect 17380 12518 17382 12570
rect 17382 12518 17434 12570
rect 17434 12518 17436 12570
rect 17380 12516 17436 12518
rect 17164 12124 17220 12180
rect 17052 11618 17108 11620
rect 17052 11566 17054 11618
rect 17054 11566 17106 11618
rect 17106 11566 17108 11618
rect 17052 11564 17108 11566
rect 17388 11676 17444 11732
rect 17612 11394 17668 11396
rect 17612 11342 17614 11394
rect 17614 11342 17666 11394
rect 17666 11342 17668 11394
rect 17612 11340 17668 11342
rect 16492 11282 16548 11284
rect 16492 11230 16494 11282
rect 16494 11230 16546 11282
rect 16546 11230 16548 11282
rect 16492 11228 16548 11230
rect 17172 11002 17228 11004
rect 17172 10950 17174 11002
rect 17174 10950 17226 11002
rect 17226 10950 17228 11002
rect 17172 10948 17228 10950
rect 17276 11002 17332 11004
rect 17276 10950 17278 11002
rect 17278 10950 17330 11002
rect 17330 10950 17332 11002
rect 17276 10948 17332 10950
rect 17380 11002 17436 11004
rect 17380 10950 17382 11002
rect 17382 10950 17434 11002
rect 17434 10950 17436 11002
rect 17380 10948 17436 10950
rect 17172 9434 17228 9436
rect 17172 9382 17174 9434
rect 17174 9382 17226 9434
rect 17226 9382 17228 9434
rect 17172 9380 17228 9382
rect 17276 9434 17332 9436
rect 17276 9382 17278 9434
rect 17278 9382 17330 9434
rect 17330 9382 17332 9434
rect 17276 9380 17332 9382
rect 17380 9434 17436 9436
rect 17380 9382 17382 9434
rect 17382 9382 17434 9434
rect 17434 9382 17436 9434
rect 17380 9380 17436 9382
rect 17948 15036 18004 15092
rect 18284 13356 18340 13412
rect 18060 12178 18116 12180
rect 18060 12126 18062 12178
rect 18062 12126 18114 12178
rect 18114 12126 18116 12178
rect 18060 12124 18116 12126
rect 17948 11452 18004 11508
rect 19516 15314 19572 15316
rect 19516 15262 19518 15314
rect 19518 15262 19570 15314
rect 19570 15262 19572 15314
rect 19516 15260 19572 15262
rect 19964 15538 20020 15540
rect 19964 15486 19966 15538
rect 19966 15486 20018 15538
rect 20018 15486 20020 15538
rect 19964 15484 20020 15486
rect 19740 15372 19796 15428
rect 20300 15314 20356 15316
rect 20300 15262 20302 15314
rect 20302 15262 20354 15314
rect 20354 15262 20356 15314
rect 20300 15260 20356 15262
rect 19740 15148 19796 15204
rect 19832 14922 19888 14924
rect 19832 14870 19834 14922
rect 19834 14870 19886 14922
rect 19886 14870 19888 14922
rect 19832 14868 19888 14870
rect 19936 14922 19992 14924
rect 19936 14870 19938 14922
rect 19938 14870 19990 14922
rect 19990 14870 19992 14922
rect 19936 14868 19992 14870
rect 20040 14922 20096 14924
rect 20040 14870 20042 14922
rect 20042 14870 20094 14922
rect 20094 14870 20096 14922
rect 20040 14868 20096 14870
rect 19180 13916 19236 13972
rect 19832 13354 19888 13356
rect 19832 13302 19834 13354
rect 19834 13302 19886 13354
rect 19886 13302 19888 13354
rect 19832 13300 19888 13302
rect 19936 13354 19992 13356
rect 19936 13302 19938 13354
rect 19938 13302 19990 13354
rect 19990 13302 19992 13354
rect 19936 13300 19992 13302
rect 20040 13354 20096 13356
rect 20040 13302 20042 13354
rect 20042 13302 20094 13354
rect 20094 13302 20096 13354
rect 20040 13300 20096 13302
rect 18396 12962 18452 12964
rect 18396 12910 18398 12962
rect 18398 12910 18450 12962
rect 18450 12910 18452 12962
rect 18396 12908 18452 12910
rect 18284 12796 18340 12852
rect 19404 12908 19460 12964
rect 19068 12850 19124 12852
rect 19068 12798 19070 12850
rect 19070 12798 19122 12850
rect 19122 12798 19124 12850
rect 19068 12796 19124 12798
rect 21644 19234 21700 19236
rect 21644 19182 21646 19234
rect 21646 19182 21698 19234
rect 21698 19182 21700 19234
rect 21644 19180 21700 19182
rect 22204 19068 22260 19124
rect 21308 19010 21364 19012
rect 21308 18958 21310 19010
rect 21310 18958 21362 19010
rect 21362 18958 21364 19010
rect 21308 18956 21364 18958
rect 21196 16882 21252 16884
rect 21196 16830 21198 16882
rect 21198 16830 21250 16882
rect 21250 16830 21252 16882
rect 21196 16828 21252 16830
rect 20972 16604 21028 16660
rect 20860 15596 20916 15652
rect 20636 15484 20692 15540
rect 20524 15426 20580 15428
rect 20524 15374 20526 15426
rect 20526 15374 20578 15426
rect 20578 15374 20580 15426
rect 20524 15372 20580 15374
rect 20636 15260 20692 15316
rect 20412 12908 20468 12964
rect 20748 12850 20804 12852
rect 20748 12798 20750 12850
rect 20750 12798 20802 12850
rect 20802 12798 20804 12850
rect 20748 12796 20804 12798
rect 21420 12796 21476 12852
rect 19292 12290 19348 12292
rect 19292 12238 19294 12290
rect 19294 12238 19346 12290
rect 19346 12238 19348 12290
rect 19292 12236 19348 12238
rect 21644 18450 21700 18452
rect 21644 18398 21646 18450
rect 21646 18398 21698 18450
rect 21698 18398 21700 18450
rect 21644 18396 21700 18398
rect 22492 18842 22548 18844
rect 22492 18790 22494 18842
rect 22494 18790 22546 18842
rect 22546 18790 22548 18842
rect 22492 18788 22548 18790
rect 22596 18842 22652 18844
rect 22596 18790 22598 18842
rect 22598 18790 22650 18842
rect 22650 18790 22652 18842
rect 22596 18788 22652 18790
rect 22700 18842 22756 18844
rect 22700 18790 22702 18842
rect 22702 18790 22754 18842
rect 22754 18790 22756 18842
rect 22700 18788 22756 18790
rect 22204 18450 22260 18452
rect 22204 18398 22206 18450
rect 22206 18398 22258 18450
rect 22258 18398 22260 18450
rect 22204 18396 22260 18398
rect 22492 17274 22548 17276
rect 22492 17222 22494 17274
rect 22494 17222 22546 17274
rect 22546 17222 22548 17274
rect 22492 17220 22548 17222
rect 22596 17274 22652 17276
rect 22596 17222 22598 17274
rect 22598 17222 22650 17274
rect 22650 17222 22652 17274
rect 22596 17220 22652 17222
rect 22700 17274 22756 17276
rect 22700 17222 22702 17274
rect 22702 17222 22754 17274
rect 22754 17222 22756 17274
rect 22700 17220 22756 17222
rect 21644 16940 21700 16996
rect 21644 13634 21700 13636
rect 21644 13582 21646 13634
rect 21646 13582 21698 13634
rect 21698 13582 21700 13634
rect 21644 13580 21700 13582
rect 21868 16156 21924 16212
rect 22316 16210 22372 16212
rect 22316 16158 22318 16210
rect 22318 16158 22370 16210
rect 22370 16158 22372 16210
rect 22316 16156 22372 16158
rect 22492 15706 22548 15708
rect 22492 15654 22494 15706
rect 22494 15654 22546 15706
rect 22546 15654 22548 15706
rect 22492 15652 22548 15654
rect 22596 15706 22652 15708
rect 22596 15654 22598 15706
rect 22598 15654 22650 15706
rect 22650 15654 22652 15706
rect 22596 15652 22652 15654
rect 22700 15706 22756 15708
rect 22700 15654 22702 15706
rect 22702 15654 22754 15706
rect 22754 15654 22756 15706
rect 22700 15652 22756 15654
rect 22492 14138 22548 14140
rect 22492 14086 22494 14138
rect 22494 14086 22546 14138
rect 22546 14086 22548 14138
rect 22492 14084 22548 14086
rect 22596 14138 22652 14140
rect 22596 14086 22598 14138
rect 22598 14086 22650 14138
rect 22650 14086 22652 14138
rect 22596 14084 22652 14086
rect 22700 14138 22756 14140
rect 22700 14086 22702 14138
rect 22702 14086 22754 14138
rect 22754 14086 22756 14138
rect 22700 14084 22756 14086
rect 18508 12124 18564 12180
rect 18396 11954 18452 11956
rect 18396 11902 18398 11954
rect 18398 11902 18450 11954
rect 18450 11902 18452 11954
rect 18396 11900 18452 11902
rect 19180 12178 19236 12180
rect 19180 12126 19182 12178
rect 19182 12126 19234 12178
rect 19234 12126 19236 12178
rect 19180 12124 19236 12126
rect 18172 11228 18228 11284
rect 21084 12460 21140 12516
rect 20412 12236 20468 12292
rect 19628 12178 19684 12180
rect 19628 12126 19630 12178
rect 19630 12126 19682 12178
rect 19682 12126 19684 12178
rect 19628 12124 19684 12126
rect 20300 12178 20356 12180
rect 20300 12126 20302 12178
rect 20302 12126 20354 12178
rect 20354 12126 20356 12178
rect 20300 12124 20356 12126
rect 19832 11786 19888 11788
rect 19832 11734 19834 11786
rect 19834 11734 19886 11786
rect 19886 11734 19888 11786
rect 19832 11732 19888 11734
rect 19936 11786 19992 11788
rect 19936 11734 19938 11786
rect 19938 11734 19990 11786
rect 19990 11734 19992 11786
rect 19936 11732 19992 11734
rect 20040 11786 20096 11788
rect 20040 11734 20042 11786
rect 20042 11734 20094 11786
rect 20094 11734 20096 11786
rect 20040 11732 20096 11734
rect 20748 12402 20804 12404
rect 20748 12350 20750 12402
rect 20750 12350 20802 12402
rect 20802 12350 20804 12402
rect 20748 12348 20804 12350
rect 20412 11900 20468 11956
rect 19404 11116 19460 11172
rect 19852 11340 19908 11396
rect 19180 9884 19236 9940
rect 21196 12348 21252 12404
rect 21644 12460 21700 12516
rect 21644 12290 21700 12292
rect 21644 12238 21646 12290
rect 21646 12238 21698 12290
rect 21698 12238 21700 12290
rect 21644 12236 21700 12238
rect 21084 12178 21140 12180
rect 21084 12126 21086 12178
rect 21086 12126 21138 12178
rect 21138 12126 21140 12178
rect 21084 12124 21140 12126
rect 19832 10218 19888 10220
rect 19832 10166 19834 10218
rect 19834 10166 19886 10218
rect 19886 10166 19888 10218
rect 19832 10164 19888 10166
rect 19936 10218 19992 10220
rect 19936 10166 19938 10218
rect 19938 10166 19990 10218
rect 19990 10166 19992 10218
rect 19936 10164 19992 10166
rect 20040 10218 20096 10220
rect 20040 10166 20042 10218
rect 20042 10166 20094 10218
rect 20094 10166 20096 10218
rect 20040 10164 20096 10166
rect 22204 13580 22260 13636
rect 22204 13244 22260 13300
rect 22492 12570 22548 12572
rect 22492 12518 22494 12570
rect 22494 12518 22546 12570
rect 22546 12518 22548 12570
rect 22492 12516 22548 12518
rect 22596 12570 22652 12572
rect 22596 12518 22598 12570
rect 22598 12518 22650 12570
rect 22650 12518 22652 12570
rect 22596 12516 22652 12518
rect 22700 12570 22756 12572
rect 22700 12518 22702 12570
rect 22702 12518 22754 12570
rect 22754 12518 22756 12570
rect 22700 12516 22756 12518
rect 21980 12124 22036 12180
rect 20972 10668 21028 10724
rect 20188 9884 20244 9940
rect 17836 8316 17892 8372
rect 16604 8258 16660 8260
rect 16604 8206 16606 8258
rect 16606 8206 16658 8258
rect 16658 8206 16660 8258
rect 16604 8204 16660 8206
rect 16380 7868 16436 7924
rect 18060 8092 18116 8148
rect 17172 7866 17228 7868
rect 17172 7814 17174 7866
rect 17174 7814 17226 7866
rect 17226 7814 17228 7866
rect 17172 7812 17228 7814
rect 17276 7866 17332 7868
rect 17276 7814 17278 7866
rect 17278 7814 17330 7866
rect 17330 7814 17332 7866
rect 17276 7812 17332 7814
rect 17380 7866 17436 7868
rect 17380 7814 17382 7866
rect 17382 7814 17434 7866
rect 17434 7814 17436 7866
rect 17380 7812 17436 7814
rect 18284 8092 18340 8148
rect 15708 7420 15764 7476
rect 14512 7082 14568 7084
rect 14512 7030 14514 7082
rect 14514 7030 14566 7082
rect 14566 7030 14568 7082
rect 14512 7028 14568 7030
rect 14616 7082 14672 7084
rect 14616 7030 14618 7082
rect 14618 7030 14670 7082
rect 14670 7030 14672 7082
rect 14616 7028 14672 7030
rect 14720 7082 14776 7084
rect 14720 7030 14722 7082
rect 14722 7030 14774 7082
rect 14774 7030 14776 7082
rect 14720 7028 14776 7030
rect 19068 8146 19124 8148
rect 19068 8094 19070 8146
rect 19070 8094 19122 8146
rect 19122 8094 19124 8146
rect 19068 8092 19124 8094
rect 19964 9826 20020 9828
rect 19964 9774 19966 9826
rect 19966 9774 20018 9826
rect 20018 9774 20020 9826
rect 19964 9772 20020 9774
rect 19628 9714 19684 9716
rect 19628 9662 19630 9714
rect 19630 9662 19682 9714
rect 19682 9662 19684 9714
rect 19628 9660 19684 9662
rect 20076 9714 20132 9716
rect 20076 9662 20078 9714
rect 20078 9662 20130 9714
rect 20130 9662 20132 9714
rect 20076 9660 20132 9662
rect 19832 8650 19888 8652
rect 19832 8598 19834 8650
rect 19834 8598 19886 8650
rect 19886 8598 19888 8650
rect 19832 8596 19888 8598
rect 19936 8650 19992 8652
rect 19936 8598 19938 8650
rect 19938 8598 19990 8650
rect 19990 8598 19992 8650
rect 19936 8596 19992 8598
rect 20040 8650 20096 8652
rect 20040 8598 20042 8650
rect 20042 8598 20094 8650
rect 20094 8598 20096 8650
rect 20040 8596 20096 8598
rect 19740 8258 19796 8260
rect 19740 8206 19742 8258
rect 19742 8206 19794 8258
rect 19794 8206 19796 8258
rect 19740 8204 19796 8206
rect 19404 7698 19460 7700
rect 19404 7646 19406 7698
rect 19406 7646 19458 7698
rect 19458 7646 19460 7698
rect 19404 7644 19460 7646
rect 18956 7586 19012 7588
rect 18956 7534 18958 7586
rect 18958 7534 19010 7586
rect 19010 7534 19012 7586
rect 18956 7532 19012 7534
rect 17948 7308 18004 7364
rect 17724 6524 17780 6580
rect 11340 6412 11396 6468
rect 16044 6466 16100 6468
rect 16044 6414 16046 6466
rect 16046 6414 16098 6466
rect 16098 6414 16100 6466
rect 16044 6412 16100 6414
rect 11852 6298 11908 6300
rect 11852 6246 11854 6298
rect 11854 6246 11906 6298
rect 11906 6246 11908 6298
rect 11852 6244 11908 6246
rect 11956 6298 12012 6300
rect 11956 6246 11958 6298
rect 11958 6246 12010 6298
rect 12010 6246 12012 6298
rect 11956 6244 12012 6246
rect 12060 6298 12116 6300
rect 12060 6246 12062 6298
rect 12062 6246 12114 6298
rect 12114 6246 12116 6298
rect 12060 6244 12116 6246
rect 17172 6298 17228 6300
rect 17172 6246 17174 6298
rect 17174 6246 17226 6298
rect 17226 6246 17228 6298
rect 17172 6244 17228 6246
rect 17276 6298 17332 6300
rect 17276 6246 17278 6298
rect 17278 6246 17330 6298
rect 17330 6246 17332 6298
rect 17276 6244 17332 6246
rect 17380 6298 17436 6300
rect 17380 6246 17382 6298
rect 17382 6246 17434 6298
rect 17434 6246 17436 6298
rect 17380 6244 17436 6246
rect 19180 7474 19236 7476
rect 19180 7422 19182 7474
rect 19182 7422 19234 7474
rect 19234 7422 19236 7474
rect 19180 7420 19236 7422
rect 19068 7362 19124 7364
rect 19068 7310 19070 7362
rect 19070 7310 19122 7362
rect 19122 7310 19124 7362
rect 19068 7308 19124 7310
rect 20524 8258 20580 8260
rect 20524 8206 20526 8258
rect 20526 8206 20578 8258
rect 20578 8206 20580 8258
rect 20524 8204 20580 8206
rect 21420 8146 21476 8148
rect 21420 8094 21422 8146
rect 21422 8094 21474 8146
rect 21474 8094 21476 8146
rect 21420 8092 21476 8094
rect 21308 8034 21364 8036
rect 21308 7982 21310 8034
rect 21310 7982 21362 8034
rect 21362 7982 21364 8034
rect 21308 7980 21364 7982
rect 22492 11002 22548 11004
rect 22492 10950 22494 11002
rect 22494 10950 22546 11002
rect 22546 10950 22548 11002
rect 22492 10948 22548 10950
rect 22596 11002 22652 11004
rect 22596 10950 22598 11002
rect 22598 10950 22650 11002
rect 22650 10950 22652 11002
rect 22596 10948 22652 10950
rect 22700 11002 22756 11004
rect 22700 10950 22702 11002
rect 22702 10950 22754 11002
rect 22754 10950 22756 11002
rect 22700 10948 22756 10950
rect 21868 10722 21924 10724
rect 21868 10670 21870 10722
rect 21870 10670 21922 10722
rect 21922 10670 21924 10722
rect 21868 10668 21924 10670
rect 21644 10332 21700 10388
rect 22204 10332 22260 10388
rect 22492 9434 22548 9436
rect 22492 9382 22494 9434
rect 22494 9382 22546 9434
rect 22546 9382 22548 9434
rect 22492 9380 22548 9382
rect 22596 9434 22652 9436
rect 22596 9382 22598 9434
rect 22598 9382 22650 9434
rect 22650 9382 22652 9434
rect 22596 9380 22652 9382
rect 22700 9434 22756 9436
rect 22700 9382 22702 9434
rect 22702 9382 22754 9434
rect 22754 9382 22756 9434
rect 22700 9380 22756 9382
rect 22876 8204 22932 8260
rect 21868 8146 21924 8148
rect 21868 8094 21870 8146
rect 21870 8094 21922 8146
rect 21922 8094 21924 8146
rect 21868 8092 21924 8094
rect 20188 7586 20244 7588
rect 20188 7534 20190 7586
rect 20190 7534 20242 7586
rect 20242 7534 20244 7586
rect 20188 7532 20244 7534
rect 21308 7644 21364 7700
rect 19964 7420 20020 7476
rect 19832 7082 19888 7084
rect 19832 7030 19834 7082
rect 19834 7030 19886 7082
rect 19886 7030 19888 7082
rect 19832 7028 19888 7030
rect 19936 7082 19992 7084
rect 19936 7030 19938 7082
rect 19938 7030 19990 7082
rect 19990 7030 19992 7082
rect 19936 7028 19992 7030
rect 20040 7082 20096 7084
rect 20040 7030 20042 7082
rect 20042 7030 20094 7082
rect 20094 7030 20096 7082
rect 20040 7028 20096 7030
rect 18284 6524 18340 6580
rect 22492 7866 22548 7868
rect 22492 7814 22494 7866
rect 22494 7814 22546 7866
rect 22546 7814 22548 7866
rect 22492 7812 22548 7814
rect 22596 7866 22652 7868
rect 22596 7814 22598 7866
rect 22598 7814 22650 7866
rect 22650 7814 22652 7866
rect 22596 7812 22652 7814
rect 22700 7866 22756 7868
rect 22700 7814 22702 7866
rect 22702 7814 22754 7866
rect 22754 7814 22756 7866
rect 22700 7812 22756 7814
rect 22204 7474 22260 7476
rect 22204 7422 22206 7474
rect 22206 7422 22258 7474
rect 22258 7422 22260 7474
rect 22204 7420 22260 7422
rect 17836 6466 17892 6468
rect 17836 6414 17838 6466
rect 17838 6414 17890 6466
rect 17890 6414 17892 6466
rect 17836 6412 17892 6414
rect 17948 6076 18004 6132
rect 11228 5964 11284 6020
rect 18508 6130 18564 6132
rect 18508 6078 18510 6130
rect 18510 6078 18562 6130
rect 18562 6078 18564 6130
rect 18508 6076 18564 6078
rect 21532 6076 21588 6132
rect 21868 5964 21924 6020
rect 3872 5514 3928 5516
rect 3872 5462 3874 5514
rect 3874 5462 3926 5514
rect 3926 5462 3928 5514
rect 3872 5460 3928 5462
rect 3976 5514 4032 5516
rect 3976 5462 3978 5514
rect 3978 5462 4030 5514
rect 4030 5462 4032 5514
rect 3976 5460 4032 5462
rect 4080 5514 4136 5516
rect 4080 5462 4082 5514
rect 4082 5462 4134 5514
rect 4134 5462 4136 5514
rect 4080 5460 4136 5462
rect 9192 5514 9248 5516
rect 9192 5462 9194 5514
rect 9194 5462 9246 5514
rect 9246 5462 9248 5514
rect 9192 5460 9248 5462
rect 9296 5514 9352 5516
rect 9296 5462 9298 5514
rect 9298 5462 9350 5514
rect 9350 5462 9352 5514
rect 9296 5460 9352 5462
rect 9400 5514 9456 5516
rect 9400 5462 9402 5514
rect 9402 5462 9454 5514
rect 9454 5462 9456 5514
rect 9400 5460 9456 5462
rect 14512 5514 14568 5516
rect 14512 5462 14514 5514
rect 14514 5462 14566 5514
rect 14566 5462 14568 5514
rect 14512 5460 14568 5462
rect 14616 5514 14672 5516
rect 14616 5462 14618 5514
rect 14618 5462 14670 5514
rect 14670 5462 14672 5514
rect 14616 5460 14672 5462
rect 14720 5514 14776 5516
rect 14720 5462 14722 5514
rect 14722 5462 14774 5514
rect 14774 5462 14776 5514
rect 14720 5460 14776 5462
rect 19832 5514 19888 5516
rect 19832 5462 19834 5514
rect 19834 5462 19886 5514
rect 19886 5462 19888 5514
rect 19832 5460 19888 5462
rect 19936 5514 19992 5516
rect 19936 5462 19938 5514
rect 19938 5462 19990 5514
rect 19990 5462 19992 5514
rect 19936 5460 19992 5462
rect 20040 5514 20096 5516
rect 20040 5462 20042 5514
rect 20042 5462 20094 5514
rect 20094 5462 20096 5514
rect 20040 5460 20096 5462
rect 21644 5122 21700 5124
rect 21644 5070 21646 5122
rect 21646 5070 21698 5122
rect 21698 5070 21700 5122
rect 21644 5068 21700 5070
rect 6532 4730 6588 4732
rect 6532 4678 6534 4730
rect 6534 4678 6586 4730
rect 6586 4678 6588 4730
rect 6532 4676 6588 4678
rect 6636 4730 6692 4732
rect 6636 4678 6638 4730
rect 6638 4678 6690 4730
rect 6690 4678 6692 4730
rect 6636 4676 6692 4678
rect 6740 4730 6796 4732
rect 6740 4678 6742 4730
rect 6742 4678 6794 4730
rect 6794 4678 6796 4730
rect 6740 4676 6796 4678
rect 11852 4730 11908 4732
rect 11852 4678 11854 4730
rect 11854 4678 11906 4730
rect 11906 4678 11908 4730
rect 11852 4676 11908 4678
rect 11956 4730 12012 4732
rect 11956 4678 11958 4730
rect 11958 4678 12010 4730
rect 12010 4678 12012 4730
rect 11956 4676 12012 4678
rect 12060 4730 12116 4732
rect 12060 4678 12062 4730
rect 12062 4678 12114 4730
rect 12114 4678 12116 4730
rect 12060 4676 12116 4678
rect 17172 4730 17228 4732
rect 17172 4678 17174 4730
rect 17174 4678 17226 4730
rect 17226 4678 17228 4730
rect 17172 4676 17228 4678
rect 17276 4730 17332 4732
rect 17276 4678 17278 4730
rect 17278 4678 17330 4730
rect 17330 4678 17332 4730
rect 17276 4676 17332 4678
rect 17380 4730 17436 4732
rect 17380 4678 17382 4730
rect 17382 4678 17434 4730
rect 17434 4678 17436 4730
rect 17380 4676 17436 4678
rect 3872 3946 3928 3948
rect 3872 3894 3874 3946
rect 3874 3894 3926 3946
rect 3926 3894 3928 3946
rect 3872 3892 3928 3894
rect 3976 3946 4032 3948
rect 3976 3894 3978 3946
rect 3978 3894 4030 3946
rect 4030 3894 4032 3946
rect 3976 3892 4032 3894
rect 4080 3946 4136 3948
rect 4080 3894 4082 3946
rect 4082 3894 4134 3946
rect 4134 3894 4136 3946
rect 4080 3892 4136 3894
rect 9192 3946 9248 3948
rect 9192 3894 9194 3946
rect 9194 3894 9246 3946
rect 9246 3894 9248 3946
rect 9192 3892 9248 3894
rect 9296 3946 9352 3948
rect 9296 3894 9298 3946
rect 9298 3894 9350 3946
rect 9350 3894 9352 3946
rect 9296 3892 9352 3894
rect 9400 3946 9456 3948
rect 9400 3894 9402 3946
rect 9402 3894 9454 3946
rect 9454 3894 9456 3946
rect 9400 3892 9456 3894
rect 14512 3946 14568 3948
rect 14512 3894 14514 3946
rect 14514 3894 14566 3946
rect 14566 3894 14568 3946
rect 14512 3892 14568 3894
rect 14616 3946 14672 3948
rect 14616 3894 14618 3946
rect 14618 3894 14670 3946
rect 14670 3894 14672 3946
rect 14616 3892 14672 3894
rect 14720 3946 14776 3948
rect 14720 3894 14722 3946
rect 14722 3894 14774 3946
rect 14774 3894 14776 3946
rect 14720 3892 14776 3894
rect 19832 3946 19888 3948
rect 19832 3894 19834 3946
rect 19834 3894 19886 3946
rect 19886 3894 19888 3946
rect 19832 3892 19888 3894
rect 19936 3946 19992 3948
rect 19936 3894 19938 3946
rect 19938 3894 19990 3946
rect 19990 3894 19992 3946
rect 19936 3892 19992 3894
rect 20040 3946 20096 3948
rect 20040 3894 20042 3946
rect 20042 3894 20094 3946
rect 20094 3894 20096 3946
rect 20040 3892 20096 3894
rect 6532 3162 6588 3164
rect 6532 3110 6534 3162
rect 6534 3110 6586 3162
rect 6586 3110 6588 3162
rect 6532 3108 6588 3110
rect 6636 3162 6692 3164
rect 6636 3110 6638 3162
rect 6638 3110 6690 3162
rect 6690 3110 6692 3162
rect 6636 3108 6692 3110
rect 6740 3162 6796 3164
rect 6740 3110 6742 3162
rect 6742 3110 6794 3162
rect 6794 3110 6796 3162
rect 6740 3108 6796 3110
rect 11852 3162 11908 3164
rect 11852 3110 11854 3162
rect 11854 3110 11906 3162
rect 11906 3110 11908 3162
rect 11852 3108 11908 3110
rect 11956 3162 12012 3164
rect 11956 3110 11958 3162
rect 11958 3110 12010 3162
rect 12010 3110 12012 3162
rect 11956 3108 12012 3110
rect 12060 3162 12116 3164
rect 12060 3110 12062 3162
rect 12062 3110 12114 3162
rect 12114 3110 12116 3162
rect 12060 3108 12116 3110
rect 17172 3162 17228 3164
rect 17172 3110 17174 3162
rect 17174 3110 17226 3162
rect 17226 3110 17228 3162
rect 17172 3108 17228 3110
rect 17276 3162 17332 3164
rect 17276 3110 17278 3162
rect 17278 3110 17330 3162
rect 17330 3110 17332 3162
rect 17276 3108 17332 3110
rect 17380 3162 17436 3164
rect 17380 3110 17382 3162
rect 17382 3110 17434 3162
rect 17434 3110 17436 3162
rect 17380 3108 17436 3110
rect 22492 6298 22548 6300
rect 22492 6246 22494 6298
rect 22494 6246 22546 6298
rect 22546 6246 22548 6298
rect 22492 6244 22548 6246
rect 22596 6298 22652 6300
rect 22596 6246 22598 6298
rect 22598 6246 22650 6298
rect 22650 6246 22652 6298
rect 22596 6244 22652 6246
rect 22700 6298 22756 6300
rect 22700 6246 22702 6298
rect 22702 6246 22754 6298
rect 22754 6246 22756 6298
rect 22700 6244 22756 6246
rect 22204 5122 22260 5124
rect 22204 5070 22206 5122
rect 22206 5070 22258 5122
rect 22258 5070 22260 5122
rect 22204 5068 22260 5070
rect 22492 4730 22548 4732
rect 22492 4678 22494 4730
rect 22494 4678 22546 4730
rect 22546 4678 22548 4730
rect 22492 4676 22548 4678
rect 22596 4730 22652 4732
rect 22596 4678 22598 4730
rect 22598 4678 22650 4730
rect 22650 4678 22652 4730
rect 22596 4676 22652 4678
rect 22700 4730 22756 4732
rect 22700 4678 22702 4730
rect 22702 4678 22754 4730
rect 22754 4678 22756 4730
rect 22700 4676 22756 4678
rect 22204 4508 22260 4564
rect 22492 3162 22548 3164
rect 22492 3110 22494 3162
rect 22494 3110 22546 3162
rect 22546 3110 22548 3162
rect 22492 3108 22548 3110
rect 22596 3162 22652 3164
rect 22596 3110 22598 3162
rect 22598 3110 22650 3162
rect 22650 3110 22652 3162
rect 22596 3108 22652 3110
rect 22700 3162 22756 3164
rect 22700 3110 22702 3162
rect 22702 3110 22754 3162
rect 22754 3110 22756 3162
rect 22700 3108 22756 3110
rect 22092 1596 22148 1652
<< metal3 >>
rect 23200 22036 24000 22064
rect 20066 21980 20076 22036
rect 20132 21980 24000 22036
rect 23200 21952 24000 21980
rect 6522 20356 6532 20412
rect 6588 20356 6636 20412
rect 6692 20356 6740 20412
rect 6796 20356 6806 20412
rect 11842 20356 11852 20412
rect 11908 20356 11956 20412
rect 12012 20356 12060 20412
rect 12116 20356 12126 20412
rect 17162 20356 17172 20412
rect 17228 20356 17276 20412
rect 17332 20356 17380 20412
rect 17436 20356 17446 20412
rect 22482 20356 22492 20412
rect 22548 20356 22596 20412
rect 22652 20356 22700 20412
rect 22756 20356 22766 20412
rect 19730 20076 19740 20132
rect 19796 20076 20748 20132
rect 20804 20076 20814 20132
rect 13570 19964 13580 20020
rect 13636 19964 18508 20020
rect 18564 19964 18574 20020
rect 11330 19852 11340 19908
rect 11396 19852 19852 19908
rect 19908 19852 19918 19908
rect 13682 19740 13692 19796
rect 13748 19740 17948 19796
rect 18004 19740 18014 19796
rect 3862 19572 3872 19628
rect 3928 19572 3976 19628
rect 4032 19572 4080 19628
rect 4136 19572 4146 19628
rect 9182 19572 9192 19628
rect 9248 19572 9296 19628
rect 9352 19572 9400 19628
rect 9456 19572 9466 19628
rect 14502 19572 14512 19628
rect 14568 19572 14616 19628
rect 14672 19572 14720 19628
rect 14776 19572 14786 19628
rect 19822 19572 19832 19628
rect 19888 19572 19936 19628
rect 19992 19572 20040 19628
rect 20096 19572 20106 19628
rect 3042 19180 3052 19236
rect 3108 19180 4172 19236
rect 4228 19180 6748 19236
rect 6804 19180 6814 19236
rect 11666 19180 11676 19236
rect 11732 19180 13468 19236
rect 13524 19180 13534 19236
rect 17938 19180 17948 19236
rect 18004 19180 19292 19236
rect 19348 19180 19358 19236
rect 20626 19180 20636 19236
rect 20692 19180 21644 19236
rect 21700 19180 21710 19236
rect 23200 19124 24000 19152
rect 4610 19068 4620 19124
rect 4676 19068 10780 19124
rect 10836 19068 10846 19124
rect 18386 19068 18396 19124
rect 18452 19068 19180 19124
rect 19236 19068 19246 19124
rect 22194 19068 22204 19124
rect 22260 19068 24000 19124
rect 23200 19040 24000 19068
rect 6626 18956 6636 19012
rect 6692 18956 7084 19012
rect 7140 18956 7150 19012
rect 7410 18956 7420 19012
rect 7476 18956 7980 19012
rect 8036 18956 9548 19012
rect 9604 18956 9614 19012
rect 19394 18956 19404 19012
rect 19460 18956 21308 19012
rect 21364 18956 21374 19012
rect 6522 18788 6532 18844
rect 6588 18788 6636 18844
rect 6692 18788 6740 18844
rect 6796 18788 6806 18844
rect 11842 18788 11852 18844
rect 11908 18788 11956 18844
rect 12012 18788 12060 18844
rect 12116 18788 12126 18844
rect 17162 18788 17172 18844
rect 17228 18788 17276 18844
rect 17332 18788 17380 18844
rect 17436 18788 17446 18844
rect 22482 18788 22492 18844
rect 22548 18788 22596 18844
rect 22652 18788 22700 18844
rect 22756 18788 22766 18844
rect 10882 18620 10892 18676
rect 10948 18620 13692 18676
rect 13748 18620 14028 18676
rect 14084 18620 14094 18676
rect 3154 18508 3164 18564
rect 3220 18508 3836 18564
rect 3892 18508 3902 18564
rect 5954 18396 5964 18452
rect 6020 18396 6972 18452
rect 7028 18396 7644 18452
rect 7700 18396 7710 18452
rect 13234 18396 13244 18452
rect 13300 18396 14140 18452
rect 14196 18396 14206 18452
rect 14354 18396 14364 18452
rect 14420 18396 15596 18452
rect 15652 18396 16044 18452
rect 16100 18396 16110 18452
rect 21634 18396 21644 18452
rect 21700 18396 22204 18452
rect 22260 18396 22270 18452
rect 6850 18284 6860 18340
rect 6916 18284 10892 18340
rect 10948 18284 11228 18340
rect 11284 18284 11294 18340
rect 11666 18284 11676 18340
rect 11732 18284 15932 18340
rect 15988 18284 16268 18340
rect 16324 18284 16334 18340
rect 3378 18172 3388 18228
rect 3444 18172 5068 18228
rect 5124 18172 7868 18228
rect 7924 18172 8428 18228
rect 8484 18172 16604 18228
rect 16660 18172 19516 18228
rect 19572 18172 19582 18228
rect 3862 18004 3872 18060
rect 3928 18004 3976 18060
rect 4032 18004 4080 18060
rect 4136 18004 4146 18060
rect 9182 18004 9192 18060
rect 9248 18004 9296 18060
rect 9352 18004 9400 18060
rect 9456 18004 9466 18060
rect 14502 18004 14512 18060
rect 14568 18004 14616 18060
rect 14672 18004 14720 18060
rect 14776 18004 14786 18060
rect 19822 18004 19832 18060
rect 19888 18004 19936 18060
rect 19992 18004 20040 18060
rect 20096 18004 20106 18060
rect 3042 17836 3052 17892
rect 3108 17836 3556 17892
rect 19842 17836 19852 17892
rect 19908 17836 20636 17892
rect 20692 17836 20702 17892
rect 3500 17668 3556 17836
rect 19506 17724 19516 17780
rect 19572 17724 19964 17780
rect 20020 17724 20030 17780
rect 3490 17612 3500 17668
rect 3556 17612 3566 17668
rect 11106 17500 11116 17556
rect 11172 17500 11564 17556
rect 11620 17500 11630 17556
rect 3154 17388 3164 17444
rect 3220 17388 4620 17444
rect 4676 17388 4686 17444
rect 6626 17388 6636 17444
rect 6692 17388 8428 17444
rect 8484 17388 8494 17444
rect 9538 17388 9548 17444
rect 9604 17388 10332 17444
rect 10388 17388 10668 17444
rect 10724 17388 11228 17444
rect 11284 17388 11294 17444
rect 6522 17220 6532 17276
rect 6588 17220 6636 17276
rect 6692 17220 6740 17276
rect 6796 17220 6806 17276
rect 11842 17220 11852 17276
rect 11908 17220 11956 17276
rect 12012 17220 12060 17276
rect 12116 17220 12126 17276
rect 17162 17220 17172 17276
rect 17228 17220 17276 17276
rect 17332 17220 17380 17276
rect 17436 17220 17446 17276
rect 22482 17220 22492 17276
rect 22548 17220 22596 17276
rect 22652 17220 22700 17276
rect 22756 17220 22766 17276
rect 9650 16940 9660 16996
rect 9716 16940 9726 16996
rect 10882 16940 10892 16996
rect 10948 16940 11788 16996
rect 11844 16940 13132 16996
rect 13188 16940 13198 16996
rect 20514 16940 20524 16996
rect 20580 16940 21644 16996
rect 21700 16940 21710 16996
rect 9660 16772 9716 16940
rect 8866 16716 8876 16772
rect 8932 16716 9716 16772
rect 9772 16828 11004 16884
rect 11060 16828 11070 16884
rect 11330 16828 11340 16884
rect 11396 16828 12236 16884
rect 12292 16828 12302 16884
rect 19394 16828 19404 16884
rect 19460 16828 20188 16884
rect 20244 16828 21196 16884
rect 21252 16828 21262 16884
rect 9772 16548 9828 16828
rect 10434 16716 10444 16772
rect 10500 16716 11452 16772
rect 11508 16716 11518 16772
rect 19730 16604 19740 16660
rect 19796 16604 20300 16660
rect 20356 16604 20972 16660
rect 21028 16604 21038 16660
rect 9762 16492 9772 16548
rect 9828 16492 9838 16548
rect 3862 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4146 16492
rect 9182 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9466 16492
rect 14502 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14786 16492
rect 19822 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20106 16492
rect 4386 16268 4396 16324
rect 4452 16268 4844 16324
rect 4900 16268 5292 16324
rect 5348 16268 15036 16324
rect 15092 16268 15102 16324
rect 15474 16268 15484 16324
rect 15540 16268 15932 16324
rect 15988 16268 19740 16324
rect 19796 16268 19806 16324
rect 23200 16212 24000 16240
rect 19618 16156 19628 16212
rect 19684 16156 21868 16212
rect 21924 16156 21934 16212
rect 22306 16156 22316 16212
rect 22372 16156 24000 16212
rect 23200 16128 24000 16156
rect 2930 16044 2940 16100
rect 2996 16044 4620 16100
rect 4676 16044 8876 16100
rect 8932 16044 8942 16100
rect 14130 16044 14140 16100
rect 14196 16044 14924 16100
rect 14980 16044 19180 16100
rect 19236 16044 19246 16100
rect 6522 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6806 15708
rect 11842 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12126 15708
rect 17162 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17446 15708
rect 22482 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22766 15708
rect 20850 15596 20860 15652
rect 20916 15596 20926 15652
rect 19954 15484 19964 15540
rect 20020 15484 20636 15540
rect 20692 15484 20702 15540
rect 11442 15372 11452 15428
rect 11508 15372 14476 15428
rect 14532 15372 14542 15428
rect 19730 15372 19740 15428
rect 19796 15372 20524 15428
rect 20580 15372 20590 15428
rect 20860 15316 20916 15596
rect 18834 15260 18844 15316
rect 18900 15260 19516 15316
rect 19572 15260 20300 15316
rect 20356 15260 20366 15316
rect 20626 15260 20636 15316
rect 20692 15260 20916 15316
rect 9986 15148 9996 15204
rect 10052 15148 11004 15204
rect 11060 15148 11070 15204
rect 15026 15148 15036 15204
rect 15092 15148 17612 15204
rect 17668 15148 17678 15204
rect 17826 15148 17836 15204
rect 17892 15148 19740 15204
rect 19796 15148 19806 15204
rect 15810 15036 15820 15092
rect 15876 15036 17948 15092
rect 18004 15036 18014 15092
rect 15474 14924 15484 14980
rect 15540 14924 16044 14980
rect 16100 14924 16940 14980
rect 16996 14924 17006 14980
rect 3862 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4146 14924
rect 9182 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9466 14924
rect 14502 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14786 14924
rect 19822 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20106 14924
rect 3602 14476 3612 14532
rect 3668 14476 4844 14532
rect 4900 14476 4910 14532
rect 9090 14476 9100 14532
rect 9156 14476 9772 14532
rect 9828 14476 9838 14532
rect 13794 14476 13804 14532
rect 13860 14476 14700 14532
rect 14756 14476 14766 14532
rect 15092 14476 15372 14532
rect 15428 14476 15438 14532
rect 15092 14420 15148 14476
rect 3332 14364 4620 14420
rect 4676 14364 6076 14420
rect 6132 14364 8652 14420
rect 8708 14364 8718 14420
rect 14130 14364 14140 14420
rect 14196 14364 15148 14420
rect 3332 14196 3388 14364
rect 3826 14252 3836 14308
rect 3892 14252 3902 14308
rect 4162 14252 4172 14308
rect 4228 14252 4564 14308
rect 8866 14252 8876 14308
rect 8932 14252 10892 14308
rect 10948 14252 10958 14308
rect 14466 14252 14476 14308
rect 14532 14252 15036 14308
rect 15092 14252 15708 14308
rect 15764 14252 15774 14308
rect 3042 14140 3052 14196
rect 3108 14140 3388 14196
rect 3836 13860 3892 14252
rect 4508 14196 4564 14252
rect 4498 14140 4508 14196
rect 4564 14140 4574 14196
rect 6522 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6806 14140
rect 11842 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12126 14140
rect 17162 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17446 14140
rect 22482 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22766 14140
rect 9650 13916 9660 13972
rect 9716 13916 19180 13972
rect 19236 13916 19246 13972
rect 3490 13804 3500 13860
rect 3556 13804 3892 13860
rect 2370 13692 2380 13748
rect 2436 13692 3052 13748
rect 3108 13692 3118 13748
rect 4246 13692 4284 13748
rect 4340 13692 4350 13748
rect 5394 13580 5404 13636
rect 5460 13580 6188 13636
rect 6244 13580 9100 13636
rect 9156 13580 9884 13636
rect 9940 13580 9950 13636
rect 21634 13580 21644 13636
rect 21700 13580 22204 13636
rect 22260 13580 22270 13636
rect 4284 13468 4732 13524
rect 4788 13468 5516 13524
rect 5572 13468 5582 13524
rect 10210 13468 10220 13524
rect 10276 13468 12236 13524
rect 12292 13468 14140 13524
rect 14196 13468 14206 13524
rect 3862 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4146 13356
rect 4284 13188 4340 13468
rect 10546 13356 10556 13412
rect 10612 13356 11116 13412
rect 11172 13356 11182 13412
rect 14914 13356 14924 13412
rect 14980 13356 17500 13412
rect 17556 13356 18284 13412
rect 18340 13356 18350 13412
rect 9182 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9466 13356
rect 14502 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14786 13356
rect 19822 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20106 13356
rect 23200 13300 24000 13328
rect 22194 13244 22204 13300
rect 22260 13244 24000 13300
rect 23200 13216 24000 13244
rect 4162 13132 4172 13188
rect 4228 13132 4340 13188
rect 14242 13132 14252 13188
rect 14308 13132 14588 13188
rect 14644 13132 15372 13188
rect 15428 13132 15438 13188
rect 10434 12908 10444 12964
rect 10500 12908 11452 12964
rect 11508 12908 11518 12964
rect 15922 12908 15932 12964
rect 15988 12908 18396 12964
rect 18452 12908 18462 12964
rect 19394 12908 19404 12964
rect 19460 12908 20412 12964
rect 20468 12908 20478 12964
rect 4946 12796 4956 12852
rect 5012 12796 14476 12852
rect 14532 12796 14542 12852
rect 15932 12740 15988 12908
rect 18274 12796 18284 12852
rect 18340 12796 19068 12852
rect 19124 12796 19134 12852
rect 20738 12796 20748 12852
rect 20804 12796 21420 12852
rect 21476 12796 21486 12852
rect 8530 12684 8540 12740
rect 8596 12684 9212 12740
rect 9268 12684 9278 12740
rect 15138 12684 15148 12740
rect 15204 12684 15988 12740
rect 4386 12572 4396 12628
rect 4452 12572 4462 12628
rect 4396 12404 4452 12572
rect 6522 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6806 12572
rect 11842 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12126 12572
rect 17162 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17446 12572
rect 22482 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22766 12572
rect 9986 12460 9996 12516
rect 10052 12460 10444 12516
rect 10500 12460 10510 12516
rect 21074 12460 21084 12516
rect 21140 12460 21644 12516
rect 21700 12460 21710 12516
rect 4358 12348 4396 12404
rect 4452 12348 4620 12404
rect 4676 12348 4686 12404
rect 20738 12348 20748 12404
rect 20804 12348 21196 12404
rect 21252 12348 21262 12404
rect 4274 12236 4284 12292
rect 4340 12236 4508 12292
rect 4564 12236 4574 12292
rect 15362 12236 15372 12292
rect 15428 12236 16268 12292
rect 16324 12236 19292 12292
rect 19348 12236 19358 12292
rect 20402 12236 20412 12292
rect 20468 12236 21644 12292
rect 21700 12236 21710 12292
rect 4274 12124 4284 12180
rect 4340 12124 4620 12180
rect 4676 12124 4686 12180
rect 9986 12124 9996 12180
rect 10052 12124 10444 12180
rect 10500 12124 15260 12180
rect 15316 12124 16156 12180
rect 16212 12124 16222 12180
rect 17154 12124 17164 12180
rect 17220 12124 18060 12180
rect 18116 12124 18126 12180
rect 18498 12124 18508 12180
rect 18564 12124 19180 12180
rect 19236 12124 19246 12180
rect 19618 12124 19628 12180
rect 19684 12124 20300 12180
rect 20356 12124 20366 12180
rect 21074 12124 21084 12180
rect 21140 12124 21980 12180
rect 22036 12124 22046 12180
rect 10770 12012 10780 12068
rect 10836 12012 11340 12068
rect 11396 12012 13804 12068
rect 13860 12012 13870 12068
rect 8642 11900 8652 11956
rect 8708 11900 10892 11956
rect 10948 11900 11228 11956
rect 11284 11900 11294 11956
rect 18386 11900 18396 11956
rect 18452 11900 20412 11956
rect 20468 11900 20478 11956
rect 9762 11788 9772 11844
rect 9828 11788 10612 11844
rect 3862 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4146 11788
rect 9182 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9466 11788
rect 10556 11620 10612 11788
rect 14502 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14786 11788
rect 19822 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20106 11788
rect 11554 11676 11564 11732
rect 11620 11676 12572 11732
rect 12628 11676 13692 11732
rect 13748 11676 13758 11732
rect 14914 11676 14924 11732
rect 14980 11676 16156 11732
rect 16212 11676 17388 11732
rect 17444 11676 17454 11732
rect 10546 11564 10556 11620
rect 10612 11564 11676 11620
rect 11732 11564 17052 11620
rect 17108 11564 17118 11620
rect 13682 11452 13692 11508
rect 13748 11452 15484 11508
rect 15540 11452 15550 11508
rect 15810 11452 15820 11508
rect 15876 11452 17948 11508
rect 18004 11452 18014 11508
rect 3154 11340 3164 11396
rect 3220 11340 3612 11396
rect 3668 11340 3678 11396
rect 17602 11340 17612 11396
rect 17668 11340 19852 11396
rect 19908 11340 19918 11396
rect 10322 11228 10332 11284
rect 10388 11228 13468 11284
rect 13524 11228 13860 11284
rect 14242 11228 14252 11284
rect 14308 11228 14924 11284
rect 14980 11228 16492 11284
rect 16548 11228 18172 11284
rect 18228 11228 18238 11284
rect 13804 11172 13860 11228
rect 10770 11116 10780 11172
rect 10836 11116 13580 11172
rect 13636 11116 13646 11172
rect 13804 11116 19404 11172
rect 19460 11116 19470 11172
rect 3378 11004 3388 11060
rect 3444 11004 3454 11060
rect 15026 11004 15036 11060
rect 15092 11004 15260 11060
rect 15316 11004 15326 11060
rect 3388 10948 3444 11004
rect 6522 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6806 11004
rect 11842 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12126 11004
rect 17162 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17446 11004
rect 22482 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22766 11004
rect 3388 10892 3612 10948
rect 3668 10892 3678 10948
rect 3266 10780 3276 10836
rect 3332 10780 4284 10836
rect 4340 10780 4350 10836
rect 8530 10780 8540 10836
rect 8596 10780 9548 10836
rect 9604 10780 9614 10836
rect 12450 10780 12460 10836
rect 12516 10780 14476 10836
rect 14532 10780 15148 10836
rect 2930 10668 2940 10724
rect 2996 10668 3724 10724
rect 3780 10668 3790 10724
rect 15092 10500 15148 10780
rect 20962 10668 20972 10724
rect 21028 10668 21868 10724
rect 21924 10668 21934 10724
rect 15092 10444 15316 10500
rect 15260 10388 15316 10444
rect 23200 10388 24000 10416
rect 15250 10332 15260 10388
rect 15316 10332 15326 10388
rect 21634 10332 21644 10388
rect 21700 10332 22204 10388
rect 22260 10332 24000 10388
rect 23200 10304 24000 10332
rect 3862 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4146 10220
rect 9182 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9466 10220
rect 14502 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14786 10220
rect 19822 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20106 10220
rect 9548 10108 9772 10164
rect 9828 10108 12572 10164
rect 12628 10108 12638 10164
rect 9548 10052 9604 10108
rect 3154 9996 3164 10052
rect 3220 9996 3836 10052
rect 3892 9996 3902 10052
rect 9314 9996 9324 10052
rect 9380 9996 9604 10052
rect 19170 9884 19180 9940
rect 19236 9884 20188 9940
rect 20244 9884 20254 9940
rect 3378 9772 3388 9828
rect 3444 9772 4508 9828
rect 4564 9772 4574 9828
rect 9874 9772 9884 9828
rect 9940 9772 10332 9828
rect 10388 9772 10398 9828
rect 15586 9772 15596 9828
rect 15652 9772 19964 9828
rect 20020 9772 20030 9828
rect 3126 9660 3164 9716
rect 3220 9660 3230 9716
rect 9538 9660 9548 9716
rect 9604 9660 10444 9716
rect 10500 9660 10510 9716
rect 19618 9660 19628 9716
rect 19684 9660 20076 9716
rect 20132 9660 20142 9716
rect 5058 9548 5068 9604
rect 5124 9548 5740 9604
rect 5796 9548 5806 9604
rect 6522 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6806 9436
rect 11842 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12126 9436
rect 17162 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17446 9436
rect 22482 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22766 9436
rect 4834 9212 4844 9268
rect 4900 9212 5964 9268
rect 6020 9212 6030 9268
rect 3332 9100 3948 9156
rect 4004 9100 9996 9156
rect 10052 9100 10062 9156
rect 3332 8820 3388 9100
rect 3602 8988 3612 9044
rect 3668 8988 4956 9044
rect 5012 8988 5022 9044
rect 6514 8988 6524 9044
rect 6580 8988 11116 9044
rect 11172 8988 11182 9044
rect 5058 8876 5068 8932
rect 5124 8876 5516 8932
rect 5572 8876 5582 8932
rect 6066 8876 6076 8932
rect 6132 8876 10668 8932
rect 10724 8876 10734 8932
rect 3042 8764 3052 8820
rect 3108 8764 3388 8820
rect 4162 8764 4172 8820
rect 4228 8764 6188 8820
rect 6244 8764 9436 8820
rect 9492 8764 9502 8820
rect 10098 8764 10108 8820
rect 10164 8764 10332 8820
rect 10388 8764 14252 8820
rect 14308 8764 14318 8820
rect 10434 8652 10444 8708
rect 10500 8652 11004 8708
rect 11060 8652 11070 8708
rect 3862 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4146 8652
rect 9182 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9466 8652
rect 14502 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14786 8652
rect 19822 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20106 8652
rect 4498 8540 4508 8596
rect 4564 8540 6076 8596
rect 6132 8540 6142 8596
rect 5954 8428 5964 8484
rect 6020 8428 10108 8484
rect 10164 8428 10174 8484
rect 10434 8428 10444 8484
rect 10500 8428 14364 8484
rect 14420 8428 14430 8484
rect 8978 8316 8988 8372
rect 9044 8316 9884 8372
rect 9940 8316 10668 8372
rect 10724 8316 11340 8372
rect 11396 8316 11406 8372
rect 15372 8316 17836 8372
rect 17892 8316 17902 8372
rect 15372 8260 15428 8316
rect 5058 8204 5068 8260
rect 5124 8204 5740 8260
rect 5796 8204 5806 8260
rect 9650 8204 9660 8260
rect 9716 8204 10332 8260
rect 10388 8204 10398 8260
rect 11554 8204 11564 8260
rect 11620 8204 15148 8260
rect 15362 8204 15372 8260
rect 15428 8204 15438 8260
rect 16258 8204 16268 8260
rect 16324 8204 16334 8260
rect 16594 8204 16604 8260
rect 16660 8204 19740 8260
rect 19796 8204 19806 8260
rect 20514 8204 20524 8260
rect 20580 8204 22876 8260
rect 22932 8204 22942 8260
rect 15092 8148 15148 8204
rect 16268 8148 16324 8204
rect 3154 8092 3164 8148
rect 3220 8092 6076 8148
rect 6132 8092 7028 8148
rect 10210 8092 10220 8148
rect 10276 8092 11004 8148
rect 11060 8092 11070 8148
rect 15092 8092 15484 8148
rect 15540 8092 15550 8148
rect 16268 8092 18060 8148
rect 18116 8092 18126 8148
rect 18274 8092 18284 8148
rect 18340 8092 19068 8148
rect 19124 8092 19134 8148
rect 21410 8092 21420 8148
rect 21476 8092 21868 8148
rect 21924 8092 21934 8148
rect 6972 7924 7028 8092
rect 10098 7980 10108 8036
rect 10164 7980 10668 8036
rect 10724 7980 11116 8036
rect 11172 7980 14588 8036
rect 14644 7980 16268 8036
rect 16324 7980 16334 8036
rect 21298 7980 21308 8036
rect 21364 7980 21374 8036
rect 6972 7868 11004 7924
rect 11060 7868 11070 7924
rect 6522 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6806 7868
rect 11842 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12126 7868
rect 15092 7700 15148 7924
rect 15204 7868 16380 7924
rect 16436 7868 16446 7924
rect 17162 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17446 7868
rect 21308 7812 21364 7980
rect 22482 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22766 7868
rect 11778 7644 11788 7700
rect 11844 7644 15148 7700
rect 18284 7756 21364 7812
rect 18284 7588 18340 7756
rect 19394 7644 19404 7700
rect 19460 7644 21308 7700
rect 21364 7644 21374 7700
rect 11330 7532 11340 7588
rect 11396 7532 18340 7588
rect 18946 7532 18956 7588
rect 19012 7532 20188 7588
rect 20244 7532 20254 7588
rect 23200 7476 24000 7504
rect 15698 7420 15708 7476
rect 15764 7420 19180 7476
rect 19236 7420 19964 7476
rect 20020 7420 20030 7476
rect 22194 7420 22204 7476
rect 22260 7420 24000 7476
rect 23200 7392 24000 7420
rect 4946 7308 4956 7364
rect 5012 7308 5628 7364
rect 5684 7308 9660 7364
rect 9716 7308 9726 7364
rect 17938 7308 17948 7364
rect 18004 7308 19068 7364
rect 19124 7308 19134 7364
rect 3862 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4146 7084
rect 9182 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9466 7084
rect 14502 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14786 7084
rect 19822 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20106 7084
rect 4834 6972 4844 7028
rect 4900 6972 5628 7028
rect 5684 6972 5694 7028
rect 9426 6860 9436 6916
rect 9492 6860 9996 6916
rect 10052 6860 10062 6916
rect 10322 6860 10332 6916
rect 10388 6860 10892 6916
rect 10948 6860 10958 6916
rect 4834 6748 4844 6804
rect 4900 6748 5740 6804
rect 5796 6748 5806 6804
rect 10210 6636 10220 6692
rect 10276 6636 11452 6692
rect 11508 6636 11518 6692
rect 5954 6524 5964 6580
rect 6020 6524 6412 6580
rect 6468 6524 17724 6580
rect 17780 6524 18284 6580
rect 18340 6524 18350 6580
rect 10882 6412 10892 6468
rect 10948 6412 11340 6468
rect 11396 6412 16044 6468
rect 16100 6412 17836 6468
rect 17892 6412 17902 6468
rect 6522 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6806 6300
rect 11842 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12126 6300
rect 17162 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17446 6300
rect 22482 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22766 6300
rect 8530 6076 8540 6132
rect 8596 6076 17948 6132
rect 18004 6076 18508 6132
rect 18564 6076 21532 6132
rect 21588 6076 21598 6132
rect 9874 5964 9884 6020
rect 9940 5964 10332 6020
rect 10388 5964 11228 6020
rect 11284 5964 21868 6020
rect 21924 5964 21934 6020
rect 3862 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4146 5516
rect 9182 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9466 5516
rect 14502 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14786 5516
rect 19822 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20106 5516
rect 21634 5068 21644 5124
rect 21700 5068 22204 5124
rect 22260 5068 22270 5124
rect 6522 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6806 4732
rect 11842 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12126 4732
rect 17162 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17446 4732
rect 22482 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22766 4732
rect 23200 4564 24000 4592
rect 22194 4508 22204 4564
rect 22260 4508 24000 4564
rect 23200 4480 24000 4508
rect 3862 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4146 3948
rect 9182 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9466 3948
rect 14502 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14786 3948
rect 19822 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20106 3948
rect 6522 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6806 3164
rect 11842 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12126 3164
rect 17162 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17446 3164
rect 22482 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22766 3164
rect 23200 1652 24000 1680
rect 22082 1596 22092 1652
rect 22148 1596 24000 1652
rect 23200 1568 24000 1596
<< via3 >>
rect 6532 20356 6588 20412
rect 6636 20356 6692 20412
rect 6740 20356 6796 20412
rect 11852 20356 11908 20412
rect 11956 20356 12012 20412
rect 12060 20356 12116 20412
rect 17172 20356 17228 20412
rect 17276 20356 17332 20412
rect 17380 20356 17436 20412
rect 22492 20356 22548 20412
rect 22596 20356 22652 20412
rect 22700 20356 22756 20412
rect 3872 19572 3928 19628
rect 3976 19572 4032 19628
rect 4080 19572 4136 19628
rect 9192 19572 9248 19628
rect 9296 19572 9352 19628
rect 9400 19572 9456 19628
rect 14512 19572 14568 19628
rect 14616 19572 14672 19628
rect 14720 19572 14776 19628
rect 19832 19572 19888 19628
rect 19936 19572 19992 19628
rect 20040 19572 20096 19628
rect 6532 18788 6588 18844
rect 6636 18788 6692 18844
rect 6740 18788 6796 18844
rect 11852 18788 11908 18844
rect 11956 18788 12012 18844
rect 12060 18788 12116 18844
rect 17172 18788 17228 18844
rect 17276 18788 17332 18844
rect 17380 18788 17436 18844
rect 22492 18788 22548 18844
rect 22596 18788 22652 18844
rect 22700 18788 22756 18844
rect 3872 18004 3928 18060
rect 3976 18004 4032 18060
rect 4080 18004 4136 18060
rect 9192 18004 9248 18060
rect 9296 18004 9352 18060
rect 9400 18004 9456 18060
rect 14512 18004 14568 18060
rect 14616 18004 14672 18060
rect 14720 18004 14776 18060
rect 19832 18004 19888 18060
rect 19936 18004 19992 18060
rect 20040 18004 20096 18060
rect 6532 17220 6588 17276
rect 6636 17220 6692 17276
rect 6740 17220 6796 17276
rect 11852 17220 11908 17276
rect 11956 17220 12012 17276
rect 12060 17220 12116 17276
rect 17172 17220 17228 17276
rect 17276 17220 17332 17276
rect 17380 17220 17436 17276
rect 22492 17220 22548 17276
rect 22596 17220 22652 17276
rect 22700 17220 22756 17276
rect 3872 16436 3928 16492
rect 3976 16436 4032 16492
rect 4080 16436 4136 16492
rect 9192 16436 9248 16492
rect 9296 16436 9352 16492
rect 9400 16436 9456 16492
rect 14512 16436 14568 16492
rect 14616 16436 14672 16492
rect 14720 16436 14776 16492
rect 19832 16436 19888 16492
rect 19936 16436 19992 16492
rect 20040 16436 20096 16492
rect 6532 15652 6588 15708
rect 6636 15652 6692 15708
rect 6740 15652 6796 15708
rect 11852 15652 11908 15708
rect 11956 15652 12012 15708
rect 12060 15652 12116 15708
rect 17172 15652 17228 15708
rect 17276 15652 17332 15708
rect 17380 15652 17436 15708
rect 22492 15652 22548 15708
rect 22596 15652 22652 15708
rect 22700 15652 22756 15708
rect 3872 14868 3928 14924
rect 3976 14868 4032 14924
rect 4080 14868 4136 14924
rect 9192 14868 9248 14924
rect 9296 14868 9352 14924
rect 9400 14868 9456 14924
rect 14512 14868 14568 14924
rect 14616 14868 14672 14924
rect 14720 14868 14776 14924
rect 19832 14868 19888 14924
rect 19936 14868 19992 14924
rect 20040 14868 20096 14924
rect 6532 14084 6588 14140
rect 6636 14084 6692 14140
rect 6740 14084 6796 14140
rect 11852 14084 11908 14140
rect 11956 14084 12012 14140
rect 12060 14084 12116 14140
rect 17172 14084 17228 14140
rect 17276 14084 17332 14140
rect 17380 14084 17436 14140
rect 22492 14084 22548 14140
rect 22596 14084 22652 14140
rect 22700 14084 22756 14140
rect 4284 13692 4340 13748
rect 3872 13300 3928 13356
rect 3976 13300 4032 13356
rect 4080 13300 4136 13356
rect 9192 13300 9248 13356
rect 9296 13300 9352 13356
rect 9400 13300 9456 13356
rect 14512 13300 14568 13356
rect 14616 13300 14672 13356
rect 14720 13300 14776 13356
rect 19832 13300 19888 13356
rect 19936 13300 19992 13356
rect 20040 13300 20096 13356
rect 6532 12516 6588 12572
rect 6636 12516 6692 12572
rect 6740 12516 6796 12572
rect 11852 12516 11908 12572
rect 11956 12516 12012 12572
rect 12060 12516 12116 12572
rect 17172 12516 17228 12572
rect 17276 12516 17332 12572
rect 17380 12516 17436 12572
rect 22492 12516 22548 12572
rect 22596 12516 22652 12572
rect 22700 12516 22756 12572
rect 4284 12236 4340 12292
rect 3872 11732 3928 11788
rect 3976 11732 4032 11788
rect 4080 11732 4136 11788
rect 9192 11732 9248 11788
rect 9296 11732 9352 11788
rect 9400 11732 9456 11788
rect 14512 11732 14568 11788
rect 14616 11732 14672 11788
rect 14720 11732 14776 11788
rect 19832 11732 19888 11788
rect 19936 11732 19992 11788
rect 20040 11732 20096 11788
rect 3164 11340 3220 11396
rect 6532 10948 6588 11004
rect 6636 10948 6692 11004
rect 6740 10948 6796 11004
rect 11852 10948 11908 11004
rect 11956 10948 12012 11004
rect 12060 10948 12116 11004
rect 17172 10948 17228 11004
rect 17276 10948 17332 11004
rect 17380 10948 17436 11004
rect 22492 10948 22548 11004
rect 22596 10948 22652 11004
rect 22700 10948 22756 11004
rect 3872 10164 3928 10220
rect 3976 10164 4032 10220
rect 4080 10164 4136 10220
rect 9192 10164 9248 10220
rect 9296 10164 9352 10220
rect 9400 10164 9456 10220
rect 14512 10164 14568 10220
rect 14616 10164 14672 10220
rect 14720 10164 14776 10220
rect 19832 10164 19888 10220
rect 19936 10164 19992 10220
rect 20040 10164 20096 10220
rect 3164 9660 3220 9716
rect 6532 9380 6588 9436
rect 6636 9380 6692 9436
rect 6740 9380 6796 9436
rect 11852 9380 11908 9436
rect 11956 9380 12012 9436
rect 12060 9380 12116 9436
rect 17172 9380 17228 9436
rect 17276 9380 17332 9436
rect 17380 9380 17436 9436
rect 22492 9380 22548 9436
rect 22596 9380 22652 9436
rect 22700 9380 22756 9436
rect 3872 8596 3928 8652
rect 3976 8596 4032 8652
rect 4080 8596 4136 8652
rect 9192 8596 9248 8652
rect 9296 8596 9352 8652
rect 9400 8596 9456 8652
rect 14512 8596 14568 8652
rect 14616 8596 14672 8652
rect 14720 8596 14776 8652
rect 19832 8596 19888 8652
rect 19936 8596 19992 8652
rect 20040 8596 20096 8652
rect 6532 7812 6588 7868
rect 6636 7812 6692 7868
rect 6740 7812 6796 7868
rect 11852 7812 11908 7868
rect 11956 7812 12012 7868
rect 12060 7812 12116 7868
rect 17172 7812 17228 7868
rect 17276 7812 17332 7868
rect 17380 7812 17436 7868
rect 22492 7812 22548 7868
rect 22596 7812 22652 7868
rect 22700 7812 22756 7868
rect 3872 7028 3928 7084
rect 3976 7028 4032 7084
rect 4080 7028 4136 7084
rect 9192 7028 9248 7084
rect 9296 7028 9352 7084
rect 9400 7028 9456 7084
rect 14512 7028 14568 7084
rect 14616 7028 14672 7084
rect 14720 7028 14776 7084
rect 19832 7028 19888 7084
rect 19936 7028 19992 7084
rect 20040 7028 20096 7084
rect 6532 6244 6588 6300
rect 6636 6244 6692 6300
rect 6740 6244 6796 6300
rect 11852 6244 11908 6300
rect 11956 6244 12012 6300
rect 12060 6244 12116 6300
rect 17172 6244 17228 6300
rect 17276 6244 17332 6300
rect 17380 6244 17436 6300
rect 22492 6244 22548 6300
rect 22596 6244 22652 6300
rect 22700 6244 22756 6300
rect 3872 5460 3928 5516
rect 3976 5460 4032 5516
rect 4080 5460 4136 5516
rect 9192 5460 9248 5516
rect 9296 5460 9352 5516
rect 9400 5460 9456 5516
rect 14512 5460 14568 5516
rect 14616 5460 14672 5516
rect 14720 5460 14776 5516
rect 19832 5460 19888 5516
rect 19936 5460 19992 5516
rect 20040 5460 20096 5516
rect 6532 4676 6588 4732
rect 6636 4676 6692 4732
rect 6740 4676 6796 4732
rect 11852 4676 11908 4732
rect 11956 4676 12012 4732
rect 12060 4676 12116 4732
rect 17172 4676 17228 4732
rect 17276 4676 17332 4732
rect 17380 4676 17436 4732
rect 22492 4676 22548 4732
rect 22596 4676 22652 4732
rect 22700 4676 22756 4732
rect 3872 3892 3928 3948
rect 3976 3892 4032 3948
rect 4080 3892 4136 3948
rect 9192 3892 9248 3948
rect 9296 3892 9352 3948
rect 9400 3892 9456 3948
rect 14512 3892 14568 3948
rect 14616 3892 14672 3948
rect 14720 3892 14776 3948
rect 19832 3892 19888 3948
rect 19936 3892 19992 3948
rect 20040 3892 20096 3948
rect 6532 3108 6588 3164
rect 6636 3108 6692 3164
rect 6740 3108 6796 3164
rect 11852 3108 11908 3164
rect 11956 3108 12012 3164
rect 12060 3108 12116 3164
rect 17172 3108 17228 3164
rect 17276 3108 17332 3164
rect 17380 3108 17436 3164
rect 22492 3108 22548 3164
rect 22596 3108 22652 3164
rect 22700 3108 22756 3164
<< metal4 >>
rect 3844 19628 4164 20444
rect 3844 19572 3872 19628
rect 3928 19572 3976 19628
rect 4032 19572 4080 19628
rect 4136 19572 4164 19628
rect 3844 18060 4164 19572
rect 3844 18004 3872 18060
rect 3928 18004 3976 18060
rect 4032 18004 4080 18060
rect 4136 18004 4164 18060
rect 3844 16492 4164 18004
rect 3844 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4164 16492
rect 3844 14924 4164 16436
rect 3844 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4164 14924
rect 3844 13356 4164 14868
rect 6504 20412 6824 20444
rect 6504 20356 6532 20412
rect 6588 20356 6636 20412
rect 6692 20356 6740 20412
rect 6796 20356 6824 20412
rect 6504 18844 6824 20356
rect 6504 18788 6532 18844
rect 6588 18788 6636 18844
rect 6692 18788 6740 18844
rect 6796 18788 6824 18844
rect 6504 17276 6824 18788
rect 6504 17220 6532 17276
rect 6588 17220 6636 17276
rect 6692 17220 6740 17276
rect 6796 17220 6824 17276
rect 6504 15708 6824 17220
rect 6504 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6824 15708
rect 6504 14140 6824 15652
rect 6504 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6824 14140
rect 3844 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4164 13356
rect 3844 11788 4164 13300
rect 4284 13748 4340 13758
rect 4284 12292 4340 13692
rect 4284 12226 4340 12236
rect 6504 12572 6824 14084
rect 6504 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6824 12572
rect 3844 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4164 11788
rect 3164 11396 3220 11406
rect 3164 9716 3220 11340
rect 3164 9650 3220 9660
rect 3844 10220 4164 11732
rect 3844 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4164 10220
rect 3844 8652 4164 10164
rect 3844 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4164 8652
rect 3844 7084 4164 8596
rect 3844 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4164 7084
rect 3844 5516 4164 7028
rect 3844 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4164 5516
rect 3844 3948 4164 5460
rect 3844 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4164 3948
rect 3844 3076 4164 3892
rect 6504 11004 6824 12516
rect 6504 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6824 11004
rect 6504 9436 6824 10948
rect 6504 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6824 9436
rect 6504 7868 6824 9380
rect 6504 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6824 7868
rect 6504 6300 6824 7812
rect 6504 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6824 6300
rect 6504 4732 6824 6244
rect 6504 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6824 4732
rect 6504 3164 6824 4676
rect 6504 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6824 3164
rect 6504 3076 6824 3108
rect 9164 19628 9484 20444
rect 9164 19572 9192 19628
rect 9248 19572 9296 19628
rect 9352 19572 9400 19628
rect 9456 19572 9484 19628
rect 9164 18060 9484 19572
rect 9164 18004 9192 18060
rect 9248 18004 9296 18060
rect 9352 18004 9400 18060
rect 9456 18004 9484 18060
rect 9164 16492 9484 18004
rect 9164 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9484 16492
rect 9164 14924 9484 16436
rect 9164 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9484 14924
rect 9164 13356 9484 14868
rect 9164 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9484 13356
rect 9164 11788 9484 13300
rect 9164 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9484 11788
rect 9164 10220 9484 11732
rect 9164 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9484 10220
rect 9164 8652 9484 10164
rect 9164 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9484 8652
rect 9164 7084 9484 8596
rect 9164 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9484 7084
rect 9164 5516 9484 7028
rect 9164 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9484 5516
rect 9164 3948 9484 5460
rect 9164 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9484 3948
rect 9164 3076 9484 3892
rect 11824 20412 12144 20444
rect 11824 20356 11852 20412
rect 11908 20356 11956 20412
rect 12012 20356 12060 20412
rect 12116 20356 12144 20412
rect 11824 18844 12144 20356
rect 11824 18788 11852 18844
rect 11908 18788 11956 18844
rect 12012 18788 12060 18844
rect 12116 18788 12144 18844
rect 11824 17276 12144 18788
rect 11824 17220 11852 17276
rect 11908 17220 11956 17276
rect 12012 17220 12060 17276
rect 12116 17220 12144 17276
rect 11824 15708 12144 17220
rect 11824 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12144 15708
rect 11824 14140 12144 15652
rect 11824 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12144 14140
rect 11824 12572 12144 14084
rect 11824 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12144 12572
rect 11824 11004 12144 12516
rect 11824 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12144 11004
rect 11824 9436 12144 10948
rect 11824 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12144 9436
rect 11824 7868 12144 9380
rect 11824 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12144 7868
rect 11824 6300 12144 7812
rect 11824 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12144 6300
rect 11824 4732 12144 6244
rect 11824 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12144 4732
rect 11824 3164 12144 4676
rect 11824 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12144 3164
rect 11824 3076 12144 3108
rect 14484 19628 14804 20444
rect 14484 19572 14512 19628
rect 14568 19572 14616 19628
rect 14672 19572 14720 19628
rect 14776 19572 14804 19628
rect 14484 18060 14804 19572
rect 14484 18004 14512 18060
rect 14568 18004 14616 18060
rect 14672 18004 14720 18060
rect 14776 18004 14804 18060
rect 14484 16492 14804 18004
rect 14484 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14804 16492
rect 14484 14924 14804 16436
rect 14484 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14804 14924
rect 14484 13356 14804 14868
rect 14484 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14804 13356
rect 14484 11788 14804 13300
rect 14484 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14804 11788
rect 14484 10220 14804 11732
rect 14484 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14804 10220
rect 14484 8652 14804 10164
rect 14484 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14804 8652
rect 14484 7084 14804 8596
rect 14484 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14804 7084
rect 14484 5516 14804 7028
rect 14484 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14804 5516
rect 14484 3948 14804 5460
rect 14484 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14804 3948
rect 14484 3076 14804 3892
rect 17144 20412 17464 20444
rect 17144 20356 17172 20412
rect 17228 20356 17276 20412
rect 17332 20356 17380 20412
rect 17436 20356 17464 20412
rect 17144 18844 17464 20356
rect 17144 18788 17172 18844
rect 17228 18788 17276 18844
rect 17332 18788 17380 18844
rect 17436 18788 17464 18844
rect 17144 17276 17464 18788
rect 17144 17220 17172 17276
rect 17228 17220 17276 17276
rect 17332 17220 17380 17276
rect 17436 17220 17464 17276
rect 17144 15708 17464 17220
rect 17144 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17464 15708
rect 17144 14140 17464 15652
rect 17144 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17464 14140
rect 17144 12572 17464 14084
rect 17144 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17464 12572
rect 17144 11004 17464 12516
rect 17144 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17464 11004
rect 17144 9436 17464 10948
rect 17144 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17464 9436
rect 17144 7868 17464 9380
rect 17144 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17464 7868
rect 17144 6300 17464 7812
rect 17144 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17464 6300
rect 17144 4732 17464 6244
rect 17144 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17464 4732
rect 17144 3164 17464 4676
rect 17144 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17464 3164
rect 17144 3076 17464 3108
rect 19804 19628 20124 20444
rect 19804 19572 19832 19628
rect 19888 19572 19936 19628
rect 19992 19572 20040 19628
rect 20096 19572 20124 19628
rect 19804 18060 20124 19572
rect 19804 18004 19832 18060
rect 19888 18004 19936 18060
rect 19992 18004 20040 18060
rect 20096 18004 20124 18060
rect 19804 16492 20124 18004
rect 19804 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20124 16492
rect 19804 14924 20124 16436
rect 19804 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20124 14924
rect 19804 13356 20124 14868
rect 19804 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20124 13356
rect 19804 11788 20124 13300
rect 19804 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20124 11788
rect 19804 10220 20124 11732
rect 19804 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20124 10220
rect 19804 8652 20124 10164
rect 19804 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20124 8652
rect 19804 7084 20124 8596
rect 19804 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20124 7084
rect 19804 5516 20124 7028
rect 19804 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20124 5516
rect 19804 3948 20124 5460
rect 19804 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20124 3948
rect 19804 3076 20124 3892
rect 22464 20412 22784 20444
rect 22464 20356 22492 20412
rect 22548 20356 22596 20412
rect 22652 20356 22700 20412
rect 22756 20356 22784 20412
rect 22464 18844 22784 20356
rect 22464 18788 22492 18844
rect 22548 18788 22596 18844
rect 22652 18788 22700 18844
rect 22756 18788 22784 18844
rect 22464 17276 22784 18788
rect 22464 17220 22492 17276
rect 22548 17220 22596 17276
rect 22652 17220 22700 17276
rect 22756 17220 22784 17276
rect 22464 15708 22784 17220
rect 22464 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22784 15708
rect 22464 14140 22784 15652
rect 22464 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22784 14140
rect 22464 12572 22784 14084
rect 22464 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22784 12572
rect 22464 11004 22784 12516
rect 22464 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22784 11004
rect 22464 9436 22784 10948
rect 22464 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22784 9436
rect 22464 7868 22784 9380
rect 22464 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22784 7868
rect 22464 6300 22784 7812
rect 22464 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22784 6300
rect 22464 4732 22784 6244
rect 22464 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22784 4732
rect 22464 3164 22784 4676
rect 22464 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22784 3164
rect 22464 3076 22784 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _100_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10528 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698431365
transform -1 0 16128 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _103_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _104_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13776 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698431365
transform -1 0 19600 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _106_
timestamp 1698431365
transform -1 0 18704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698431365
transform -1 0 18256 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698431365
transform -1 0 18592 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _109_
timestamp 1698431365
transform -1 0 20160 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698431365
transform 1 0 9520 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _111_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15680 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _113_
timestamp 1698431365
transform -1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698431365
transform -1 0 16240 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _115_
timestamp 1698431365
transform -1 0 20384 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698431365
transform -1 0 14784 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698431365
transform 1 0 14784 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _118_
timestamp 1698431365
transform -1 0 15792 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _119_
timestamp 1698431365
transform -1 0 16688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698431365
transform -1 0 14784 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698431365
transform -1 0 16688 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _122_
timestamp 1698431365
transform -1 0 17808 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698431365
transform -1 0 16016 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _124_
timestamp 1698431365
transform -1 0 12880 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _125_
timestamp 1698431365
transform -1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _126_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11200 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698431365
transform -1 0 11312 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698431365
transform -1 0 10080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _130_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _131_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _132_
timestamp 1698431365
transform -1 0 20832 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698431365
transform 1 0 17920 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _134_
timestamp 1698431365
transform -1 0 19824 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698431365
transform 1 0 13888 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _136_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15456 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698431365
transform -1 0 5152 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _138_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1698431365
transform -1 0 21840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _140_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _141_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _142_
timestamp 1698431365
transform -1 0 20160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _143_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698431365
transform 1 0 4592 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1698431365
transform 1 0 4368 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1698431365
transform -1 0 6160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698431365
transform 1 0 4368 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _149_
timestamp 1698431365
transform -1 0 5712 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698431365
transform -1 0 14336 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _151_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698431365
transform 1 0 16128 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _154_
timestamp 1698431365
transform -1 0 9856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _155_
timestamp 1698431365
transform -1 0 10752 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _156_
timestamp 1698431365
transform -1 0 9184 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _157_
timestamp 1698431365
transform 1 0 6384 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _158_
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _159_
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _160_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1698431365
transform -1 0 21616 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _162_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _163_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7280 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _164_
timestamp 1698431365
transform -1 0 6384 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _165_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4704 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _166_
timestamp 1698431365
transform 1 0 2576 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _167_
timestamp 1698431365
transform -1 0 11536 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _168_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698431365
transform -1 0 3920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _170_
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_
timestamp 1698431365
transform -1 0 4704 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _172_
timestamp 1698431365
transform -1 0 9968 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _173_
timestamp 1698431365
transform 1 0 10192 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _174_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _175_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _176_
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _177_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _178_
timestamp 1698431365
transform 1 0 10640 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _179_
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _180_
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _181_
timestamp 1698431365
transform -1 0 15344 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _182_
timestamp 1698431365
transform -1 0 10640 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698431365
transform 1 0 4592 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _184_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _185_
timestamp 1698431365
transform -1 0 11984 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _186_
timestamp 1698431365
transform 1 0 9968 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _187_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _188_
timestamp 1698431365
transform 1 0 4144 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _189_
timestamp 1698431365
transform 1 0 4368 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _190_
timestamp 1698431365
transform -1 0 21840 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _191_
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _192_
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _193_
timestamp 1698431365
transform 1 0 20160 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _194_
timestamp 1698431365
transform -1 0 19936 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _195_
timestamp 1698431365
transform 1 0 19936 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _196_
timestamp 1698431365
transform -1 0 20608 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _197_
timestamp 1698431365
transform 1 0 20832 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _198_
timestamp 1698431365
transform -1 0 21616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _199_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17808 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10192 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _201_
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _202_
timestamp 1698431365
transform 1 0 19936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _203_
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _204_
timestamp 1698431365
transform 1 0 18816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _205_
timestamp 1698431365
transform -1 0 18144 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _206_
timestamp 1698431365
transform -1 0 7056 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _207_
timestamp 1698431365
transform -1 0 6384 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _208_
timestamp 1698431365
transform 1 0 5712 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _209_
timestamp 1698431365
transform -1 0 16576 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _210_
timestamp 1698431365
transform 1 0 15008 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _211_
timestamp 1698431365
transform -1 0 15232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _212_
timestamp 1698431365
transform -1 0 13440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _213_
timestamp 1698431365
transform 1 0 10864 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _214_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _215_
timestamp 1698431365
transform 1 0 12320 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _216_
timestamp 1698431365
transform 1 0 11088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _217_
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _218_
timestamp 1698431365
transform 1 0 11312 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _219_
timestamp 1698431365
transform 1 0 20160 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _220_
timestamp 1698431365
transform 1 0 2688 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _221_
timestamp 1698431365
transform 1 0 2800 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _222_
timestamp 1698431365
transform 1 0 2912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _223_
timestamp 1698431365
transform -1 0 4816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _224_
timestamp 1698431365
transform 1 0 3696 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _225_
timestamp 1698431365
transform -1 0 3696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _226_
timestamp 1698431365
transform 1 0 3472 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _227_
timestamp 1698431365
transform 1 0 3920 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _228_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2800 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _229_
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _230_
timestamp 1698431365
transform 1 0 19040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _231_
timestamp 1698431365
transform 1 0 17808 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _232_
timestamp 1698431365
transform 1 0 19040 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _233_
timestamp 1698431365
transform -1 0 16128 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _234_
timestamp 1698431365
transform -1 0 15456 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _235_
timestamp 1698431365
transform -1 0 15680 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _236_
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _238_
timestamp 1698431365
transform -1 0 19040 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _239_
timestamp 1698431365
transform 1 0 18256 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__I
timestamp 1698431365
transform 1 0 18480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1698431365
transform -1 0 8736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__A1
timestamp 1698431365
transform 1 0 9408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__A1
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__B
timestamp 1698431365
transform 1 0 10304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__A1
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__A1
timestamp 1698431365
transform 1 0 19488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__B
timestamp 1698431365
transform 1 0 12208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__A1
timestamp 1698431365
transform -1 0 4032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A1
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 22176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 21728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 21728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 22400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 21728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 21728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_174 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_182
timestamp 1698431365
transform 1 0 21728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_186 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_179
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_82
timestamp 1698431365
transform 1 0 10528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_84
timestamp 1698431365
transform 1 0 10752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_91
timestamp 1698431365
transform 1 0 11536 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_123
timestamp 1698431365
transform 1 0 15120 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_144
timestamp 1698431365
transform 1 0 17472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_151
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_155
timestamp 1698431365
transform 1 0 18704 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_187
timestamp 1698431365
transform 1 0 22288 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_18
timestamp 1698431365
transform 1 0 3360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_26
timestamp 1698431365
transform 1 0 4256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_28
timestamp 1698431365
transform 1 0 4480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_43
timestamp 1698431365
transform 1 0 6160 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_59
timestamp 1698431365
transform 1 0 7952 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_67
timestamp 1698431365
transform 1 0 8848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_88
timestamp 1698431365
transform 1 0 11200 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_95
timestamp 1698431365
transform 1 0 11984 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_133
timestamp 1698431365
transform 1 0 16240 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_141
timestamp 1698431365
transform 1 0 17136 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_145
timestamp 1698431365
transform 1 0 17584 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_150
timestamp 1698431365
transform 1 0 18144 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_166
timestamp 1698431365
transform 1 0 19936 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_183
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_187
timestamp 1698431365
transform 1 0 22288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_18
timestamp 1698431365
transform 1 0 3360 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_26
timestamp 1698431365
transform 1 0 4256 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_36
timestamp 1698431365
transform 1 0 5376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_40
timestamp 1698431365
transform 1 0 5824 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_56
timestamp 1698431365
transform 1 0 7616 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_64
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_89
timestamp 1698431365
transform 1 0 11312 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_105
timestamp 1698431365
transform 1 0 13104 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_113
timestamp 1698431365
transform 1 0 14000 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_117
timestamp 1698431365
transform 1 0 14448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_119
timestamp 1698431365
transform 1 0 14672 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_126
timestamp 1698431365
transform 1 0 15456 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_134
timestamp 1698431365
transform 1 0 16352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_146
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_154
timestamp 1698431365
transform 1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_170
timestamp 1698431365
transform 1 0 20384 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_18
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_22
timestamp 1698431365
transform 1 0 3808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_24
timestamp 1698431365
transform 1 0 4032 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_47
timestamp 1698431365
transform 1 0 6608 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_63
timestamp 1698431365
transform 1 0 8400 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_71
timestamp 1698431365
transform 1 0 9296 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_94
timestamp 1698431365
transform 1 0 11872 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_102
timestamp 1698431365
transform 1 0 12768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_111
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_113
timestamp 1698431365
transform 1 0 14000 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_120
timestamp 1698431365
transform 1 0 14784 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_137
timestamp 1698431365
transform 1 0 16688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_153
timestamp 1698431365
transform 1 0 18480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_173
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_35
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_48
timestamp 1698431365
transform 1 0 6720 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_64
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_74
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_87
timestamp 1698431365
transform 1 0 11088 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_119
timestamp 1698431365
transform 1 0 14672 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_135
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_168
timestamp 1698431365
transform 1 0 20160 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_184
timestamp 1698431365
transform 1 0 21952 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_10
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_30
timestamp 1698431365
transform 1 0 4704 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_43
timestamp 1698431365
transform 1 0 6160 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_59
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_67
timestamp 1698431365
transform 1 0 8848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_81
timestamp 1698431365
transform 1 0 10416 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_97
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_139
timestamp 1698431365
transform 1 0 16912 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_155
timestamp 1698431365
transform 1 0 18704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_187
timestamp 1698431365
transform 1 0 22288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_10
timestamp 1698431365
transform 1 0 2464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_21
timestamp 1698431365
transform 1 0 3696 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_53
timestamp 1698431365
transform 1 0 7280 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_76
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_108
timestamp 1698431365
transform 1 0 13440 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_112
timestamp 1698431365
transform 1 0 13888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_162
timestamp 1698431365
transform 1 0 19488 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_168
timestamp 1698431365
transform 1 0 20160 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_176
timestamp 1698431365
transform 1 0 21056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_23
timestamp 1698431365
transform 1 0 3920 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_73
timestamp 1698431365
transform 1 0 9520 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_75
timestamp 1698431365
transform 1 0 9744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_84
timestamp 1698431365
transform 1 0 10752 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_92
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_94
timestamp 1698431365
transform 1 0 11872 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_137
timestamp 1698431365
transform 1 0 16688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_147
timestamp 1698431365
transform 1 0 17808 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_154
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_162
timestamp 1698431365
transform 1 0 19488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_166
timestamp 1698431365
transform 1 0 19936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_26
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_50
timestamp 1698431365
transform 1 0 6944 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_58
timestamp 1698431365
transform 1 0 7840 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_95
timestamp 1698431365
transform 1 0 11984 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_127
timestamp 1698431365
transform 1 0 15568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_135
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_155
timestamp 1698431365
transform 1 0 18704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_165
timestamp 1698431365
transform 1 0 19824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_167
timestamp 1698431365
transform 1 0 20048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_186
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_43
timestamp 1698431365
transform 1 0 6160 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_59
timestamp 1698431365
transform 1 0 7952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_70
timestamp 1698431365
transform 1 0 9184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_74
timestamp 1698431365
transform 1 0 9632 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_76
timestamp 1698431365
transform 1 0 9856 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_115
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_136
timestamp 1698431365
transform 1 0 16576 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_144
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_146
timestamp 1698431365
transform 1 0 17696 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_163
timestamp 1698431365
transform 1 0 19600 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_10
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_43
timestamp 1698431365
transform 1 0 6160 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_59
timestamp 1698431365
transform 1 0 7952 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_79
timestamp 1698431365
transform 1 0 10192 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_111
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_127
timestamp 1698431365
transform 1 0 15568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_135
timestamp 1698431365
transform 1 0 16464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_174
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_178
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_33
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_63
timestamp 1698431365
transform 1 0 8400 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_73
timestamp 1698431365
transform 1 0 9520 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_77
timestamp 1698431365
transform 1 0 9968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_79
timestamp 1698431365
transform 1 0 10192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_82
timestamp 1698431365
transform 1 0 10528 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_98
timestamp 1698431365
transform 1 0 12320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_102
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_124
timestamp 1698431365
transform 1 0 15232 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_156
timestamp 1698431365
transform 1 0 18816 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_10
timestamp 1698431365
transform 1 0 2464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_14
timestamp 1698431365
transform 1 0 2912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_16
timestamp 1698431365
transform 1 0 3136 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_21
timestamp 1698431365
transform 1 0 3696 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_53
timestamp 1698431365
transform 1 0 7280 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_61
timestamp 1698431365
transform 1 0 8176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_63
timestamp 1698431365
transform 1 0 8400 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_88
timestamp 1698431365
transform 1 0 11200 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698431365
transform 1 0 13440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_132
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_152
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_156
timestamp 1698431365
transform 1 0 18816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_182
timestamp 1698431365
transform 1 0 21728 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_186
timestamp 1698431365
transform 1 0 22176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_18
timestamp 1698431365
transform 1 0 3360 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_26
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_33
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_77
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_119
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_128
timestamp 1698431365
transform 1 0 15680 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_144
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_152
timestamp 1698431365
transform 1 0 18368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_156
timestamp 1698431365
transform 1 0 18816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_181
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_25
timestamp 1698431365
transform 1 0 4144 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_57
timestamp 1698431365
transform 1 0 7728 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_65
timestamp 1698431365
transform 1 0 8624 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_82
timestamp 1698431365
transform 1 0 10528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_84
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_95
timestamp 1698431365
transform 1 0 11984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_99
timestamp 1698431365
transform 1 0 12432 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_115
timestamp 1698431365
transform 1 0 14224 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_119
timestamp 1698431365
transform 1 0 14672 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_132
timestamp 1698431365
transform 1 0 16128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698431365
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_10
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_12
timestamp 1698431365
transform 1 0 2688 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_69
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_77
timestamp 1698431365
transform 1 0 9968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_79
timestamp 1698431365
transform 1 0 10192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_155
timestamp 1698431365
transform 1 0 18704 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_159
timestamp 1698431365
transform 1 0 19152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_161
timestamp 1698431365
transform 1 0 19376 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_12
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_29
timestamp 1698431365
transform 1 0 4592 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_37
timestamp 1698431365
transform 1 0 5488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_61
timestamp 1698431365
transform 1 0 8176 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_65
timestamp 1698431365
transform 1 0 8624 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_95
timestamp 1698431365
transform 1 0 11984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_97
timestamp 1698431365
transform 1 0 12208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_108
timestamp 1698431365
transform 1 0 13440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_110
timestamp 1698431365
transform 1 0 13664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_119
timestamp 1698431365
transform 1 0 14672 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_123
timestamp 1698431365
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_125
timestamp 1698431365
transform 1 0 15344 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_156
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_172
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_10
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_20
timestamp 1698431365
transform 1 0 3584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_24
timestamp 1698431365
transform 1 0 4032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_57
timestamp 1698431365
transform 1 0 7728 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_73
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_80
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_88
timestamp 1698431365
transform 1 0 11200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_95
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_113
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_121
timestamp 1698431365
transform 1 0 14896 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_128
timestamp 1698431365
transform 1 0 15680 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_144
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_146
timestamp 1698431365
transform 1 0 17696 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_157
timestamp 1698431365
transform 1 0 18928 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_166
timestamp 1698431365
transform 1 0 19936 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_187
timestamp 1698431365
transform 1 0 22288 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_4
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_11
timestamp 1698431365
transform 1 0 2576 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_19
timestamp 1698431365
transform 1 0 3472 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_23
timestamp 1698431365
transform 1 0 3920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_31
timestamp 1698431365
transform 1 0 4816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_33
timestamp 1698431365
transform 1 0 5040 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_36
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_44
timestamp 1698431365
transform 1 0 6272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_51
timestamp 1698431365
transform 1 0 7056 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_76
timestamp 1698431365
transform 1 0 9856 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_84
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_91
timestamp 1698431365
transform 1 0 11536 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_99
timestamp 1698431365
transform 1 0 12432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_101
timestamp 1698431365
transform 1 0 12656 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_104
timestamp 1698431365
transform 1 0 12992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_111
timestamp 1698431365
transform 1 0 13776 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_119
timestamp 1698431365
transform 1 0 14672 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_123
timestamp 1698431365
transform 1 0 15120 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_131
timestamp 1698431365
transform 1 0 16016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_135
timestamp 1698431365
transform 1 0 16464 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_138
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698431365
transform 1 0 17472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_151
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_153
timestamp 1698431365
transform 1 0 18480 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_158
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_162
timestamp 1698431365
transform 1 0 19488 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_178
timestamp 1698431365
transform 1 0 21280 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 22400 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 22400 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 22400 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 22400 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 22400 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform -1 0 22400 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output7
timestamp 1698431365
transform 1 0 19712 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output8
timestamp 1698431365
transform -1 0 2576 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output9
timestamp 1698431365
transform -1 0 4816 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output10
timestamp 1698431365
transform -1 0 7056 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output11
timestamp 1698431365
transform -1 0 9856 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output12
timestamp 1698431365
transform -1 0 11536 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output13
timestamp 1698431365
transform -1 0 13776 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output14
timestamp 1698431365
transform -1 0 16016 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output15
timestamp 1698431365
transform -1 0 18256 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output16
timestamp 1698431365
transform -1 0 21280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output17
timestamp 1698431365
transform 1 0 21728 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_22 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 22624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_23
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 22624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_24
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 22624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_25
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 22624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_26
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 22624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_27
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 22624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_28
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 22624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_29
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_30
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 22624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_31
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_32
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 22624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_33
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_34
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 22624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_35
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 22624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_36
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 22624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_37
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_38
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_39
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 22624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_40
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 22624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_41
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 22624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_42
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_43
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 22624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_46
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_47
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_48
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_51
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_52
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_54
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_55
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_56
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_57
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_58
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_59
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_60
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_61
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_62
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_63
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_64
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_65
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_66
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_67
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_68
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_69
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_70
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_71
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_72
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_73
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_74
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_75
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_76
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_77
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_78
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_79
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_80
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_81
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_82
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_83
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_84
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_85
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_86
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_87
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_88
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_89
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_90
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_91
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_92
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_93
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_94
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_95
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_96
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_97
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_98
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_99
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_100
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_101
timestamp 1698431365
transform 1 0 12768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_102
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_103
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -86 -86 310 870
<< labels >>
flabel metal3 s 23200 1568 24000 1680 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 23200 7392 24000 7504 0 FreeSans 448 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 23200 10304 24000 10416 0 FreeSans 448 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 23200 13216 24000 13328 0 FreeSans 448 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 23200 16128 24000 16240 0 FreeSans 448 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 23200 19040 24000 19152 0 FreeSans 448 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal3 s 23200 21952 24000 22064 0 FreeSans 448 0 0 0 io_oeb
port 6 nsew signal tristate
flabel metal2 s 1792 23200 1904 24000 0 FreeSans 448 90 0 0 io_out[0]
port 7 nsew signal tristate
flabel metal2 s 4032 23200 4144 24000 0 FreeSans 448 90 0 0 io_out[1]
port 8 nsew signal tristate
flabel metal2 s 6272 23200 6384 24000 0 FreeSans 448 90 0 0 io_out[2]
port 9 nsew signal tristate
flabel metal2 s 8512 23200 8624 24000 0 FreeSans 448 90 0 0 io_out[3]
port 10 nsew signal tristate
flabel metal2 s 10752 23200 10864 24000 0 FreeSans 448 90 0 0 io_out[4]
port 11 nsew signal tristate
flabel metal2 s 12992 23200 13104 24000 0 FreeSans 448 90 0 0 io_out[5]
port 12 nsew signal tristate
flabel metal2 s 15232 23200 15344 24000 0 FreeSans 448 90 0 0 io_out[6]
port 13 nsew signal tristate
flabel metal2 s 17472 23200 17584 24000 0 FreeSans 448 90 0 0 io_out[7]
port 14 nsew signal tristate
flabel metal2 s 19712 23200 19824 24000 0 FreeSans 448 90 0 0 io_out[8]
port 15 nsew signal tristate
flabel metal2 s 21952 23200 22064 24000 0 FreeSans 448 90 0 0 io_out[9]
port 16 nsew signal tristate
flabel metal3 s 23200 4480 24000 4592 0 FreeSans 448 0 0 0 rst_n
port 17 nsew signal input
flabel metal4 s 3844 3076 4164 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 9164 3076 9484 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 14484 3076 14804 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 19804 3076 20124 20444 0 FreeSans 1280 90 0 0 vdd
port 18 nsew power bidirectional
flabel metal4 s 6504 3076 6824 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 11824 3076 12144 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 17144 3076 17464 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
flabel metal4 s 22464 3076 22784 20444 0 FreeSans 1280 90 0 0 vss
port 19 nsew ground bidirectional
rlabel metal1 11984 19600 11984 19600 0 vdd
rlabel via1 12064 20384 12064 20384 0 vss
rlabel metal2 15288 12824 15288 12824 0 _000_
rlabel metal3 17360 11256 17360 11256 0 _001_
rlabel metal2 16184 11480 16184 11480 0 _002_
rlabel metal2 15512 11368 15512 11368 0 _003_
rlabel metal3 10528 15176 10528 15176 0 _004_
rlabel metal2 10864 15064 10864 15064 0 _005_
rlabel metal2 10528 15512 10528 15512 0 _006_
rlabel metal2 2968 16856 2968 16856 0 _007_
rlabel metal2 9856 15512 9856 15512 0 _008_
rlabel metal3 10136 17416 10136 17416 0 _009_
rlabel metal2 20328 11872 20328 11872 0 _010_
rlabel metal3 15960 12824 15960 12824 0 _011_
rlabel metal2 15624 12936 15624 12936 0 _012_
rlabel metal2 4984 12600 4984 12600 0 _013_
rlabel metal2 20216 10024 20216 10024 0 _014_
rlabel metal2 21448 18984 21448 18984 0 _015_
rlabel metal2 19544 10248 19544 10248 0 _016_
rlabel metal2 4872 6720 4872 6720 0 _017_
rlabel metal2 15064 16632 15064 16632 0 _018_
rlabel metal2 5768 13720 5768 13720 0 _019_
rlabel metal2 4984 9072 4984 9072 0 _020_
rlabel metal2 18256 15400 18256 15400 0 _021_
rlabel metal2 16632 18368 16632 18368 0 _022_
rlabel metal2 8512 12040 8512 12040 0 _023_
rlabel metal2 10024 10416 10024 10416 0 _024_
rlabel metal2 6664 17808 6664 17808 0 _025_
rlabel metal2 7112 18760 7112 18760 0 _026_
rlabel metal2 7560 18872 7560 18872 0 _027_
rlabel metal2 9240 14672 9240 14672 0 _028_
rlabel metal3 18312 7672 18312 7672 0 _029_
rlabel metal2 6888 18480 6888 18480 0 _030_
rlabel metal2 6216 16744 6216 16744 0 _031_
rlabel metal2 3528 13776 3528 13776 0 _032_
rlabel metal2 3416 10192 3416 10192 0 _033_
rlabel metal2 10416 7224 10416 7224 0 _034_
rlabel metal2 3080 9240 3080 9240 0 _035_
rlabel metal2 2968 10640 2968 10640 0 _036_
rlabel metal2 3192 10248 3192 10248 0 _037_
rlabel metal2 4760 8064 4760 8064 0 _038_
rlabel metal2 10248 7672 10248 7672 0 _039_
rlabel metal2 10472 12432 10472 12432 0 _040_
rlabel metal2 10808 10192 10808 10192 0 _041_
rlabel metal3 8400 8904 8400 8904 0 _042_
rlabel metal2 5656 7952 5656 7952 0 _043_
rlabel metal2 4312 8512 4312 8512 0 _044_
rlabel metal2 11144 8680 11144 8680 0 _045_
rlabel metal2 5824 9688 5824 9688 0 _046_
rlabel metal2 6328 9464 6328 9464 0 _047_
rlabel metal2 10472 8400 10472 8400 0 _048_
rlabel metal2 5992 8736 5992 8736 0 _049_
rlabel metal2 5544 8960 5544 8960 0 _050_
rlabel metal2 4872 8848 4872 8848 0 _051_
rlabel metal3 9968 11928 9968 11928 0 _052_
rlabel metal2 3584 14056 3584 14056 0 _053_
rlabel metal3 5432 8232 5432 8232 0 _054_
rlabel metal2 4648 7728 4648 7728 0 _055_
rlabel metal2 21728 16856 21728 16856 0 _056_
rlabel metal2 21560 12488 21560 12488 0 _057_
rlabel metal2 20216 16464 20216 16464 0 _058_
rlabel metal2 20328 17360 20328 17360 0 _059_
rlabel metal2 21280 16072 21280 16072 0 _060_
rlabel metal3 19208 15288 19208 15288 0 _061_
rlabel metal2 19208 14616 19208 14616 0 _062_
rlabel metal2 20664 15736 20664 15736 0 _063_
rlabel metal2 17976 7000 17976 7000 0 _064_
rlabel metal2 5880 18928 5880 18928 0 _065_
rlabel metal2 15288 18144 15288 18144 0 _066_
rlabel metal2 11480 16464 11480 16464 0 _067_
rlabel metal2 11816 16912 11816 16912 0 _068_
rlabel metal3 11368 17528 11368 17528 0 _069_
rlabel metal2 12040 18144 12040 18144 0 _070_
rlabel metal2 11760 18536 11760 18536 0 _071_
rlabel metal2 11032 18480 11032 18480 0 _072_
rlabel metal2 3192 16408 3192 16408 0 _073_
rlabel metal2 3528 18032 3528 18032 0 _074_
rlabel metal2 3192 18760 3192 18760 0 _075_
rlabel metal2 4536 18088 4536 18088 0 _076_
rlabel metal2 3304 16184 3304 16184 0 _077_
rlabel metal2 4536 13944 4536 13944 0 _078_
rlabel metal2 3808 16632 3808 16632 0 _079_
rlabel metal2 3080 17416 3080 17416 0 _080_
rlabel metal3 18648 19208 18648 19208 0 _081_
rlabel metal2 15960 16464 15960 16464 0 _082_
rlabel metal2 15456 16632 15456 16632 0 _083_
rlabel metal2 9408 15960 9408 15960 0 _084_
rlabel metal2 18760 19488 18760 19488 0 _085_
rlabel metal2 9800 7056 9800 7056 0 _086_
rlabel metal2 15960 18368 15960 18368 0 _087_
rlabel metal2 15624 18480 15624 18480 0 _088_
rlabel metal2 13944 18872 13944 18872 0 _089_
rlabel metal2 18312 12768 18312 12768 0 _090_
rlabel metal2 17752 6328 17752 6328 0 _091_
rlabel metal2 19320 12600 19320 12600 0 _092_
rlabel metal3 17808 9800 17808 9800 0 _093_
rlabel metal2 16184 12544 16184 12544 0 _094_
rlabel metal2 18032 15176 18032 15176 0 _095_
rlabel metal2 15512 8176 15512 8176 0 _096_
rlabel metal3 18200 8232 18200 8232 0 _097_
rlabel metal2 14280 7840 14280 7840 0 _098_
rlabel metal2 19768 15232 19768 15232 0 _099_
rlabel metal3 22666 1624 22666 1624 0 clk
rlabel metal3 22722 7448 22722 7448 0 io_in[0]
rlabel metal2 22232 10472 22232 10472 0 io_in[1]
rlabel metal2 22232 13496 22232 13496 0 io_in[2]
rlabel metal3 22778 16184 22778 16184 0 io_in[3]
rlabel metal2 22232 18760 22232 18760 0 io_in[4]
rlabel metal3 21658 22008 21658 22008 0 io_oeb
rlabel metal2 1848 21686 1848 21686 0 io_out[0]
rlabel metal2 4312 20888 4312 20888 0 io_out[1]
rlabel metal2 6552 20160 6552 20160 0 io_out[2]
rlabel metal2 9352 21672 9352 21672 0 io_out[3]
rlabel metal2 11032 20888 11032 20888 0 io_out[4]
rlabel metal2 13272 20888 13272 20888 0 io_out[5]
rlabel metal2 15288 21686 15288 21686 0 io_out[6]
rlabel metal2 17528 21686 17528 21686 0 io_out[7]
rlabel metal2 19768 21658 19768 21658 0 io_out[8]
rlabel metal2 22008 21686 22008 21686 0 io_out[9]
rlabel metal2 18648 18816 18648 18816 0 main.GATES_100.input2
rlabel metal2 15400 10416 15400 10416 0 main.GATES_102.input1
rlabel metal2 18032 11368 18032 11368 0 main.GATES_102.input2
rlabel metal2 13832 14784 13832 14784 0 main.GATES_102.input3
rlabel metal2 5992 18816 5992 18816 0 main.GATES_103.input2
rlabel metal2 6384 19320 6384 19320 0 main.GATES_105.input3
rlabel metal2 13048 18424 13048 18424 0 main.GATES_106.input2
rlabel metal2 19432 11760 19432 11760 0 main.GATES_107.input2
rlabel metal2 5824 13160 5824 13160 0 main.GATES_108.input1
rlabel metal2 11704 19264 11704 19264 0 main.GATES_109.input2
rlabel metal2 11144 7840 11144 7840 0 main.GATES_11.input2
rlabel metal2 5880 15484 5880 15484 0 main.GATES_110.input1
rlabel metal2 5656 6944 5656 6944 0 main.GATES_113.input1
rlabel metal2 3752 11536 3752 11536 0 main.GATES_114.input2
rlabel metal2 20440 11592 20440 11592 0 main.GATES_115.input2
rlabel metal2 11704 11760 11704 11760 0 main.GATES_116.input1
rlabel metal2 15400 14784 15400 14784 0 main.GATES_116.input3
rlabel metal2 5880 11368 5880 11368 0 main.GATES_119.result
rlabel metal3 16968 6440 16968 6440 0 main.GATES_124.input2
rlabel metal2 19880 11088 19880 11088 0 main.GATES_127.result
rlabel metal2 3976 17360 3976 17360 0 main.GATES_132.input1
rlabel metal3 19880 9688 19880 9688 0 main.GATES_15.input3
rlabel metal2 18256 19096 18256 19096 0 main.GATES_16.input1
rlabel metal2 20216 17248 20216 17248 0 main.GATES_18.result
rlabel metal3 14560 16072 14560 16072 0 main.GATES_19.input1
rlabel metal2 15288 15680 15288 15680 0 main.GATES_20.result
rlabel metal2 20216 7784 20216 7784 0 main.GATES_26.input3
rlabel metal2 21336 12376 21336 12376 0 main.GATES_29.input3
rlabel metal2 21000 16744 21000 16744 0 main.GATES_46.input3
rlabel metal3 21672 8120 21672 8120 0 net1
rlabel metal2 4312 10304 4312 10304 0 net10
rlabel metal3 8512 18984 8512 18984 0 net11
rlabel metal2 10136 19264 10136 19264 0 net12
rlabel metal2 18536 19656 18536 19656 0 net13
rlabel metal2 15568 19096 15568 19096 0 net14
rlabel metal2 17976 19880 17976 19880 0 net15
rlabel metal2 20664 15232 20664 15232 0 net16
rlabel metal2 21672 19600 21672 19600 0 net17
rlabel metal2 20832 9800 20832 9800 0 net2
rlabel metal3 21560 12152 21560 12152 0 net3
rlabel metal2 21896 16576 21896 16576 0 net4
rlabel metal2 22400 17416 22400 17416 0 net5
rlabel metal2 21896 5488 21896 5488 0 net6
rlabel metal2 19880 19936 19880 19936 0 net7
rlabel metal3 2744 13720 2744 13720 0 net8
rlabel metal2 4536 19712 4536 19712 0 net9
rlabel metal2 22232 4816 22232 4816 0 rst_n
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
