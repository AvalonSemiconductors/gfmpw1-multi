magic
tech gf180mcuD
magscale 1 10
timestamp 1702048942
<< metal1 >>
rect 8754 66782 8766 66834
rect 8818 66831 8830 66834
rect 9314 66831 9326 66834
rect 8818 66785 9326 66831
rect 8818 66782 8830 66785
rect 9314 66782 9326 66785
rect 9378 66782 9390 66834
rect 1344 66666 58576 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 58576 66666
rect 1344 66580 58576 66614
rect 26126 66498 26178 66510
rect 26126 66434 26178 66446
rect 40798 66498 40850 66510
rect 40798 66434 40850 66446
rect 43822 66498 43874 66510
rect 43822 66434 43874 66446
rect 48414 66498 48466 66510
rect 48414 66434 48466 66446
rect 52222 66498 52274 66510
rect 52222 66434 52274 66446
rect 56030 66498 56082 66510
rect 56030 66434 56082 66446
rect 18834 66334 18846 66386
rect 18898 66334 18910 66386
rect 22866 66334 22878 66386
rect 22930 66334 22942 66386
rect 36978 66334 36990 66386
rect 37042 66334 37054 66386
rect 17602 66222 17614 66274
rect 17666 66222 17678 66274
rect 23538 66222 23550 66274
rect 23602 66222 23614 66274
rect 25106 66222 25118 66274
rect 25170 66222 25182 66274
rect 39218 66222 39230 66274
rect 39282 66222 39294 66274
rect 39778 66222 39790 66274
rect 39842 66222 39854 66274
rect 46162 66222 46174 66274
rect 46226 66222 46238 66274
rect 47394 66222 47406 66274
rect 47458 66222 47470 66274
rect 51202 66222 51214 66274
rect 51266 66222 51278 66274
rect 55010 66222 55022 66274
rect 55074 66222 55086 66274
rect 2942 66162 2994 66174
rect 2942 66098 2994 66110
rect 5518 66162 5570 66174
rect 5518 66098 5570 66110
rect 6974 66162 7026 66174
rect 6974 66098 7026 66110
rect 9326 66162 9378 66174
rect 9326 66098 9378 66110
rect 11006 66162 11058 66174
rect 11006 66098 11058 66110
rect 13134 66162 13186 66174
rect 13134 66098 13186 66110
rect 15038 66162 15090 66174
rect 15038 66098 15090 66110
rect 17054 66162 17106 66174
rect 17054 66098 17106 66110
rect 29150 66162 29202 66174
rect 29150 66098 29202 66110
rect 31166 66162 31218 66174
rect 31166 66098 31218 66110
rect 33182 66162 33234 66174
rect 33182 66098 33234 66110
rect 35198 66162 35250 66174
rect 35198 66098 35250 66110
rect 43038 66162 43090 66174
rect 43038 66098 43090 66110
rect 1344 65882 58576 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 58576 65882
rect 1344 65796 58576 65830
rect 34862 65602 34914 65614
rect 34862 65538 34914 65550
rect 57822 65602 57874 65614
rect 57822 65538 57874 65550
rect 35534 65490 35586 65502
rect 57598 65490 57650 65502
rect 20178 65438 20190 65490
rect 20242 65438 20254 65490
rect 21858 65438 21870 65490
rect 21922 65438 21934 65490
rect 29698 65438 29710 65490
rect 29762 65438 29774 65490
rect 36642 65438 36654 65490
rect 36706 65438 36718 65490
rect 44370 65438 44382 65490
rect 44434 65438 44446 65490
rect 44818 65438 44830 65490
rect 44882 65438 44894 65490
rect 48850 65438 48862 65490
rect 48914 65438 48926 65490
rect 54898 65438 54910 65490
rect 54962 65438 54974 65490
rect 35534 65426 35586 65438
rect 57598 65426 57650 65438
rect 58158 65490 58210 65502
rect 58158 65426 58210 65438
rect 8878 65378 8930 65390
rect 8878 65314 8930 65326
rect 12462 65378 12514 65390
rect 20862 65378 20914 65390
rect 25454 65378 25506 65390
rect 17378 65326 17390 65378
rect 17442 65326 17454 65378
rect 19506 65326 19518 65378
rect 19570 65326 19582 65378
rect 22530 65326 22542 65378
rect 22594 65326 22606 65378
rect 24658 65326 24670 65378
rect 24722 65326 24734 65378
rect 12462 65314 12514 65326
rect 20862 65314 20914 65326
rect 25454 65314 25506 65326
rect 27358 65378 27410 65390
rect 27358 65314 27410 65326
rect 30270 65378 30322 65390
rect 30270 65314 30322 65326
rect 34974 65378 35026 65390
rect 40126 65378 40178 65390
rect 37426 65326 37438 65378
rect 37490 65326 37502 65378
rect 39554 65326 39566 65378
rect 39618 65326 39630 65378
rect 34974 65314 35026 65326
rect 40126 65314 40178 65326
rect 41134 65378 41186 65390
rect 55470 65378 55522 65390
rect 41570 65326 41582 65378
rect 41634 65326 41646 65378
rect 43698 65326 43710 65378
rect 43762 65326 43774 65378
rect 45602 65326 45614 65378
rect 45666 65326 45678 65378
rect 47730 65326 47742 65378
rect 47794 65326 47806 65378
rect 49522 65326 49534 65378
rect 49586 65326 49598 65378
rect 51650 65326 51662 65378
rect 51714 65326 51726 65378
rect 51986 65326 51998 65378
rect 52050 65326 52062 65378
rect 54114 65326 54126 65378
rect 54178 65326 54190 65378
rect 41134 65314 41186 65326
rect 55470 65314 55522 65326
rect 35086 65266 35138 65278
rect 35086 65202 35138 65214
rect 1344 65098 58576 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 58576 65098
rect 1344 65012 58576 65046
rect 23550 64930 23602 64942
rect 23550 64866 23602 64878
rect 42702 64930 42754 64942
rect 42702 64866 42754 64878
rect 47518 64930 47570 64942
rect 47518 64866 47570 64878
rect 50206 64930 50258 64942
rect 50206 64866 50258 64878
rect 51774 64930 51826 64942
rect 51774 64866 51826 64878
rect 44942 64818 44994 64830
rect 8530 64766 8542 64818
rect 8594 64766 8606 64818
rect 12114 64766 12126 64818
rect 12178 64766 12190 64818
rect 20738 64766 20750 64818
rect 20802 64766 20814 64818
rect 26898 64766 26910 64818
rect 26962 64766 26974 64818
rect 33506 64766 33518 64818
rect 33570 64766 33582 64818
rect 35634 64766 35646 64818
rect 35698 64766 35710 64818
rect 41346 64766 41358 64818
rect 41410 64766 41422 64818
rect 44942 64754 44994 64766
rect 45390 64818 45442 64830
rect 55234 64766 55246 64818
rect 55298 64766 55310 64818
rect 45390 64754 45442 64766
rect 27918 64706 27970 64718
rect 5730 64654 5742 64706
rect 5794 64654 5806 64706
rect 9314 64654 9326 64706
rect 9378 64654 9390 64706
rect 13458 64654 13470 64706
rect 13522 64654 13534 64706
rect 17938 64654 17950 64706
rect 18002 64654 18014 64706
rect 23986 64654 23998 64706
rect 24050 64654 24062 64706
rect 27918 64642 27970 64654
rect 29038 64706 29090 64718
rect 29038 64642 29090 64654
rect 29486 64706 29538 64718
rect 29486 64642 29538 64654
rect 30382 64706 30434 64718
rect 37102 64706 37154 64718
rect 36418 64654 36430 64706
rect 36482 64654 36494 64706
rect 38546 64654 38558 64706
rect 38610 64654 38622 64706
rect 41682 64654 41694 64706
rect 41746 64654 41758 64706
rect 49410 64654 49422 64706
rect 49474 64654 49486 64706
rect 54562 64654 54574 64706
rect 54626 64654 54638 64706
rect 58034 64654 58046 64706
rect 58098 64654 58110 64706
rect 30382 64642 30434 64654
rect 37102 64642 37154 64654
rect 12686 64594 12738 64606
rect 6402 64542 6414 64594
rect 6466 64542 6478 64594
rect 9986 64542 9998 64594
rect 10050 64542 10062 64594
rect 12686 64530 12738 64542
rect 13806 64594 13858 64606
rect 23662 64594 23714 64606
rect 30942 64594 30994 64606
rect 18610 64542 18622 64594
rect 18674 64542 18686 64594
rect 24770 64542 24782 64594
rect 24834 64542 24846 64594
rect 13806 64530 13858 64542
rect 23662 64530 23714 64542
rect 30942 64530 30994 64542
rect 32510 64594 32562 64606
rect 32510 64530 32562 64542
rect 32622 64594 32674 64606
rect 32622 64530 32674 64542
rect 32958 64594 33010 64606
rect 50318 64594 50370 64606
rect 39218 64542 39230 64594
rect 39282 64542 39294 64594
rect 32958 64530 33010 64542
rect 50318 64530 50370 64542
rect 51662 64594 51714 64606
rect 57362 64542 57374 64594
rect 57426 64542 57438 64594
rect 51662 64530 51714 64542
rect 12798 64482 12850 64494
rect 12798 64418 12850 64430
rect 13022 64482 13074 64494
rect 13022 64418 13074 64430
rect 13694 64482 13746 64494
rect 13694 64418 13746 64430
rect 21422 64482 21474 64494
rect 21422 64418 21474 64430
rect 23214 64482 23266 64494
rect 23214 64418 23266 64430
rect 27246 64482 27298 64494
rect 27246 64418 27298 64430
rect 27358 64482 27410 64494
rect 27358 64418 27410 64430
rect 27470 64482 27522 64494
rect 27470 64418 27522 64430
rect 28702 64482 28754 64494
rect 28702 64418 28754 64430
rect 29598 64482 29650 64494
rect 29598 64418 29650 64430
rect 29710 64482 29762 64494
rect 29710 64418 29762 64430
rect 30830 64482 30882 64494
rect 30830 64418 30882 64430
rect 31054 64482 31106 64494
rect 31054 64418 31106 64430
rect 31502 64482 31554 64494
rect 31502 64418 31554 64430
rect 32286 64482 32338 64494
rect 32286 64418 32338 64430
rect 33070 64482 33122 64494
rect 33070 64418 33122 64430
rect 33294 64482 33346 64494
rect 33294 64418 33346 64430
rect 52782 64482 52834 64494
rect 52782 64418 52834 64430
rect 54014 64482 54066 64494
rect 54014 64418 54066 64430
rect 54350 64482 54402 64494
rect 54350 64418 54402 64430
rect 1344 64314 58576 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 58576 64314
rect 1344 64228 58576 64262
rect 17614 64146 17666 64158
rect 12786 64094 12798 64146
rect 12850 64094 12862 64146
rect 17614 64082 17666 64094
rect 27806 64146 27858 64158
rect 27806 64082 27858 64094
rect 32286 64146 32338 64158
rect 32286 64082 32338 64094
rect 41582 64146 41634 64158
rect 41582 64082 41634 64094
rect 42030 64146 42082 64158
rect 42030 64082 42082 64094
rect 46734 64146 46786 64158
rect 46734 64082 46786 64094
rect 50430 64146 50482 64158
rect 50430 64082 50482 64094
rect 52334 64146 52386 64158
rect 52334 64082 52386 64094
rect 54574 64146 54626 64158
rect 54574 64082 54626 64094
rect 8542 64034 8594 64046
rect 17726 64034 17778 64046
rect 11442 63982 11454 64034
rect 11506 63982 11518 64034
rect 8542 63970 8594 63982
rect 17726 63970 17778 63982
rect 27470 64034 27522 64046
rect 27470 63970 27522 63982
rect 27582 64034 27634 64046
rect 46846 64034 46898 64046
rect 56030 64034 56082 64046
rect 31938 63982 31950 64034
rect 32002 63982 32014 64034
rect 35186 63982 35198 64034
rect 35250 63982 35262 64034
rect 50866 63982 50878 64034
rect 50930 64031 50942 64034
rect 51202 64031 51214 64034
rect 50930 63985 51214 64031
rect 50930 63982 50942 63985
rect 51202 63982 51214 63985
rect 51266 63982 51278 64034
rect 27582 63970 27634 63982
rect 46846 63970 46898 63982
rect 56030 63970 56082 63982
rect 56814 64034 56866 64046
rect 56814 63970 56866 63982
rect 16830 63922 16882 63934
rect 11778 63870 11790 63922
rect 11842 63870 11854 63922
rect 12450 63870 12462 63922
rect 12514 63870 12526 63922
rect 13570 63870 13582 63922
rect 13634 63870 13646 63922
rect 16830 63858 16882 63870
rect 17278 63922 17330 63934
rect 17278 63858 17330 63870
rect 17838 63922 17890 63934
rect 23438 63922 23490 63934
rect 32510 63922 32562 63934
rect 39454 63922 39506 63934
rect 43822 63922 43874 63934
rect 20178 63870 20190 63922
rect 20242 63870 20254 63922
rect 26674 63870 26686 63922
rect 26738 63870 26750 63922
rect 28018 63870 28030 63922
rect 28082 63870 28094 63922
rect 32050 63870 32062 63922
rect 32114 63870 32126 63922
rect 33506 63870 33518 63922
rect 33570 63870 33582 63922
rect 34626 63870 34638 63922
rect 34690 63870 34702 63922
rect 43362 63870 43374 63922
rect 43426 63870 43438 63922
rect 17838 63858 17890 63870
rect 23438 63858 23490 63870
rect 32510 63858 32562 63870
rect 39454 63858 39506 63870
rect 43822 63858 43874 63870
rect 46398 63922 46450 63934
rect 46398 63858 46450 63870
rect 47070 63922 47122 63934
rect 47070 63858 47122 63870
rect 49534 63922 49586 63934
rect 49534 63858 49586 63870
rect 49646 63922 49698 63934
rect 49646 63858 49698 63870
rect 49982 63922 50034 63934
rect 49982 63858 50034 63870
rect 50094 63922 50146 63934
rect 54126 63922 54178 63934
rect 51314 63870 51326 63922
rect 51378 63870 51390 63922
rect 50094 63858 50146 63870
rect 54126 63858 54178 63870
rect 54798 63922 54850 63934
rect 54798 63858 54850 63870
rect 27134 63810 27186 63822
rect 50430 63810 50482 63822
rect 14242 63758 14254 63810
rect 14306 63758 14318 63810
rect 16370 63758 16382 63810
rect 16434 63758 16446 63810
rect 20850 63758 20862 63810
rect 20914 63758 20926 63810
rect 22978 63758 22990 63810
rect 23042 63758 23054 63810
rect 26338 63758 26350 63810
rect 26402 63758 26414 63810
rect 28802 63758 28814 63810
rect 28866 63758 28878 63810
rect 30930 63758 30942 63810
rect 30994 63758 31006 63810
rect 31714 63758 31726 63810
rect 31778 63758 31790 63810
rect 33170 63758 33182 63810
rect 33234 63758 33246 63810
rect 27134 63746 27186 63758
rect 50430 63746 50482 63758
rect 50766 63810 50818 63822
rect 50766 63746 50818 63758
rect 54686 63810 54738 63822
rect 54686 63746 54738 63758
rect 8430 63698 8482 63710
rect 8430 63634 8482 63646
rect 43038 63698 43090 63710
rect 43038 63634 43090 63646
rect 43374 63698 43426 63710
rect 43374 63634 43426 63646
rect 56590 63698 56642 63710
rect 56590 63634 56642 63646
rect 56926 63698 56978 63710
rect 56926 63634 56978 63646
rect 1344 63530 58576 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 58576 63530
rect 1344 63444 58576 63478
rect 12014 63362 12066 63374
rect 12014 63298 12066 63310
rect 12350 63362 12402 63374
rect 12350 63298 12402 63310
rect 12686 63362 12738 63374
rect 12686 63298 12738 63310
rect 19630 63362 19682 63374
rect 19630 63298 19682 63310
rect 22318 63362 22370 63374
rect 22318 63298 22370 63310
rect 31278 63362 31330 63374
rect 31278 63298 31330 63310
rect 53566 63362 53618 63374
rect 54450 63310 54462 63362
rect 54514 63310 54526 63362
rect 53566 63298 53618 63310
rect 6638 63250 6690 63262
rect 6638 63186 6690 63198
rect 11902 63250 11954 63262
rect 11902 63186 11954 63198
rect 17502 63250 17554 63262
rect 17502 63186 17554 63198
rect 26238 63250 26290 63262
rect 45166 63250 45218 63262
rect 32050 63198 32062 63250
rect 32114 63198 32126 63250
rect 26238 63186 26290 63198
rect 45166 63186 45218 63198
rect 47742 63250 47794 63262
rect 47742 63186 47794 63198
rect 51438 63250 51490 63262
rect 51438 63186 51490 63198
rect 51662 63250 51714 63262
rect 51662 63186 51714 63198
rect 53006 63250 53058 63262
rect 53006 63186 53058 63198
rect 53902 63250 53954 63262
rect 53902 63186 53954 63198
rect 54910 63250 54962 63262
rect 55234 63198 55246 63250
rect 55298 63198 55310 63250
rect 57362 63198 57374 63250
rect 57426 63198 57438 63250
rect 54910 63186 54962 63198
rect 6750 63138 6802 63150
rect 26686 63138 26738 63150
rect 7858 63086 7870 63138
rect 7922 63086 7934 63138
rect 8082 63086 8094 63138
rect 8146 63086 8158 63138
rect 15474 63086 15486 63138
rect 15538 63086 15550 63138
rect 16258 63086 16270 63138
rect 16322 63086 16334 63138
rect 19618 63086 19630 63138
rect 19682 63086 19694 63138
rect 21298 63086 21310 63138
rect 21362 63086 21374 63138
rect 6750 63074 6802 63086
rect 26686 63074 26738 63086
rect 27134 63138 27186 63150
rect 27806 63138 27858 63150
rect 27570 63086 27582 63138
rect 27634 63086 27646 63138
rect 27134 63074 27186 63086
rect 27806 63074 27858 63086
rect 28142 63138 28194 63150
rect 30382 63138 30434 63150
rect 43486 63138 43538 63150
rect 30146 63086 30158 63138
rect 30210 63086 30222 63138
rect 32162 63086 32174 63138
rect 32226 63086 32238 63138
rect 32386 63086 32398 63138
rect 32450 63086 32462 63138
rect 41234 63086 41246 63138
rect 41298 63086 41310 63138
rect 28142 63074 28194 63086
rect 30382 63074 30434 63086
rect 43486 63074 43538 63086
rect 44046 63138 44098 63150
rect 44046 63074 44098 63086
rect 44942 63138 44994 63150
rect 50654 63138 50706 63150
rect 46050 63086 46062 63138
rect 46114 63086 46126 63138
rect 46498 63086 46510 63138
rect 46562 63086 46574 63138
rect 44942 63074 44994 63086
rect 50654 63074 50706 63086
rect 50766 63138 50818 63150
rect 50766 63074 50818 63086
rect 51102 63138 51154 63150
rect 51102 63074 51154 63086
rect 51214 63138 51266 63150
rect 51214 63074 51266 63086
rect 51774 63138 51826 63150
rect 51774 63074 51826 63086
rect 53230 63138 53282 63150
rect 53230 63074 53282 63086
rect 54126 63138 54178 63150
rect 58034 63086 58046 63138
rect 58098 63086 58110 63138
rect 54126 63074 54178 63086
rect 6526 63026 6578 63038
rect 6526 62962 6578 62974
rect 7086 63026 7138 63038
rect 7086 62962 7138 62974
rect 7646 63026 7698 63038
rect 7646 62962 7698 62974
rect 14814 63026 14866 63038
rect 17614 63026 17666 63038
rect 16370 62974 16382 63026
rect 16434 62974 16446 63026
rect 14814 62962 14866 62974
rect 17614 62962 17666 62974
rect 19966 63026 20018 63038
rect 19966 62962 20018 62974
rect 26126 63026 26178 63038
rect 26126 62962 26178 62974
rect 26462 63026 26514 63038
rect 26462 62962 26514 62974
rect 28030 63026 28082 63038
rect 28030 62962 28082 62974
rect 29486 63026 29538 63038
rect 29486 62962 29538 62974
rect 31166 63026 31218 63038
rect 31166 62962 31218 62974
rect 31278 63026 31330 63038
rect 31278 62962 31330 62974
rect 31950 63026 32002 63038
rect 44158 63026 44210 63038
rect 41010 62974 41022 63026
rect 41074 62974 41086 63026
rect 42242 62974 42254 63026
rect 42306 62974 42318 63026
rect 31950 62962 32002 62974
rect 44158 62962 44210 62974
rect 45054 63026 45106 63038
rect 45054 62962 45106 62974
rect 45502 63026 45554 63038
rect 45502 62962 45554 62974
rect 45838 63026 45890 63038
rect 45838 62962 45890 62974
rect 12462 62914 12514 62926
rect 12462 62850 12514 62862
rect 13694 62914 13746 62926
rect 13694 62850 13746 62862
rect 17390 62914 17442 62926
rect 17390 62850 17442 62862
rect 17838 62914 17890 62926
rect 17838 62850 17890 62862
rect 18510 62914 18562 62926
rect 18510 62850 18562 62862
rect 27022 62914 27074 62926
rect 27022 62850 27074 62862
rect 27246 62914 27298 62926
rect 27246 62850 27298 62862
rect 28590 62914 28642 62926
rect 28590 62850 28642 62862
rect 32846 62914 32898 62926
rect 42926 62914 42978 62926
rect 42466 62862 42478 62914
rect 42530 62862 42542 62914
rect 32846 62850 32898 62862
rect 42926 62850 42978 62862
rect 44382 62914 44434 62926
rect 44382 62850 44434 62862
rect 45278 62914 45330 62926
rect 45278 62850 45330 62862
rect 47182 62914 47234 62926
rect 47182 62850 47234 62862
rect 1344 62746 58576 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 58576 62746
rect 1344 62660 58576 62694
rect 7198 62578 7250 62590
rect 7198 62514 7250 62526
rect 7310 62578 7362 62590
rect 7310 62514 7362 62526
rect 7982 62578 8034 62590
rect 14926 62578 14978 62590
rect 13906 62526 13918 62578
rect 13970 62526 13982 62578
rect 7982 62514 8034 62526
rect 14926 62514 14978 62526
rect 16494 62578 16546 62590
rect 16494 62514 16546 62526
rect 16718 62578 16770 62590
rect 16718 62514 16770 62526
rect 19406 62578 19458 62590
rect 19406 62514 19458 62526
rect 19966 62578 20018 62590
rect 19966 62514 20018 62526
rect 29038 62578 29090 62590
rect 29038 62514 29090 62526
rect 44046 62578 44098 62590
rect 44046 62514 44098 62526
rect 44718 62578 44770 62590
rect 44718 62514 44770 62526
rect 45502 62578 45554 62590
rect 45502 62514 45554 62526
rect 45614 62578 45666 62590
rect 45614 62514 45666 62526
rect 47182 62578 47234 62590
rect 47182 62514 47234 62526
rect 52110 62578 52162 62590
rect 52110 62514 52162 62526
rect 6862 62466 6914 62478
rect 6862 62402 6914 62414
rect 8542 62466 8594 62478
rect 14814 62466 14866 62478
rect 10882 62414 10894 62466
rect 10946 62414 10958 62466
rect 13122 62414 13134 62466
rect 13186 62414 13198 62466
rect 8542 62402 8594 62414
rect 14814 62402 14866 62414
rect 18958 62466 19010 62478
rect 18958 62402 19010 62414
rect 28926 62466 28978 62478
rect 28926 62402 28978 62414
rect 37886 62466 37938 62478
rect 37886 62402 37938 62414
rect 39454 62466 39506 62478
rect 39454 62402 39506 62414
rect 41918 62466 41970 62478
rect 41918 62402 41970 62414
rect 43262 62466 43314 62478
rect 43262 62402 43314 62414
rect 47294 62466 47346 62478
rect 47294 62402 47346 62414
rect 52446 62466 52498 62478
rect 52446 62402 52498 62414
rect 56926 62466 56978 62478
rect 56926 62402 56978 62414
rect 57374 62466 57426 62478
rect 57374 62402 57426 62414
rect 7086 62354 7138 62366
rect 7086 62290 7138 62302
rect 7870 62354 7922 62366
rect 7870 62290 7922 62302
rect 8206 62354 8258 62366
rect 8206 62290 8258 62302
rect 8430 62354 8482 62366
rect 8430 62290 8482 62302
rect 8766 62354 8818 62366
rect 16382 62354 16434 62366
rect 9426 62302 9438 62354
rect 9490 62302 9502 62354
rect 10210 62302 10222 62354
rect 10274 62302 10286 62354
rect 12898 62302 12910 62354
rect 12962 62302 12974 62354
rect 13794 62302 13806 62354
rect 13858 62302 13870 62354
rect 15138 62302 15150 62354
rect 15202 62302 15214 62354
rect 8766 62290 8818 62302
rect 16382 62290 16434 62302
rect 19182 62354 19234 62366
rect 19182 62290 19234 62302
rect 19518 62354 19570 62366
rect 19518 62290 19570 62302
rect 19854 62354 19906 62366
rect 19854 62290 19906 62302
rect 20078 62354 20130 62366
rect 29150 62354 29202 62366
rect 20402 62302 20414 62354
rect 20466 62302 20478 62354
rect 20078 62290 20130 62302
rect 29150 62290 29202 62302
rect 29374 62354 29426 62366
rect 43486 62354 43538 62366
rect 37202 62302 37214 62354
rect 37266 62302 37278 62354
rect 38770 62302 38782 62354
rect 38834 62302 38846 62354
rect 41234 62302 41246 62354
rect 41298 62302 41310 62354
rect 42802 62302 42814 62354
rect 42866 62302 42878 62354
rect 29374 62290 29426 62302
rect 43486 62290 43538 62302
rect 43934 62354 43986 62366
rect 43934 62290 43986 62302
rect 44158 62354 44210 62366
rect 44158 62290 44210 62302
rect 44606 62354 44658 62366
rect 44606 62290 44658 62302
rect 44942 62354 44994 62366
rect 44942 62290 44994 62302
rect 45054 62354 45106 62366
rect 45054 62290 45106 62302
rect 45726 62354 45778 62366
rect 45726 62290 45778 62302
rect 45950 62354 46002 62366
rect 45950 62290 46002 62302
rect 46286 62354 46338 62366
rect 46286 62290 46338 62302
rect 46510 62354 46562 62366
rect 57150 62354 57202 62366
rect 46946 62302 46958 62354
rect 47010 62302 47022 62354
rect 48850 62302 48862 62354
rect 48914 62302 48926 62354
rect 53442 62302 53454 62354
rect 53506 62302 53518 62354
rect 56690 62302 56702 62354
rect 56754 62302 56766 62354
rect 46510 62290 46562 62302
rect 57150 62290 57202 62302
rect 57486 62354 57538 62366
rect 57486 62290 57538 62302
rect 15598 62242 15650 62254
rect 10546 62190 10558 62242
rect 10610 62190 10622 62242
rect 15598 62178 15650 62190
rect 20862 62242 20914 62254
rect 20862 62178 20914 62190
rect 27694 62242 27746 62254
rect 27694 62178 27746 62190
rect 30830 62242 30882 62254
rect 30830 62178 30882 62190
rect 31278 62242 31330 62254
rect 46174 62242 46226 62254
rect 37538 62190 37550 62242
rect 37602 62190 37614 62242
rect 38546 62190 38558 62242
rect 38610 62190 38622 62242
rect 41010 62190 41022 62242
rect 41074 62190 41086 62242
rect 42466 62190 42478 62242
rect 42530 62190 42542 62242
rect 49522 62190 49534 62242
rect 49586 62190 49598 62242
rect 51650 62190 51662 62242
rect 51714 62190 51726 62242
rect 52882 62190 52894 62242
rect 52946 62190 52958 62242
rect 55346 62190 55358 62242
rect 55410 62190 55422 62242
rect 31278 62178 31330 62190
rect 46174 62178 46226 62190
rect 1344 61962 58576 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 58576 61962
rect 1344 61876 58576 61910
rect 20302 61794 20354 61806
rect 20302 61730 20354 61742
rect 38222 61794 38274 61806
rect 38222 61730 38274 61742
rect 43374 61794 43426 61806
rect 43374 61730 43426 61742
rect 49198 61794 49250 61806
rect 49198 61730 49250 61742
rect 56366 61794 56418 61806
rect 56366 61730 56418 61742
rect 7534 61682 7586 61694
rect 7534 61618 7586 61630
rect 12238 61682 12290 61694
rect 35870 61682 35922 61694
rect 24546 61630 24558 61682
rect 24610 61630 24622 61682
rect 12238 61618 12290 61630
rect 35870 61618 35922 61630
rect 37438 61682 37490 61694
rect 52770 61630 52782 61682
rect 52834 61630 52846 61682
rect 55010 61630 55022 61682
rect 55074 61630 55086 61682
rect 37438 61618 37490 61630
rect 21746 61518 21758 61570
rect 21810 61518 21822 61570
rect 35634 61518 35646 61570
rect 35698 61518 35710 61570
rect 38546 61518 38558 61570
rect 38610 61518 38622 61570
rect 43362 61518 43374 61570
rect 43426 61518 43438 61570
rect 53106 61518 53118 61570
rect 53170 61518 53182 61570
rect 54338 61518 54350 61570
rect 54402 61518 54414 61570
rect 55458 61518 55470 61570
rect 55522 61518 55534 61570
rect 6414 61458 6466 61470
rect 6414 61394 6466 61406
rect 6750 61458 6802 61470
rect 6750 61394 6802 61406
rect 19966 61458 20018 61470
rect 24894 61458 24946 61470
rect 20402 61406 20414 61458
rect 20466 61455 20478 61458
rect 20626 61455 20638 61458
rect 20466 61409 20638 61455
rect 20466 61406 20478 61409
rect 20626 61406 20638 61409
rect 20690 61406 20702 61458
rect 22418 61406 22430 61458
rect 22482 61406 22494 61458
rect 19966 61394 20018 61406
rect 24894 61394 24946 61406
rect 32734 61458 32786 61470
rect 32734 61394 32786 61406
rect 34414 61458 34466 61470
rect 34414 61394 34466 61406
rect 34974 61458 35026 61470
rect 34974 61394 35026 61406
rect 35982 61458 36034 61470
rect 35982 61394 36034 61406
rect 36990 61458 37042 61470
rect 36990 61394 37042 61406
rect 37214 61458 37266 61470
rect 37214 61394 37266 61406
rect 37550 61458 37602 61470
rect 37550 61394 37602 61406
rect 43710 61458 43762 61470
rect 43710 61394 43762 61406
rect 49086 61458 49138 61470
rect 49086 61394 49138 61406
rect 6190 61346 6242 61358
rect 6190 61282 6242 61294
rect 6302 61346 6354 61358
rect 6302 61282 6354 61294
rect 6862 61346 6914 61358
rect 6862 61282 6914 61294
rect 7086 61346 7138 61358
rect 7086 61282 7138 61294
rect 20190 61346 20242 61358
rect 20190 61282 20242 61294
rect 20750 61346 20802 61358
rect 20750 61282 20802 61294
rect 25006 61346 25058 61358
rect 25006 61282 25058 61294
rect 25566 61346 25618 61358
rect 25566 61282 25618 61294
rect 25902 61346 25954 61358
rect 25902 61282 25954 61294
rect 32398 61346 32450 61358
rect 32398 61282 32450 61294
rect 32622 61346 32674 61358
rect 32622 61282 32674 61294
rect 34526 61346 34578 61358
rect 34526 61282 34578 61294
rect 34750 61346 34802 61358
rect 34750 61282 34802 61294
rect 35086 61346 35138 61358
rect 35086 61282 35138 61294
rect 35198 61346 35250 61358
rect 35198 61282 35250 61294
rect 38334 61346 38386 61358
rect 38334 61282 38386 61294
rect 44942 61346 44994 61358
rect 44942 61282 44994 61294
rect 1344 61178 58576 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 58576 61178
rect 1344 61092 58576 61126
rect 25454 61010 25506 61022
rect 7858 60958 7870 61010
rect 7922 60958 7934 61010
rect 25454 60946 25506 60958
rect 26014 61010 26066 61022
rect 37326 61010 37378 61022
rect 42702 61010 42754 61022
rect 32274 60958 32286 61010
rect 32338 60958 32350 61010
rect 40002 60958 40014 61010
rect 40066 60958 40078 61010
rect 26014 60946 26066 60958
rect 37326 60946 37378 60958
rect 42702 60946 42754 60958
rect 49086 61010 49138 61022
rect 49086 60946 49138 60958
rect 49646 61010 49698 61022
rect 57934 61010 57986 61022
rect 50978 60958 50990 61010
rect 51042 60958 51054 61010
rect 57026 60958 57038 61010
rect 57090 60958 57102 61010
rect 49646 60946 49698 60958
rect 57934 60946 57986 60958
rect 11006 60898 11058 60910
rect 6290 60846 6302 60898
rect 6354 60846 6366 60898
rect 11006 60834 11058 60846
rect 13022 60898 13074 60910
rect 13022 60834 13074 60846
rect 13246 60898 13298 60910
rect 13246 60834 13298 60846
rect 17502 60898 17554 60910
rect 17502 60834 17554 60846
rect 17950 60898 18002 60910
rect 17950 60834 18002 60846
rect 18062 60898 18114 60910
rect 27246 60898 27298 60910
rect 20962 60846 20974 60898
rect 21026 60846 21038 60898
rect 18062 60834 18114 60846
rect 27246 60834 27298 60846
rect 27806 60898 27858 60910
rect 27806 60834 27858 60846
rect 29598 60898 29650 60910
rect 29598 60834 29650 60846
rect 35422 60898 35474 60910
rect 35422 60834 35474 60846
rect 36766 60898 36818 60910
rect 57374 60898 57426 60910
rect 39106 60846 39118 60898
rect 39170 60846 39182 60898
rect 54450 60846 54462 60898
rect 54514 60846 54526 60898
rect 55794 60846 55806 60898
rect 55858 60846 55870 60898
rect 57138 60846 57150 60898
rect 57202 60846 57214 60898
rect 36766 60834 36818 60846
rect 57374 60834 57426 60846
rect 10782 60786 10834 60798
rect 13358 60786 13410 60798
rect 2818 60734 2830 60786
rect 2882 60734 2894 60786
rect 6738 60734 6750 60786
rect 6802 60734 6814 60786
rect 7522 60734 7534 60786
rect 7586 60734 7598 60786
rect 11554 60734 11566 60786
rect 11618 60734 11630 60786
rect 11890 60734 11902 60786
rect 11954 60734 11966 60786
rect 12562 60734 12574 60786
rect 12626 60734 12638 60786
rect 10782 60722 10834 60734
rect 13358 60722 13410 60734
rect 17390 60786 17442 60798
rect 17390 60722 17442 60734
rect 17726 60786 17778 60798
rect 25902 60786 25954 60798
rect 21746 60734 21758 60786
rect 21810 60734 21822 60786
rect 22642 60734 22654 60786
rect 22706 60734 22718 60786
rect 17726 60722 17778 60734
rect 25902 60722 25954 60734
rect 26238 60786 26290 60798
rect 26238 60722 26290 60734
rect 27134 60786 27186 60798
rect 27134 60722 27186 60734
rect 27470 60786 27522 60798
rect 27470 60722 27522 60734
rect 27694 60786 27746 60798
rect 27694 60722 27746 60734
rect 27918 60786 27970 60798
rect 27918 60722 27970 60734
rect 28366 60786 28418 60798
rect 31950 60786 32002 60798
rect 35870 60786 35922 60798
rect 41358 60786 41410 60798
rect 50094 60786 50146 60798
rect 53006 60786 53058 60798
rect 57710 60786 57762 60798
rect 28914 60734 28926 60786
rect 28978 60734 28990 60786
rect 33394 60734 33406 60786
rect 33458 60734 33470 60786
rect 34738 60734 34750 60786
rect 34802 60734 34814 60786
rect 36082 60734 36094 60786
rect 36146 60734 36158 60786
rect 37762 60734 37774 60786
rect 37826 60734 37838 60786
rect 38994 60734 39006 60786
rect 39058 60734 39070 60786
rect 39890 60734 39902 60786
rect 39954 60734 39966 60786
rect 42466 60734 42478 60786
rect 42530 60734 42542 60786
rect 48850 60734 48862 60786
rect 48914 60734 48926 60786
rect 49298 60734 49310 60786
rect 49362 60734 49374 60786
rect 49634 60734 49646 60786
rect 49698 60734 49710 60786
rect 51202 60734 51214 60786
rect 51266 60734 51278 60786
rect 53330 60734 53342 60786
rect 53394 60734 53406 60786
rect 54674 60734 54686 60786
rect 54738 60734 54750 60786
rect 56690 60734 56702 60786
rect 56754 60734 56766 60786
rect 28366 60722 28418 60734
rect 31950 60722 32002 60734
rect 35870 60722 35922 60734
rect 41358 60722 41410 60734
rect 50094 60722 50146 60734
rect 53006 60722 53058 60734
rect 57710 60722 57762 60734
rect 13918 60674 13970 60686
rect 3490 60622 3502 60674
rect 3554 60622 3566 60674
rect 5618 60622 5630 60674
rect 5682 60622 5694 60674
rect 11106 60622 11118 60674
rect 11170 60622 11182 60674
rect 12674 60622 12686 60674
rect 12738 60622 12750 60674
rect 13918 60610 13970 60622
rect 14254 60674 14306 60686
rect 30046 60674 30098 60686
rect 18834 60622 18846 60674
rect 18898 60622 18910 60674
rect 23202 60622 23214 60674
rect 23266 60622 23278 60674
rect 28690 60622 28702 60674
rect 28754 60622 28766 60674
rect 14254 60610 14306 60622
rect 30046 60610 30098 60622
rect 30494 60674 30546 60686
rect 30494 60610 30546 60622
rect 31614 60674 31666 60686
rect 34078 60674 34130 60686
rect 38558 60674 38610 60686
rect 33170 60622 33182 60674
rect 33234 60622 33246 60674
rect 34514 60622 34526 60674
rect 34578 60622 34590 60674
rect 37874 60622 37886 60674
rect 37938 60622 37950 60674
rect 31614 60610 31666 60622
rect 34078 60610 34130 60622
rect 38558 60610 38610 60622
rect 41918 60674 41970 60686
rect 41918 60610 41970 60622
rect 49758 60674 49810 60686
rect 49758 60610 49810 60622
rect 56030 60674 56082 60686
rect 56030 60610 56082 60622
rect 18062 60562 18114 60574
rect 18062 60498 18114 60510
rect 25230 60562 25282 60574
rect 25230 60498 25282 60510
rect 25566 60562 25618 60574
rect 25566 60498 25618 60510
rect 29934 60562 29986 60574
rect 29934 60498 29986 60510
rect 41470 60562 41522 60574
rect 41470 60498 41522 60510
rect 42814 60562 42866 60574
rect 42814 60498 42866 60510
rect 56926 60562 56978 60574
rect 56926 60498 56978 60510
rect 58046 60562 58098 60574
rect 58046 60498 58098 60510
rect 1344 60394 58576 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 58576 60394
rect 1344 60308 58576 60342
rect 22654 60226 22706 60238
rect 6962 60174 6974 60226
rect 7026 60174 7038 60226
rect 17602 60174 17614 60226
rect 17666 60174 17678 60226
rect 18946 60174 18958 60226
rect 19010 60174 19022 60226
rect 22654 60162 22706 60174
rect 28366 60226 28418 60238
rect 28366 60162 28418 60174
rect 32510 60226 32562 60238
rect 32510 60162 32562 60174
rect 34414 60226 34466 60238
rect 44270 60226 44322 60238
rect 34738 60174 34750 60226
rect 34802 60174 34814 60226
rect 34414 60162 34466 60174
rect 44270 60162 44322 60174
rect 5854 60114 5906 60126
rect 15710 60114 15762 60126
rect 27806 60114 27858 60126
rect 9090 60062 9102 60114
rect 9154 60062 9166 60114
rect 11218 60062 11230 60114
rect 11282 60062 11294 60114
rect 11778 60062 11790 60114
rect 11842 60062 11854 60114
rect 17154 60062 17166 60114
rect 17218 60062 17230 60114
rect 25442 60062 25454 60114
rect 25506 60062 25518 60114
rect 5854 60050 5906 60062
rect 15710 60050 15762 60062
rect 27806 60050 27858 60062
rect 32062 60114 32114 60126
rect 32062 60050 32114 60062
rect 34190 60114 34242 60126
rect 34190 60050 34242 60062
rect 38670 60114 38722 60126
rect 54910 60114 54962 60126
rect 42466 60062 42478 60114
rect 42530 60062 42542 60114
rect 49858 60062 49870 60114
rect 49922 60062 49934 60114
rect 55234 60062 55246 60114
rect 55298 60062 55310 60114
rect 38670 60050 38722 60062
rect 54910 60050 54962 60062
rect 12910 60002 12962 60014
rect 16494 60002 16546 60014
rect 19854 60002 19906 60014
rect 28030 60002 28082 60014
rect 6514 59950 6526 60002
rect 6578 59950 6590 60002
rect 7074 59950 7086 60002
rect 7138 59950 7150 60002
rect 7410 59950 7422 60002
rect 7474 59950 7486 60002
rect 8418 59950 8430 60002
rect 8482 59950 8494 60002
rect 11666 59950 11678 60002
rect 11730 59950 11742 60002
rect 12450 59950 12462 60002
rect 12514 59950 12526 60002
rect 14130 59950 14142 60002
rect 14194 59950 14206 60002
rect 15250 59950 15262 60002
rect 15314 59950 15326 60002
rect 16930 59950 16942 60002
rect 16994 59950 17006 60002
rect 18834 59950 18846 60002
rect 18898 59950 18910 60002
rect 20178 59950 20190 60002
rect 20242 59950 20254 60002
rect 23986 59950 23998 60002
rect 24050 59950 24062 60002
rect 25890 59950 25902 60002
rect 25954 59950 25966 60002
rect 26450 59950 26462 60002
rect 26514 59950 26526 60002
rect 12910 59938 12962 59950
rect 16494 59938 16546 59950
rect 19854 59938 19906 59950
rect 28030 59938 28082 59950
rect 29038 60002 29090 60014
rect 29038 59938 29090 59950
rect 29374 60002 29426 60014
rect 29374 59938 29426 59950
rect 31166 60002 31218 60014
rect 32846 60002 32898 60014
rect 31378 59950 31390 60002
rect 31442 59950 31454 60002
rect 31166 59938 31218 59950
rect 32846 59938 32898 59950
rect 33630 60002 33682 60014
rect 33630 59938 33682 59950
rect 40798 60002 40850 60014
rect 50990 60002 51042 60014
rect 41682 59950 41694 60002
rect 41746 59950 41758 60002
rect 47058 59950 47070 60002
rect 47122 59950 47134 60002
rect 40798 59938 40850 59950
rect 50990 59938 51042 59950
rect 51214 60002 51266 60014
rect 51886 60002 51938 60014
rect 51650 59950 51662 60002
rect 51714 59950 51726 60002
rect 51214 59938 51266 59950
rect 51886 59938 51938 59950
rect 52110 60002 52162 60014
rect 58034 59950 58046 60002
rect 58098 59950 58110 60002
rect 52110 59938 52162 59950
rect 12014 59890 12066 59902
rect 16158 59890 16210 59902
rect 13794 59838 13806 59890
rect 13858 59838 13870 59890
rect 12014 59826 12066 59838
rect 16158 59826 16210 59838
rect 16270 59890 16322 59902
rect 16270 59826 16322 59838
rect 22990 59890 23042 59902
rect 22990 59826 23042 59838
rect 23326 59890 23378 59902
rect 29262 59890 29314 59902
rect 24882 59838 24894 59890
rect 24946 59838 24958 59890
rect 26562 59838 26574 59890
rect 26626 59838 26638 59890
rect 23326 59826 23378 59838
rect 29262 59826 29314 59838
rect 32398 59890 32450 59902
rect 32398 59826 32450 59838
rect 33070 59890 33122 59902
rect 33070 59826 33122 59838
rect 33182 59890 33234 59902
rect 33182 59826 33234 59838
rect 44158 59890 44210 59902
rect 47730 59838 47742 59890
rect 47794 59838 47806 59890
rect 50194 59838 50206 59890
rect 50258 59838 50270 59890
rect 57362 59838 57374 59890
rect 57426 59838 57438 59890
rect 44158 59826 44210 59838
rect 21982 59778 22034 59790
rect 21982 59714 22034 59726
rect 22766 59778 22818 59790
rect 27470 59778 27522 59790
rect 30718 59778 30770 59790
rect 26002 59726 26014 59778
rect 26066 59726 26078 59778
rect 30370 59726 30382 59778
rect 30434 59726 30446 59778
rect 22766 59714 22818 59726
rect 27470 59714 27522 59726
rect 30718 59714 30770 59726
rect 32510 59778 32562 59790
rect 32510 59714 32562 59726
rect 40014 59778 40066 59790
rect 40014 59714 40066 59726
rect 40462 59778 40514 59790
rect 40462 59714 40514 59726
rect 40686 59778 40738 59790
rect 40686 59714 40738 59726
rect 40910 59778 40962 59790
rect 40910 59714 40962 59726
rect 50542 59778 50594 59790
rect 50542 59714 50594 59726
rect 51102 59778 51154 59790
rect 51986 59726 51998 59778
rect 52050 59726 52062 59778
rect 51102 59714 51154 59726
rect 1344 59610 58576 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 58576 59610
rect 1344 59524 58576 59558
rect 7646 59442 7698 59454
rect 7646 59378 7698 59390
rect 11342 59442 11394 59454
rect 11342 59378 11394 59390
rect 15038 59442 15090 59454
rect 15038 59378 15090 59390
rect 15150 59442 15202 59454
rect 42254 59442 42306 59454
rect 15698 59390 15710 59442
rect 15762 59390 15774 59442
rect 16706 59390 16718 59442
rect 16770 59390 16782 59442
rect 27010 59390 27022 59442
rect 27074 59390 27086 59442
rect 15150 59378 15202 59390
rect 42254 59378 42306 59390
rect 48078 59442 48130 59454
rect 48078 59378 48130 59390
rect 48862 59442 48914 59454
rect 48862 59378 48914 59390
rect 48974 59442 49026 59454
rect 48974 59378 49026 59390
rect 49534 59442 49586 59454
rect 49534 59378 49586 59390
rect 50430 59442 50482 59454
rect 50430 59378 50482 59390
rect 54686 59442 54738 59454
rect 54686 59378 54738 59390
rect 56030 59442 56082 59454
rect 56030 59378 56082 59390
rect 56814 59442 56866 59454
rect 56814 59378 56866 59390
rect 7534 59330 7586 59342
rect 7534 59266 7586 59278
rect 7758 59330 7810 59342
rect 7758 59266 7810 59278
rect 8206 59330 8258 59342
rect 41470 59330 41522 59342
rect 17602 59278 17614 59330
rect 17666 59278 17678 59330
rect 35634 59278 35646 59330
rect 35698 59278 35710 59330
rect 8206 59266 8258 59278
rect 41470 59266 41522 59278
rect 42366 59330 42418 59342
rect 42366 59266 42418 59278
rect 43038 59330 43090 59342
rect 43038 59266 43090 59278
rect 48190 59330 48242 59342
rect 48190 59266 48242 59278
rect 56926 59330 56978 59342
rect 56926 59266 56978 59278
rect 14478 59218 14530 59230
rect 12226 59166 12238 59218
rect 12290 59166 12302 59218
rect 14478 59154 14530 59166
rect 14926 59218 14978 59230
rect 27358 59218 27410 59230
rect 37102 59218 37154 59230
rect 40798 59218 40850 59230
rect 15922 59166 15934 59218
rect 15986 59166 15998 59218
rect 16482 59166 16494 59218
rect 16546 59166 16558 59218
rect 17714 59166 17726 59218
rect 17778 59166 17790 59218
rect 36530 59166 36542 59218
rect 36594 59166 36606 59218
rect 39890 59166 39902 59218
rect 39954 59166 39966 59218
rect 14926 59154 14978 59166
rect 27358 59154 27410 59166
rect 37102 59154 37154 59166
rect 40798 59154 40850 59166
rect 41246 59218 41298 59230
rect 41246 59154 41298 59166
rect 42030 59218 42082 59230
rect 42030 59154 42082 59166
rect 42142 59218 42194 59230
rect 42926 59218 42978 59230
rect 42578 59166 42590 59218
rect 42642 59166 42654 59218
rect 42142 59154 42194 59166
rect 42926 59154 42978 59166
rect 43262 59218 43314 59230
rect 49310 59218 49362 59230
rect 45266 59166 45278 59218
rect 45330 59166 45342 59218
rect 43262 59154 43314 59166
rect 49310 59154 49362 59166
rect 49422 59218 49474 59230
rect 49422 59154 49474 59166
rect 49982 59218 50034 59230
rect 58158 59218 58210 59230
rect 51426 59166 51438 59218
rect 51490 59166 51502 59218
rect 56578 59166 56590 59218
rect 56642 59166 56654 59218
rect 49982 59154 50034 59166
rect 58158 59154 58210 59166
rect 1822 59106 1874 59118
rect 27806 59106 27858 59118
rect 12786 59054 12798 59106
rect 12850 59054 12862 59106
rect 18050 59054 18062 59106
rect 18114 59054 18126 59106
rect 1822 59042 1874 59054
rect 27806 59042 27858 59054
rect 30942 59106 30994 59118
rect 30942 59042 30994 59054
rect 32286 59106 32338 59118
rect 40350 59106 40402 59118
rect 39442 59054 39454 59106
rect 39506 59054 39518 59106
rect 32286 59042 32338 59054
rect 40350 59042 40402 59054
rect 41022 59106 41074 59118
rect 41022 59042 41074 59054
rect 45726 59106 45778 59118
rect 45726 59042 45778 59054
rect 49646 59106 49698 59118
rect 55582 59106 55634 59118
rect 52098 59054 52110 59106
rect 52162 59054 52174 59106
rect 54226 59054 54238 59106
rect 54290 59054 54302 59106
rect 57698 59054 57710 59106
rect 57762 59054 57774 59106
rect 49646 59042 49698 59054
rect 55582 59042 55634 59054
rect 37214 58994 37266 59006
rect 35746 58942 35758 58994
rect 35810 58942 35822 58994
rect 37214 58930 37266 58942
rect 44942 58994 44994 59006
rect 44942 58930 44994 58942
rect 45278 58994 45330 59006
rect 55570 58942 55582 58994
rect 55634 58991 55646 58994
rect 56130 58991 56142 58994
rect 55634 58945 56142 58991
rect 55634 58942 55646 58945
rect 56130 58942 56142 58945
rect 56194 58942 56206 58994
rect 45278 58930 45330 58942
rect 1344 58826 58576 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 58576 58826
rect 1344 58740 58576 58774
rect 16382 58658 16434 58670
rect 16382 58594 16434 58606
rect 16718 58658 16770 58670
rect 35982 58658 36034 58670
rect 25778 58606 25790 58658
rect 25842 58655 25854 58658
rect 26114 58655 26126 58658
rect 25842 58609 26126 58655
rect 25842 58606 25854 58609
rect 26114 58606 26126 58609
rect 26178 58606 26190 58658
rect 16718 58594 16770 58606
rect 35982 58594 36034 58606
rect 43150 58658 43202 58670
rect 43150 58594 43202 58606
rect 52110 58658 52162 58670
rect 52110 58594 52162 58606
rect 4846 58546 4898 58558
rect 12350 58546 12402 58558
rect 10210 58494 10222 58546
rect 10274 58494 10286 58546
rect 4846 58482 4898 58494
rect 12350 58482 12402 58494
rect 14478 58546 14530 58558
rect 41806 58546 41858 58558
rect 48190 58546 48242 58558
rect 27346 58494 27358 58546
rect 27410 58494 27422 58546
rect 39218 58494 39230 58546
rect 39282 58494 39294 58546
rect 41346 58494 41358 58546
rect 41410 58494 41422 58546
rect 44818 58494 44830 58546
rect 44882 58494 44894 58546
rect 46946 58494 46958 58546
rect 47010 58494 47022 58546
rect 14478 58482 14530 58494
rect 41806 58482 41858 58494
rect 48190 58482 48242 58494
rect 51998 58546 52050 58558
rect 58270 58546 58322 58558
rect 54674 58494 54686 58546
rect 54738 58494 54750 58546
rect 51998 58482 52050 58494
rect 58270 58482 58322 58494
rect 2270 58434 2322 58446
rect 2270 58370 2322 58382
rect 4174 58434 4226 58446
rect 4174 58370 4226 58382
rect 4286 58434 4338 58446
rect 4286 58370 4338 58382
rect 5630 58434 5682 58446
rect 25678 58434 25730 58446
rect 43262 58434 43314 58446
rect 11778 58382 11790 58434
rect 11842 58382 11854 58434
rect 26674 58382 26686 58434
rect 26738 58382 26750 58434
rect 27794 58382 27806 58434
rect 27858 58382 27870 58434
rect 38546 58382 38558 58434
rect 38610 58382 38622 58434
rect 47730 58382 47742 58434
rect 47794 58382 47806 58434
rect 52994 58382 53006 58434
rect 53058 58382 53070 58434
rect 5630 58370 5682 58382
rect 25678 58370 25730 58382
rect 43262 58370 43314 58382
rect 1710 58322 1762 58334
rect 1710 58258 1762 58270
rect 3838 58322 3890 58334
rect 15822 58322 15874 58334
rect 10658 58270 10670 58322
rect 10722 58270 10734 58322
rect 13458 58270 13470 58322
rect 13522 58270 13534 58322
rect 3838 58258 3890 58270
rect 15822 58258 15874 58270
rect 16158 58322 16210 58334
rect 16158 58258 16210 58270
rect 25342 58322 25394 58334
rect 29822 58322 29874 58334
rect 28130 58270 28142 58322
rect 28194 58270 28206 58322
rect 25342 58258 25394 58270
rect 29822 58258 29874 58270
rect 30494 58322 30546 58334
rect 30494 58258 30546 58270
rect 36318 58322 36370 58334
rect 36318 58258 36370 58270
rect 43150 58322 43202 58334
rect 43150 58258 43202 58270
rect 3950 58210 4002 58222
rect 3950 58146 4002 58158
rect 5742 58210 5794 58222
rect 5742 58146 5794 58158
rect 5966 58210 6018 58222
rect 5966 58146 6018 58158
rect 13806 58210 13858 58222
rect 13806 58146 13858 58158
rect 15374 58210 15426 58222
rect 15374 58146 15426 58158
rect 25454 58210 25506 58222
rect 25454 58146 25506 58158
rect 26126 58210 26178 58222
rect 26126 58146 26178 58158
rect 29934 58210 29986 58222
rect 29934 58146 29986 58158
rect 30046 58210 30098 58222
rect 30046 58146 30098 58158
rect 30606 58210 30658 58222
rect 30606 58146 30658 58158
rect 30830 58210 30882 58222
rect 30830 58146 30882 58158
rect 36094 58210 36146 58222
rect 36094 58146 36146 58158
rect 1344 58042 58576 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 58576 58042
rect 1344 57956 58576 57990
rect 9886 57874 9938 57886
rect 6850 57822 6862 57874
rect 6914 57822 6926 57874
rect 9886 57810 9938 57822
rect 10558 57874 10610 57886
rect 10558 57810 10610 57822
rect 20526 57874 20578 57886
rect 28030 57874 28082 57886
rect 51662 57874 51714 57886
rect 25330 57822 25342 57874
rect 25394 57822 25406 57874
rect 44930 57822 44942 57874
rect 44994 57822 45006 57874
rect 20526 57810 20578 57822
rect 28030 57810 28082 57822
rect 51662 57810 51714 57822
rect 52558 57874 52610 57886
rect 52558 57810 52610 57822
rect 4958 57762 5010 57774
rect 2482 57710 2494 57762
rect 2546 57710 2558 57762
rect 4958 57698 5010 57710
rect 13806 57762 13858 57774
rect 13806 57698 13858 57710
rect 19630 57762 19682 57774
rect 19630 57698 19682 57710
rect 19742 57762 19794 57774
rect 19742 57698 19794 57710
rect 22878 57762 22930 57774
rect 23986 57710 23998 57762
rect 24050 57710 24062 57762
rect 27682 57710 27694 57762
rect 27746 57710 27758 57762
rect 30034 57710 30046 57762
rect 30098 57710 30110 57762
rect 36418 57710 36430 57762
rect 36482 57710 36494 57762
rect 38994 57710 39006 57762
rect 39058 57710 39070 57762
rect 43250 57710 43262 57762
rect 43314 57710 43326 57762
rect 22878 57698 22930 57710
rect 6302 57650 6354 57662
rect 1810 57598 1822 57650
rect 1874 57598 1886 57650
rect 5618 57598 5630 57650
rect 5682 57598 5694 57650
rect 6302 57586 6354 57598
rect 7982 57650 8034 57662
rect 7982 57586 8034 57598
rect 8318 57650 8370 57662
rect 8318 57586 8370 57598
rect 8542 57650 8594 57662
rect 8542 57586 8594 57598
rect 9438 57650 9490 57662
rect 9438 57586 9490 57598
rect 10110 57650 10162 57662
rect 10110 57586 10162 57598
rect 10334 57650 10386 57662
rect 10334 57586 10386 57598
rect 10670 57650 10722 57662
rect 10670 57586 10722 57598
rect 13918 57650 13970 57662
rect 13918 57586 13970 57598
rect 19406 57650 19458 57662
rect 19406 57586 19458 57598
rect 20078 57650 20130 57662
rect 20078 57586 20130 57598
rect 20302 57650 20354 57662
rect 20302 57586 20354 57598
rect 20750 57650 20802 57662
rect 20750 57586 20802 57598
rect 22766 57650 22818 57662
rect 25678 57650 25730 57662
rect 51438 57650 51490 57662
rect 23650 57598 23662 57650
rect 23714 57598 23726 57650
rect 24658 57598 24670 57650
rect 24722 57598 24734 57650
rect 26450 57598 26462 57650
rect 26514 57598 26526 57650
rect 27010 57598 27022 57650
rect 27074 57598 27086 57650
rect 28242 57598 28254 57650
rect 28306 57598 28318 57650
rect 30258 57598 30270 57650
rect 30322 57598 30334 57650
rect 30930 57598 30942 57650
rect 30994 57598 31006 57650
rect 32386 57598 32398 57650
rect 32450 57598 32462 57650
rect 37650 57598 37662 57650
rect 37714 57598 37726 57650
rect 42130 57598 42142 57650
rect 42194 57598 42206 57650
rect 44482 57598 44494 57650
rect 44546 57598 44558 57650
rect 51986 57598 51998 57650
rect 52050 57598 52062 57650
rect 22766 57586 22818 57598
rect 25678 57586 25730 57598
rect 51438 57586 51490 57598
rect 8094 57538 8146 57550
rect 4610 57486 4622 57538
rect 4674 57486 4686 57538
rect 5842 57486 5854 57538
rect 5906 57486 5918 57538
rect 8094 57474 8146 57486
rect 9998 57538 10050 57550
rect 9998 57474 10050 57486
rect 13358 57538 13410 57550
rect 31614 57538 31666 57550
rect 23762 57486 23774 57538
rect 23826 57486 23838 57538
rect 13358 57474 13410 57486
rect 31614 57474 31666 57486
rect 32062 57538 32114 57550
rect 32062 57474 32114 57486
rect 33182 57538 33234 57550
rect 42590 57538 42642 57550
rect 36194 57486 36206 57538
rect 36258 57486 36270 57538
rect 33182 57474 33234 57486
rect 42590 57474 42642 57486
rect 43150 57538 43202 57550
rect 43150 57474 43202 57486
rect 51102 57538 51154 57550
rect 51102 57474 51154 57486
rect 51550 57538 51602 57550
rect 51550 57474 51602 57486
rect 6526 57426 6578 57438
rect 6526 57362 6578 57374
rect 13806 57426 13858 57438
rect 13806 57362 13858 57374
rect 22654 57426 22706 57438
rect 22654 57362 22706 57374
rect 32398 57426 32450 57438
rect 32398 57362 32450 57374
rect 1344 57258 58576 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 58576 57258
rect 1344 57172 58576 57206
rect 12238 57090 12290 57102
rect 12238 57026 12290 57038
rect 24670 57090 24722 57102
rect 24670 57026 24722 57038
rect 27246 57090 27298 57102
rect 43598 57090 43650 57102
rect 29810 57038 29822 57090
rect 29874 57038 29886 57090
rect 27246 57026 27298 57038
rect 43598 57026 43650 57038
rect 4510 56978 4562 56990
rect 4510 56914 4562 56926
rect 6078 56978 6130 56990
rect 14142 56978 14194 56990
rect 7410 56926 7422 56978
rect 7474 56926 7486 56978
rect 9538 56926 9550 56978
rect 9602 56926 9614 56978
rect 10658 56926 10670 56978
rect 10722 56926 10734 56978
rect 6078 56914 6130 56926
rect 14142 56914 14194 56926
rect 15038 56978 15090 56990
rect 15038 56914 15090 56926
rect 16158 56978 16210 56990
rect 20190 56978 20242 56990
rect 34974 56978 35026 56990
rect 19394 56926 19406 56978
rect 19458 56926 19470 56978
rect 22082 56926 22094 56978
rect 22146 56926 22158 56978
rect 24210 56926 24222 56978
rect 24274 56926 24286 56978
rect 29922 56926 29934 56978
rect 29986 56926 29998 56978
rect 31602 56926 31614 56978
rect 31666 56926 31678 56978
rect 33730 56926 33742 56978
rect 33794 56926 33806 56978
rect 16158 56914 16210 56926
rect 20190 56914 20242 56926
rect 34974 56914 35026 56926
rect 36318 56978 36370 56990
rect 36318 56914 36370 56926
rect 42366 56978 42418 56990
rect 42366 56914 42418 56926
rect 42702 56978 42754 56990
rect 50430 56978 50482 56990
rect 47058 56926 47070 56978
rect 47122 56926 47134 56978
rect 55346 56926 55358 56978
rect 55410 56926 55422 56978
rect 42702 56914 42754 56926
rect 50430 56914 50482 56926
rect 4622 56866 4674 56878
rect 4622 56802 4674 56814
rect 5070 56866 5122 56878
rect 5070 56802 5122 56814
rect 5518 56866 5570 56878
rect 5518 56802 5570 56814
rect 5966 56866 6018 56878
rect 20302 56866 20354 56878
rect 6738 56814 6750 56866
rect 6802 56814 6814 56866
rect 10546 56814 10558 56866
rect 10610 56814 10622 56866
rect 16482 56814 16494 56866
rect 16546 56814 16558 56866
rect 5966 56802 6018 56814
rect 20302 56802 20354 56814
rect 20750 56866 20802 56878
rect 25454 56866 25506 56878
rect 26686 56866 26738 56878
rect 35982 56866 36034 56878
rect 21298 56814 21310 56866
rect 21362 56814 21374 56866
rect 26114 56814 26126 56866
rect 26178 56814 26190 56866
rect 30146 56814 30158 56866
rect 30210 56814 30222 56866
rect 30818 56814 30830 56866
rect 30882 56814 30894 56866
rect 34514 56814 34526 56866
rect 34578 56814 34590 56866
rect 20750 56802 20802 56814
rect 25454 56802 25506 56814
rect 26686 56802 26738 56814
rect 35982 56802 36034 56814
rect 37102 56866 37154 56878
rect 37998 56866 38050 56878
rect 37314 56814 37326 56866
rect 37378 56814 37390 56866
rect 37102 56802 37154 56814
rect 37998 56802 38050 56814
rect 42254 56866 42306 56878
rect 42254 56802 42306 56814
rect 42926 56866 42978 56878
rect 49970 56814 49982 56866
rect 50034 56814 50046 56866
rect 42926 56802 42978 56814
rect 4398 56754 4450 56766
rect 4398 56690 4450 56702
rect 9886 56754 9938 56766
rect 9886 56690 9938 56702
rect 12014 56754 12066 56766
rect 13918 56754 13970 56766
rect 13794 56702 13806 56754
rect 13858 56702 13870 56754
rect 12014 56690 12066 56702
rect 13918 56690 13970 56702
rect 14254 56754 14306 56766
rect 14254 56690 14306 56702
rect 15150 56754 15202 56766
rect 19854 56754 19906 56766
rect 17266 56702 17278 56754
rect 17330 56702 17342 56754
rect 15150 56690 15202 56702
rect 19854 56690 19906 56702
rect 24782 56754 24834 56766
rect 26798 56754 26850 56766
rect 25106 56702 25118 56754
rect 25170 56702 25182 56754
rect 24782 56690 24834 56702
rect 26798 56690 26850 56702
rect 27134 56754 27186 56766
rect 27134 56690 27186 56702
rect 36094 56754 36146 56766
rect 36094 56690 36146 56702
rect 36430 56754 36482 56766
rect 36430 56690 36482 56702
rect 42478 56754 42530 56766
rect 42478 56690 42530 56702
rect 43262 56754 43314 56766
rect 43262 56690 43314 56702
rect 43486 56754 43538 56766
rect 55582 56754 55634 56766
rect 49186 56702 49198 56754
rect 49250 56702 49262 56754
rect 43486 56690 43538 56702
rect 55582 56690 55634 56702
rect 6190 56642 6242 56654
rect 14030 56642 14082 56654
rect 12562 56590 12574 56642
rect 12626 56590 12638 56642
rect 6190 56578 6242 56590
rect 14030 56578 14082 56590
rect 14702 56642 14754 56654
rect 14702 56578 14754 56590
rect 14926 56642 14978 56654
rect 14926 56578 14978 56590
rect 20078 56642 20130 56654
rect 20078 56578 20130 56590
rect 24670 56642 24722 56654
rect 24670 56578 24722 56590
rect 27694 56642 27746 56654
rect 27694 56578 27746 56590
rect 55358 56642 55410 56654
rect 55358 56578 55410 56590
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 8654 56306 8706 56318
rect 8654 56242 8706 56254
rect 8766 56306 8818 56318
rect 8766 56242 8818 56254
rect 9774 56306 9826 56318
rect 13694 56306 13746 56318
rect 28478 56306 28530 56318
rect 46958 56306 47010 56318
rect 10770 56254 10782 56306
rect 10834 56254 10846 56306
rect 11218 56254 11230 56306
rect 11282 56254 11294 56306
rect 12114 56254 12126 56306
rect 12178 56254 12190 56306
rect 22642 56254 22654 56306
rect 22706 56254 22718 56306
rect 36530 56254 36542 56306
rect 36594 56254 36606 56306
rect 9774 56242 9826 56254
rect 13694 56242 13746 56254
rect 28478 56242 28530 56254
rect 46958 56242 47010 56254
rect 48190 56306 48242 56318
rect 48190 56242 48242 56254
rect 48862 56306 48914 56318
rect 54238 56306 54290 56318
rect 49970 56254 49982 56306
rect 50034 56254 50046 56306
rect 48862 56242 48914 56254
rect 54238 56242 54290 56254
rect 8318 56194 8370 56206
rect 8318 56130 8370 56142
rect 12910 56194 12962 56206
rect 12910 56130 12962 56142
rect 13134 56194 13186 56206
rect 13134 56130 13186 56142
rect 13358 56194 13410 56206
rect 13358 56130 13410 56142
rect 13470 56194 13522 56206
rect 13470 56130 13522 56142
rect 13918 56194 13970 56206
rect 13918 56130 13970 56142
rect 14030 56194 14082 56206
rect 14030 56130 14082 56142
rect 16046 56194 16098 56206
rect 16046 56130 16098 56142
rect 17950 56194 18002 56206
rect 48750 56194 48802 56206
rect 19058 56142 19070 56194
rect 19122 56142 19134 56194
rect 20290 56142 20302 56194
rect 20354 56142 20366 56194
rect 23874 56142 23886 56194
rect 23938 56142 23950 56194
rect 31826 56142 31838 56194
rect 31890 56142 31902 56194
rect 32498 56142 32510 56194
rect 32562 56142 32574 56194
rect 35186 56142 35198 56194
rect 35250 56142 35262 56194
rect 35634 56142 35646 56194
rect 35698 56142 35710 56194
rect 51650 56142 51662 56194
rect 51714 56142 51726 56194
rect 17950 56130 18002 56142
rect 48750 56130 48802 56142
rect 8542 56082 8594 56094
rect 8542 56018 8594 56030
rect 10222 56082 10274 56094
rect 10222 56018 10274 56030
rect 10446 56082 10498 56094
rect 10446 56018 10498 56030
rect 11566 56082 11618 56094
rect 11566 56018 11618 56030
rect 12462 56082 12514 56094
rect 12462 56018 12514 56030
rect 12798 56082 12850 56094
rect 12798 56018 12850 56030
rect 14254 56082 14306 56094
rect 14254 56018 14306 56030
rect 14590 56082 14642 56094
rect 38222 56082 38274 56094
rect 47070 56082 47122 56094
rect 15138 56030 15150 56082
rect 15202 56030 15214 56082
rect 22978 56030 22990 56082
rect 23042 56030 23054 56082
rect 32274 56030 32286 56082
rect 32338 56030 32350 56082
rect 33618 56030 33630 56082
rect 33682 56030 33694 56082
rect 34178 56030 34190 56082
rect 34242 56030 34254 56082
rect 35522 56030 35534 56082
rect 35586 56030 35598 56082
rect 37202 56030 37214 56082
rect 37266 56030 37278 56082
rect 38994 56030 39006 56082
rect 39058 56030 39070 56082
rect 14590 56018 14642 56030
rect 38222 56018 38274 56030
rect 47070 56018 47122 56030
rect 47182 56082 47234 56094
rect 48078 56082 48130 56094
rect 47618 56030 47630 56082
rect 47682 56030 47694 56082
rect 47182 56018 47234 56030
rect 48078 56018 48130 56030
rect 50318 56082 50370 56094
rect 50866 56030 50878 56082
rect 50930 56030 50942 56082
rect 54898 56030 54910 56082
rect 54962 56030 54974 56082
rect 50318 56018 50370 56030
rect 4622 55970 4674 55982
rect 4622 55906 4674 55918
rect 5182 55970 5234 55982
rect 18174 55970 18226 55982
rect 15250 55918 15262 55970
rect 15314 55918 15326 55970
rect 17826 55918 17838 55970
rect 17890 55918 17902 55970
rect 5182 55906 5234 55918
rect 18174 55906 18226 55918
rect 18734 55970 18786 55982
rect 18734 55906 18786 55918
rect 20750 55970 20802 55982
rect 25342 55970 25394 55982
rect 24434 55918 24446 55970
rect 24498 55918 24510 55970
rect 20750 55906 20802 55918
rect 25342 55906 25394 55918
rect 31390 55970 31442 55982
rect 31390 55906 31442 55918
rect 45502 55970 45554 55982
rect 45502 55906 45554 55918
rect 47854 55970 47906 55982
rect 53778 55918 53790 55970
rect 53842 55918 53854 55970
rect 55122 55918 55134 55970
rect 55186 55918 55198 55970
rect 47854 55906 47906 55918
rect 45614 55858 45666 55870
rect 30930 55806 30942 55858
rect 30994 55855 31006 55858
rect 31378 55855 31390 55858
rect 30994 55809 31390 55855
rect 30994 55806 31006 55809
rect 31378 55806 31390 55809
rect 31442 55806 31454 55858
rect 55570 55806 55582 55858
rect 55634 55806 55646 55858
rect 45614 55794 45666 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 4846 55522 4898 55534
rect 4846 55458 4898 55470
rect 32286 55522 32338 55534
rect 43150 55522 43202 55534
rect 35186 55470 35198 55522
rect 35250 55470 35262 55522
rect 32286 55458 32338 55470
rect 43150 55458 43202 55470
rect 11790 55410 11842 55422
rect 11790 55346 11842 55358
rect 23550 55410 23602 55422
rect 23762 55358 23774 55410
rect 23826 55358 23838 55410
rect 33058 55358 33070 55410
rect 33122 55358 33134 55410
rect 34850 55358 34862 55410
rect 34914 55358 34926 55410
rect 40450 55358 40462 55410
rect 40514 55358 40526 55410
rect 41570 55358 41582 55410
rect 41634 55358 41646 55410
rect 42130 55358 42142 55410
rect 42194 55358 42206 55410
rect 45602 55358 45614 55410
rect 45666 55358 45678 55410
rect 47730 55358 47742 55410
rect 47794 55358 47806 55410
rect 52770 55358 52782 55410
rect 52834 55358 52846 55410
rect 55570 55358 55582 55410
rect 55634 55358 55646 55410
rect 57698 55358 57710 55410
rect 57762 55358 57774 55410
rect 23550 55346 23602 55358
rect 2942 55298 2994 55310
rect 2942 55234 2994 55246
rect 3502 55298 3554 55310
rect 3502 55234 3554 55246
rect 3950 55298 4002 55310
rect 3950 55234 4002 55246
rect 4510 55298 4562 55310
rect 4510 55234 4562 55246
rect 11006 55298 11058 55310
rect 11006 55234 11058 55246
rect 11342 55298 11394 55310
rect 11342 55234 11394 55246
rect 14478 55298 14530 55310
rect 28366 55298 28418 55310
rect 31726 55298 31778 55310
rect 33854 55298 33906 55310
rect 42814 55298 42866 55310
rect 58158 55298 58210 55310
rect 23874 55246 23886 55298
rect 23938 55246 23950 55298
rect 29250 55246 29262 55298
rect 29314 55246 29326 55298
rect 30146 55246 30158 55298
rect 30210 55246 30222 55298
rect 30930 55246 30942 55298
rect 30994 55246 31006 55298
rect 32946 55246 32958 55298
rect 33010 55246 33022 55298
rect 34738 55246 34750 55298
rect 34802 55246 34814 55298
rect 37650 55246 37662 55298
rect 37714 55246 37726 55298
rect 41458 55246 41470 55298
rect 41522 55246 41534 55298
rect 42354 55246 42366 55298
rect 42418 55246 42430 55298
rect 44930 55246 44942 55298
rect 44994 55246 45006 55298
rect 53330 55246 53342 55298
rect 53394 55246 53406 55298
rect 54898 55246 54910 55298
rect 54962 55246 54974 55298
rect 14478 55234 14530 55246
rect 28366 55234 28418 55246
rect 31726 55234 31778 55246
rect 33854 55234 33906 55246
rect 42814 55234 42866 55246
rect 58158 55234 58210 55246
rect 3278 55186 3330 55198
rect 3278 55122 3330 55134
rect 4958 55186 5010 55198
rect 31390 55186 31442 55198
rect 29362 55134 29374 55186
rect 29426 55134 29438 55186
rect 30706 55134 30718 55186
rect 30770 55134 30782 55186
rect 4958 55122 5010 55134
rect 31390 55122 31442 55134
rect 32286 55186 32338 55198
rect 32286 55122 32338 55134
rect 32398 55186 32450 55198
rect 40798 55186 40850 55198
rect 38322 55134 38334 55186
rect 38386 55134 38398 55186
rect 49970 55134 49982 55186
rect 50034 55134 50046 55186
rect 32398 55122 32450 55134
rect 40798 55122 40850 55134
rect 3054 55074 3106 55086
rect 3054 55010 3106 55022
rect 3838 55074 3890 55086
rect 3838 55010 3890 55022
rect 4062 55074 4114 55086
rect 4062 55010 4114 55022
rect 4846 55074 4898 55086
rect 4846 55010 4898 55022
rect 11118 55074 11170 55086
rect 11118 55010 11170 55022
rect 12686 55074 12738 55086
rect 12686 55010 12738 55022
rect 13582 55074 13634 55086
rect 13582 55010 13634 55022
rect 14590 55074 14642 55086
rect 14590 55010 14642 55022
rect 18398 55074 18450 55086
rect 18398 55010 18450 55022
rect 27694 55074 27746 55086
rect 27694 55010 27746 55022
rect 27806 55074 27858 55086
rect 27806 55010 27858 55022
rect 27918 55074 27970 55086
rect 31502 55074 31554 55086
rect 30146 55022 30158 55074
rect 30210 55022 30222 55074
rect 27918 55010 27970 55022
rect 31502 55010 31554 55022
rect 43038 55074 43090 55086
rect 43038 55010 43090 55022
rect 44270 55074 44322 55086
rect 49534 55074 49586 55086
rect 49186 55022 49198 55074
rect 49250 55022 49262 55074
rect 44270 55010 44322 55022
rect 49534 55010 49586 55022
rect 50318 55074 50370 55086
rect 50318 55010 50370 55022
rect 52782 55074 52834 55086
rect 52782 55010 52834 55022
rect 52894 55074 52946 55086
rect 52894 55010 52946 55022
rect 53118 55074 53170 55086
rect 53118 55010 53170 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 5070 54738 5122 54750
rect 39566 54738 39618 54750
rect 10994 54686 11006 54738
rect 11058 54686 11070 54738
rect 29474 54686 29486 54738
rect 29538 54686 29550 54738
rect 5070 54674 5122 54686
rect 39566 54674 39618 54686
rect 41022 54738 41074 54750
rect 41022 54674 41074 54686
rect 41582 54738 41634 54750
rect 41582 54674 41634 54686
rect 41694 54738 41746 54750
rect 41694 54674 41746 54686
rect 41806 54738 41858 54750
rect 41806 54674 41858 54686
rect 42478 54738 42530 54750
rect 42478 54674 42530 54686
rect 45502 54738 45554 54750
rect 45502 54674 45554 54686
rect 45950 54738 46002 54750
rect 45950 54674 46002 54686
rect 46622 54738 46674 54750
rect 51874 54686 51886 54738
rect 51938 54686 51950 54738
rect 46622 54674 46674 54686
rect 5406 54626 5458 54638
rect 2482 54574 2494 54626
rect 2546 54574 2558 54626
rect 5406 54562 5458 54574
rect 14590 54626 14642 54638
rect 14590 54562 14642 54574
rect 26686 54626 26738 54638
rect 26686 54562 26738 54574
rect 27022 54626 27074 54638
rect 27022 54562 27074 54574
rect 31502 54626 31554 54638
rect 31502 54562 31554 54574
rect 31950 54626 32002 54638
rect 31950 54562 32002 54574
rect 39454 54626 39506 54638
rect 39454 54562 39506 54574
rect 42366 54626 42418 54638
rect 55806 54626 55858 54638
rect 51202 54574 51214 54626
rect 51266 54574 51278 54626
rect 42366 54562 42418 54574
rect 55806 54562 55858 54574
rect 4958 54514 5010 54526
rect 1810 54462 1822 54514
rect 1874 54462 1886 54514
rect 4958 54450 5010 54462
rect 5182 54514 5234 54526
rect 5182 54450 5234 54462
rect 11342 54514 11394 54526
rect 11342 54450 11394 54462
rect 14254 54514 14306 54526
rect 14254 54450 14306 54462
rect 14478 54514 14530 54526
rect 14478 54450 14530 54462
rect 14814 54514 14866 54526
rect 18286 54514 18338 54526
rect 15138 54462 15150 54514
rect 15202 54462 15214 54514
rect 15474 54462 15486 54514
rect 15538 54462 15550 54514
rect 14814 54450 14866 54462
rect 18286 54450 18338 54462
rect 27246 54514 27298 54526
rect 27246 54450 27298 54462
rect 27582 54514 27634 54526
rect 39790 54514 39842 54526
rect 28130 54462 28142 54514
rect 28194 54462 28206 54514
rect 30818 54462 30830 54514
rect 30882 54462 30894 54514
rect 27582 54450 27634 54462
rect 39790 54450 39842 54462
rect 40014 54514 40066 54526
rect 40014 54450 40066 54462
rect 41470 54514 41522 54526
rect 46062 54514 46114 54526
rect 42018 54462 42030 54514
rect 42082 54462 42094 54514
rect 41470 54450 41522 54462
rect 46062 54450 46114 54462
rect 46398 54514 46450 54526
rect 50878 54514 50930 54526
rect 56478 54514 56530 54526
rect 46610 54462 46622 54514
rect 46674 54462 46686 54514
rect 51650 54462 51662 54514
rect 51714 54462 51726 54514
rect 46398 54450 46450 54462
rect 50878 54450 50930 54462
rect 56478 54450 56530 54462
rect 56814 54514 56866 54526
rect 56814 54450 56866 54462
rect 57150 54514 57202 54526
rect 57150 54450 57202 54462
rect 26798 54402 26850 54414
rect 28926 54402 28978 54414
rect 4610 54350 4622 54402
rect 4674 54350 4686 54402
rect 16706 54350 16718 54402
rect 16770 54350 16782 54402
rect 28466 54350 28478 54402
rect 28530 54350 28542 54402
rect 26798 54338 26850 54350
rect 28926 54338 28978 54350
rect 29150 54402 29202 54414
rect 46846 54402 46898 54414
rect 30594 54350 30606 54402
rect 30658 54350 30670 54402
rect 29150 54338 29202 54350
rect 46846 54338 46898 54350
rect 47182 54402 47234 54414
rect 47182 54338 47234 54350
rect 55134 54402 55186 54414
rect 55134 54338 55186 54350
rect 55918 54402 55970 54414
rect 55918 54338 55970 54350
rect 56702 54402 56754 54414
rect 56702 54338 56754 54350
rect 54910 54290 54962 54302
rect 54562 54238 54574 54290
rect 54626 54238 54638 54290
rect 54910 54226 54962 54238
rect 56030 54290 56082 54302
rect 56030 54226 56082 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 8990 53954 9042 53966
rect 8990 53890 9042 53902
rect 23326 53954 23378 53966
rect 23326 53890 23378 53902
rect 29374 53954 29426 53966
rect 29374 53890 29426 53902
rect 29710 53954 29762 53966
rect 52670 53954 52722 53966
rect 36306 53902 36318 53954
rect 36370 53902 36382 53954
rect 29710 53890 29762 53902
rect 52670 53890 52722 53902
rect 2942 53842 2994 53854
rect 2942 53778 2994 53790
rect 18734 53842 18786 53854
rect 29150 53842 29202 53854
rect 40014 53842 40066 53854
rect 22306 53790 22318 53842
rect 22370 53790 22382 53842
rect 24098 53790 24110 53842
rect 24162 53790 24174 53842
rect 26002 53790 26014 53842
rect 26066 53790 26078 53842
rect 28130 53790 28142 53842
rect 28194 53790 28206 53842
rect 36082 53790 36094 53842
rect 36146 53790 36158 53842
rect 37090 53790 37102 53842
rect 37154 53790 37166 53842
rect 18734 53778 18786 53790
rect 29150 53778 29202 53790
rect 40014 53778 40066 53790
rect 53006 53842 53058 53854
rect 53006 53778 53058 53790
rect 53902 53842 53954 53854
rect 56018 53790 56030 53842
rect 56082 53790 56094 53842
rect 58146 53790 58158 53842
rect 58210 53790 58222 53842
rect 53902 53778 53954 53790
rect 3838 53730 3890 53742
rect 3378 53678 3390 53730
rect 3442 53678 3454 53730
rect 3838 53666 3890 53678
rect 4622 53730 4674 53742
rect 4622 53666 4674 53678
rect 5070 53730 5122 53742
rect 5070 53666 5122 53678
rect 7870 53730 7922 53742
rect 7870 53666 7922 53678
rect 8430 53730 8482 53742
rect 8430 53666 8482 53678
rect 8878 53730 8930 53742
rect 8878 53666 8930 53678
rect 17838 53730 17890 53742
rect 17838 53666 17890 53678
rect 18398 53730 18450 53742
rect 18398 53666 18450 53678
rect 19854 53730 19906 53742
rect 19854 53666 19906 53678
rect 19966 53730 20018 53742
rect 37998 53730 38050 53742
rect 23874 53678 23886 53730
rect 23938 53678 23950 53730
rect 24770 53678 24782 53730
rect 24834 53678 24846 53730
rect 25218 53678 25230 53730
rect 25282 53678 25294 53730
rect 34514 53678 34526 53730
rect 34578 53678 34590 53730
rect 35970 53678 35982 53730
rect 36034 53678 36046 53730
rect 37314 53678 37326 53730
rect 37378 53678 37390 53730
rect 19966 53666 20018 53678
rect 37998 53666 38050 53678
rect 39902 53730 39954 53742
rect 39902 53666 39954 53678
rect 40574 53730 40626 53742
rect 51426 53678 51438 53730
rect 51490 53678 51502 53730
rect 54898 53678 54910 53730
rect 54962 53678 54974 53730
rect 55234 53678 55246 53730
rect 55298 53678 55310 53730
rect 40574 53666 40626 53678
rect 4286 53618 4338 53630
rect 4286 53554 4338 53566
rect 4398 53618 4450 53630
rect 4398 53554 4450 53566
rect 7086 53618 7138 53630
rect 7086 53554 7138 53566
rect 7422 53618 7474 53630
rect 7422 53554 7474 53566
rect 7646 53618 7698 53630
rect 17950 53618 18002 53630
rect 10322 53566 10334 53618
rect 10386 53566 10398 53618
rect 7646 53554 7698 53566
rect 17950 53554 18002 53566
rect 19070 53618 19122 53630
rect 19070 53554 19122 53566
rect 20638 53618 20690 53630
rect 20638 53554 20690 53566
rect 22654 53618 22706 53630
rect 22654 53554 22706 53566
rect 23102 53618 23154 53630
rect 39566 53618 39618 53630
rect 24322 53566 24334 53618
rect 24386 53566 24398 53618
rect 30370 53566 30382 53618
rect 30434 53566 30446 53618
rect 23102 53554 23154 53566
rect 39566 53554 39618 53566
rect 40910 53618 40962 53630
rect 40910 53554 40962 53566
rect 41246 53618 41298 53630
rect 41246 53554 41298 53566
rect 41582 53618 41634 53630
rect 41582 53554 41634 53566
rect 41694 53618 41746 53630
rect 54226 53566 54238 53618
rect 54290 53566 54302 53618
rect 54786 53566 54798 53618
rect 54850 53566 54862 53618
rect 41694 53554 41746 53566
rect 7198 53506 7250 53518
rect 7198 53442 7250 53454
rect 8318 53506 8370 53518
rect 8318 53442 8370 53454
rect 8542 53506 8594 53518
rect 8542 53442 8594 53454
rect 8990 53506 9042 53518
rect 8990 53442 9042 53454
rect 10670 53506 10722 53518
rect 10670 53442 10722 53454
rect 18174 53506 18226 53518
rect 18174 53442 18226 53454
rect 18622 53506 18674 53518
rect 18622 53442 18674 53454
rect 18846 53506 18898 53518
rect 18846 53442 18898 53454
rect 19630 53506 19682 53518
rect 19630 53442 19682 53454
rect 20078 53506 20130 53518
rect 20078 53442 20130 53454
rect 20302 53506 20354 53518
rect 20302 53442 20354 53454
rect 20526 53506 20578 53518
rect 20526 53442 20578 53454
rect 22430 53506 22482 53518
rect 22430 53442 22482 53454
rect 23214 53506 23266 53518
rect 23214 53442 23266 53454
rect 30046 53506 30098 53518
rect 30046 53442 30098 53454
rect 33182 53506 33234 53518
rect 33182 53442 33234 53454
rect 40126 53506 40178 53518
rect 40126 53442 40178 53454
rect 41022 53506 41074 53518
rect 41022 53442 41074 53454
rect 41358 53506 41410 53518
rect 52782 53506 52834 53518
rect 51650 53454 51662 53506
rect 51714 53454 51726 53506
rect 41358 53442 41410 53454
rect 52782 53442 52834 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 14590 53170 14642 53182
rect 14590 53106 14642 53118
rect 23998 53170 24050 53182
rect 23998 53106 24050 53118
rect 24670 53170 24722 53182
rect 24670 53106 24722 53118
rect 25342 53170 25394 53182
rect 25342 53106 25394 53118
rect 31278 53170 31330 53182
rect 31278 53106 31330 53118
rect 36430 53170 36482 53182
rect 36430 53106 36482 53118
rect 45838 53170 45890 53182
rect 45838 53106 45890 53118
rect 46622 53170 46674 53182
rect 46622 53106 46674 53118
rect 46846 53170 46898 53182
rect 46846 53106 46898 53118
rect 47518 53170 47570 53182
rect 47518 53106 47570 53118
rect 47966 53170 48018 53182
rect 47966 53106 48018 53118
rect 55022 53170 55074 53182
rect 55022 53106 55074 53118
rect 8542 53058 8594 53070
rect 5954 53006 5966 53058
rect 6018 53006 6030 53058
rect 8542 52994 8594 53006
rect 12014 53058 12066 53070
rect 12014 52994 12066 53006
rect 12574 53058 12626 53070
rect 12574 52994 12626 53006
rect 14814 53058 14866 53070
rect 23886 53058 23938 53070
rect 18162 53006 18174 53058
rect 18226 53006 18238 53058
rect 21410 53006 21422 53058
rect 21474 53006 21486 53058
rect 14814 52994 14866 53006
rect 23886 52994 23938 53006
rect 36206 53058 36258 53070
rect 36206 52994 36258 53006
rect 36654 53058 36706 53070
rect 51538 53006 51550 53058
rect 51602 53006 51614 53058
rect 36654 52994 36706 53006
rect 8430 52946 8482 52958
rect 5170 52894 5182 52946
rect 5234 52894 5246 52946
rect 8430 52882 8482 52894
rect 8654 52946 8706 52958
rect 10334 52946 10386 52958
rect 12686 52946 12738 52958
rect 8978 52894 8990 52946
rect 9042 52894 9054 52946
rect 11554 52894 11566 52946
rect 11618 52894 11630 52946
rect 12338 52894 12350 52946
rect 12402 52894 12414 52946
rect 8654 52882 8706 52894
rect 10334 52882 10386 52894
rect 12686 52882 12738 52894
rect 14926 52946 14978 52958
rect 31614 52946 31666 52958
rect 17490 52894 17502 52946
rect 17554 52894 17566 52946
rect 20626 52894 20638 52946
rect 20690 52894 20702 52946
rect 24210 52894 24222 52946
rect 24274 52894 24286 52946
rect 14926 52882 14978 52894
rect 31614 52882 31666 52894
rect 32174 52946 32226 52958
rect 34414 52946 34466 52958
rect 36766 52946 36818 52958
rect 54126 52946 54178 52958
rect 33730 52894 33742 52946
rect 33794 52894 33806 52946
rect 35634 52894 35646 52946
rect 35698 52894 35710 52946
rect 35970 52894 35982 52946
rect 36034 52894 36046 52946
rect 42466 52894 42478 52946
rect 42530 52894 42542 52946
rect 46386 52894 46398 52946
rect 46450 52894 46462 52946
rect 47058 52894 47070 52946
rect 47122 52894 47134 52946
rect 50754 52894 50766 52946
rect 50818 52894 50830 52946
rect 32174 52882 32226 52894
rect 34414 52882 34466 52894
rect 36766 52882 36818 52894
rect 54126 52882 54178 52894
rect 54462 52946 54514 52958
rect 54462 52882 54514 52894
rect 58158 52946 58210 52958
rect 58158 52882 58210 52894
rect 9774 52834 9826 52846
rect 8082 52782 8094 52834
rect 8146 52782 8158 52834
rect 9774 52770 9826 52782
rect 10110 52834 10162 52846
rect 10110 52770 10162 52782
rect 10670 52834 10722 52846
rect 13694 52834 13746 52846
rect 31950 52834 32002 52846
rect 41022 52834 41074 52846
rect 57374 52834 57426 52846
rect 11106 52782 11118 52834
rect 11170 52782 11182 52834
rect 20290 52782 20302 52834
rect 20354 52782 20366 52834
rect 23538 52782 23550 52834
rect 23602 52782 23614 52834
rect 33506 52782 33518 52834
rect 33570 52782 33582 52834
rect 43250 52782 43262 52834
rect 43314 52782 43326 52834
rect 45378 52782 45390 52834
rect 45442 52782 45454 52834
rect 46498 52782 46510 52834
rect 46562 52782 46574 52834
rect 53666 52782 53678 52834
rect 53730 52782 53742 52834
rect 10670 52770 10722 52782
rect 13694 52770 13746 52782
rect 31950 52770 32002 52782
rect 41022 52770 41074 52782
rect 57374 52770 57426 52782
rect 57598 52834 57650 52846
rect 57598 52770 57650 52782
rect 54014 52722 54066 52734
rect 13122 52670 13134 52722
rect 13186 52670 13198 52722
rect 32498 52670 32510 52722
rect 32562 52670 32574 52722
rect 45602 52670 45614 52722
rect 45666 52719 45678 52722
rect 46162 52719 46174 52722
rect 45666 52673 46174 52719
rect 45666 52670 45678 52673
rect 46162 52670 46174 52673
rect 46226 52670 46238 52722
rect 47282 52670 47294 52722
rect 47346 52719 47358 52722
rect 47618 52719 47630 52722
rect 47346 52673 47630 52719
rect 47346 52670 47358 52673
rect 47618 52670 47630 52673
rect 47682 52670 47694 52722
rect 54014 52658 54066 52670
rect 54350 52722 54402 52734
rect 54350 52658 54402 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 8766 52386 8818 52398
rect 8766 52322 8818 52334
rect 15710 52386 15762 52398
rect 15710 52322 15762 52334
rect 16158 52386 16210 52398
rect 20414 52386 20466 52398
rect 55918 52386 55970 52398
rect 16482 52334 16494 52386
rect 16546 52334 16558 52386
rect 20738 52334 20750 52386
rect 20802 52334 20814 52386
rect 36082 52334 36094 52386
rect 36146 52334 36158 52386
rect 16158 52322 16210 52334
rect 20414 52322 20466 52334
rect 55918 52322 55970 52334
rect 56142 52386 56194 52398
rect 56142 52322 56194 52334
rect 56254 52386 56306 52398
rect 56254 52322 56306 52334
rect 7310 52274 7362 52286
rect 12350 52274 12402 52286
rect 8194 52222 8206 52274
rect 8258 52222 8270 52274
rect 7310 52210 7362 52222
rect 12350 52210 12402 52222
rect 18510 52274 18562 52286
rect 20190 52274 20242 52286
rect 19394 52222 19406 52274
rect 19458 52222 19470 52274
rect 18510 52210 18562 52222
rect 20190 52210 20242 52222
rect 21534 52274 21586 52286
rect 32398 52274 32450 52286
rect 35982 52274 36034 52286
rect 24546 52222 24558 52274
rect 24610 52222 24622 52274
rect 33618 52222 33630 52274
rect 33682 52222 33694 52274
rect 21534 52210 21586 52222
rect 32398 52210 32450 52222
rect 35982 52210 36034 52222
rect 39454 52274 39506 52286
rect 39454 52210 39506 52222
rect 43262 52274 43314 52286
rect 51774 52274 51826 52286
rect 46722 52222 46734 52274
rect 46786 52222 46798 52274
rect 47618 52222 47630 52274
rect 47682 52222 47694 52274
rect 51202 52222 51214 52274
rect 51266 52222 51278 52274
rect 43262 52210 43314 52222
rect 51774 52210 51826 52222
rect 4622 52162 4674 52174
rect 8654 52162 8706 52174
rect 7970 52110 7982 52162
rect 8034 52110 8046 52162
rect 4622 52098 4674 52110
rect 8654 52098 8706 52110
rect 9662 52162 9714 52174
rect 12910 52162 12962 52174
rect 10210 52110 10222 52162
rect 10274 52110 10286 52162
rect 9662 52098 9714 52110
rect 12910 52098 12962 52110
rect 13582 52162 13634 52174
rect 14478 52162 14530 52174
rect 13906 52110 13918 52162
rect 13970 52110 13982 52162
rect 13582 52098 13634 52110
rect 14478 52098 14530 52110
rect 14814 52162 14866 52174
rect 14814 52098 14866 52110
rect 15038 52162 15090 52174
rect 15038 52098 15090 52110
rect 15262 52162 15314 52174
rect 15262 52098 15314 52110
rect 15934 52162 15986 52174
rect 32286 52162 32338 52174
rect 38894 52162 38946 52174
rect 19170 52110 19182 52162
rect 19234 52110 19246 52162
rect 23090 52110 23102 52162
rect 23154 52110 23166 52162
rect 30930 52110 30942 52162
rect 30994 52110 31006 52162
rect 31938 52110 31950 52162
rect 32002 52110 32014 52162
rect 32722 52110 32734 52162
rect 32786 52110 32798 52162
rect 33282 52110 33294 52162
rect 33346 52110 33358 52162
rect 35634 52110 35646 52162
rect 35698 52110 35710 52162
rect 15934 52098 15986 52110
rect 32286 52098 32338 52110
rect 38894 52098 38946 52110
rect 43822 52162 43874 52174
rect 54126 52162 54178 52174
rect 46610 52110 46622 52162
rect 46674 52110 46686 52162
rect 50530 52110 50542 52162
rect 50594 52110 50606 52162
rect 50978 52110 50990 52162
rect 51042 52110 51054 52162
rect 43822 52098 43874 52110
rect 54126 52098 54178 52110
rect 8766 52050 8818 52062
rect 37662 52050 37714 52062
rect 9986 51998 9998 52050
rect 10050 51998 10062 52050
rect 11442 51998 11454 52050
rect 11506 51998 11518 52050
rect 24322 51998 24334 52050
rect 24386 51998 24398 52050
rect 30706 51998 30718 52050
rect 30770 51998 30782 52050
rect 33730 51998 33742 52050
rect 33794 51998 33806 52050
rect 8766 51986 8818 51998
rect 37662 51986 37714 51998
rect 43150 52050 43202 52062
rect 43150 51986 43202 51998
rect 44158 52050 44210 52062
rect 44158 51986 44210 51998
rect 47070 52050 47122 52062
rect 47070 51986 47122 51998
rect 47294 52050 47346 52062
rect 49746 51998 49758 52050
rect 49810 51998 49822 52050
rect 47294 51986 47346 51998
rect 11790 51938 11842 51950
rect 11790 51874 11842 51886
rect 12238 51938 12290 51950
rect 12238 51874 12290 51886
rect 12462 51938 12514 51950
rect 37998 51938 38050 51950
rect 22530 51886 22542 51938
rect 22594 51886 22606 51938
rect 12462 51874 12514 51886
rect 37998 51874 38050 51886
rect 43374 51938 43426 51950
rect 43374 51874 43426 51886
rect 46846 51938 46898 51950
rect 56254 51938 56306 51950
rect 54450 51886 54462 51938
rect 54514 51886 54526 51938
rect 46846 51874 46898 51886
rect 56254 51874 56306 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 12910 51602 12962 51614
rect 12910 51538 12962 51550
rect 13134 51602 13186 51614
rect 13134 51538 13186 51550
rect 13358 51602 13410 51614
rect 13358 51538 13410 51550
rect 32510 51602 32562 51614
rect 43262 51602 43314 51614
rect 36306 51550 36318 51602
rect 36370 51550 36382 51602
rect 32510 51538 32562 51550
rect 43262 51538 43314 51550
rect 47182 51602 47234 51614
rect 47182 51538 47234 51550
rect 48302 51602 48354 51614
rect 48302 51538 48354 51550
rect 48862 51602 48914 51614
rect 48862 51538 48914 51550
rect 51886 51602 51938 51614
rect 56702 51602 56754 51614
rect 52770 51550 52782 51602
rect 52834 51550 52846 51602
rect 55906 51550 55918 51602
rect 55970 51550 55982 51602
rect 51886 51538 51938 51550
rect 56702 51538 56754 51550
rect 3390 51490 3442 51502
rect 13470 51490 13522 51502
rect 5394 51438 5406 51490
rect 5458 51438 5470 51490
rect 3390 51426 3442 51438
rect 13470 51426 13522 51438
rect 15038 51490 15090 51502
rect 38670 51490 38722 51502
rect 37314 51438 37326 51490
rect 37378 51438 37390 51490
rect 15038 51426 15090 51438
rect 38670 51426 38722 51438
rect 41022 51490 41074 51502
rect 41022 51426 41074 51438
rect 41582 51490 41634 51502
rect 41582 51426 41634 51438
rect 41694 51490 41746 51502
rect 41694 51426 41746 51438
rect 48750 51490 48802 51502
rect 48750 51426 48802 51438
rect 53230 51490 53282 51502
rect 53230 51426 53282 51438
rect 55470 51490 55522 51502
rect 55470 51426 55522 51438
rect 3278 51378 3330 51390
rect 3278 51314 3330 51326
rect 3614 51378 3666 51390
rect 4174 51378 4226 51390
rect 3826 51326 3838 51378
rect 3890 51326 3902 51378
rect 3614 51314 3666 51326
rect 4174 51314 4226 51326
rect 4398 51378 4450 51390
rect 14590 51378 14642 51390
rect 5058 51326 5070 51378
rect 5122 51326 5134 51378
rect 5730 51326 5742 51378
rect 5794 51326 5806 51378
rect 4398 51314 4450 51326
rect 14590 51314 14642 51326
rect 15262 51378 15314 51390
rect 15262 51314 15314 51326
rect 28478 51378 28530 51390
rect 47294 51378 47346 51390
rect 29250 51326 29262 51378
rect 29314 51326 29326 51378
rect 30034 51326 30046 51378
rect 30098 51326 30110 51378
rect 36194 51326 36206 51378
rect 36258 51326 36270 51378
rect 36754 51326 36766 51378
rect 36818 51326 36830 51378
rect 37986 51326 37998 51378
rect 38050 51326 38062 51378
rect 43698 51326 43710 51378
rect 43762 51326 43774 51378
rect 46946 51326 46958 51378
rect 47010 51326 47022 51378
rect 28478 51314 28530 51326
rect 47294 51314 47346 51326
rect 47630 51378 47682 51390
rect 52446 51378 52498 51390
rect 55358 51378 55410 51390
rect 52098 51326 52110 51378
rect 52162 51326 52174 51378
rect 55122 51326 55134 51378
rect 55186 51326 55198 51378
rect 47630 51314 47682 51326
rect 52446 51314 52498 51326
rect 55358 51314 55410 51326
rect 56478 51378 56530 51390
rect 56478 51314 56530 51326
rect 56814 51378 56866 51390
rect 56814 51314 56866 51326
rect 57038 51378 57090 51390
rect 57038 51314 57090 51326
rect 4286 51266 4338 51278
rect 15150 51266 15202 51278
rect 42254 51266 42306 51278
rect 47854 51266 47906 51278
rect 5506 51214 5518 51266
rect 5570 51214 5582 51266
rect 29698 51214 29710 51266
rect 29762 51214 29774 51266
rect 37762 51214 37774 51266
rect 37826 51214 37838 51266
rect 44370 51214 44382 51266
rect 44434 51214 44446 51266
rect 46498 51214 46510 51266
rect 46562 51214 46574 51266
rect 4286 51202 4338 51214
rect 15150 51202 15202 51214
rect 42254 51202 42306 51214
rect 47854 51202 47906 51214
rect 48190 51266 48242 51278
rect 48190 51202 48242 51214
rect 28590 51154 28642 51166
rect 28590 51090 28642 51102
rect 29822 51154 29874 51166
rect 29822 51090 29874 51102
rect 40910 51154 40962 51166
rect 40910 51090 40962 51102
rect 41246 51154 41298 51166
rect 41246 51090 41298 51102
rect 41694 51154 41746 51166
rect 41694 51090 41746 51102
rect 51774 51154 51826 51166
rect 51774 51090 51826 51102
rect 53118 51154 53170 51166
rect 53118 51090 53170 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 5070 50818 5122 50830
rect 5070 50754 5122 50766
rect 5742 50818 5794 50830
rect 5742 50754 5794 50766
rect 14366 50818 14418 50830
rect 14366 50754 14418 50766
rect 41806 50818 41858 50830
rect 41806 50754 41858 50766
rect 44942 50706 44994 50718
rect 4610 50654 4622 50706
rect 4674 50654 4686 50706
rect 9314 50654 9326 50706
rect 9378 50654 9390 50706
rect 11554 50654 11566 50706
rect 11618 50654 11630 50706
rect 28354 50654 28366 50706
rect 28418 50654 28430 50706
rect 29698 50654 29710 50706
rect 29762 50654 29774 50706
rect 33170 50654 33182 50706
rect 33234 50654 33246 50706
rect 35186 50654 35198 50706
rect 35250 50654 35262 50706
rect 36306 50654 36318 50706
rect 36370 50654 36382 50706
rect 38546 50654 38558 50706
rect 38610 50654 38622 50706
rect 40674 50654 40686 50706
rect 40738 50654 40750 50706
rect 56018 50654 56030 50706
rect 56082 50654 56094 50706
rect 58146 50654 58158 50706
rect 58210 50654 58222 50706
rect 44942 50642 44994 50654
rect 4958 50594 5010 50606
rect 1810 50542 1822 50594
rect 1874 50542 1886 50594
rect 4958 50530 5010 50542
rect 5630 50594 5682 50606
rect 30158 50594 30210 50606
rect 9202 50542 9214 50594
rect 9266 50542 9278 50594
rect 9874 50542 9886 50594
rect 9938 50542 9950 50594
rect 25442 50542 25454 50594
rect 25506 50542 25518 50594
rect 29474 50542 29486 50594
rect 29538 50542 29550 50594
rect 5630 50530 5682 50542
rect 30158 50530 30210 50542
rect 30382 50594 30434 50606
rect 30382 50530 30434 50542
rect 30718 50594 30770 50606
rect 30718 50530 30770 50542
rect 30942 50594 30994 50606
rect 41918 50594 41970 50606
rect 32274 50542 32286 50594
rect 32338 50542 32350 50594
rect 32498 50542 32510 50594
rect 32562 50542 32574 50594
rect 33282 50542 33294 50594
rect 33346 50542 33358 50594
rect 35074 50542 35086 50594
rect 35138 50542 35150 50594
rect 41458 50542 41470 50594
rect 41522 50542 41534 50594
rect 30942 50530 30994 50542
rect 41918 50530 41970 50542
rect 42142 50594 42194 50606
rect 42142 50530 42194 50542
rect 42254 50594 42306 50606
rect 42254 50530 42306 50542
rect 42814 50594 42866 50606
rect 42814 50530 42866 50542
rect 44830 50594 44882 50606
rect 44830 50530 44882 50542
rect 45502 50594 45554 50606
rect 45502 50530 45554 50542
rect 45838 50594 45890 50606
rect 47182 50594 47234 50606
rect 46722 50542 46734 50594
rect 46786 50542 46798 50594
rect 47394 50542 47406 50594
rect 47458 50542 47470 50594
rect 55234 50542 55246 50594
rect 55298 50542 55310 50594
rect 45838 50530 45890 50542
rect 47182 50530 47234 50542
rect 5742 50482 5794 50494
rect 10782 50482 10834 50494
rect 2482 50430 2494 50482
rect 2546 50430 2558 50482
rect 8866 50430 8878 50482
rect 8930 50430 8942 50482
rect 5742 50418 5794 50430
rect 10782 50418 10834 50430
rect 11118 50482 11170 50494
rect 11118 50418 11170 50430
rect 14030 50482 14082 50494
rect 14030 50418 14082 50430
rect 19630 50482 19682 50494
rect 19630 50418 19682 50430
rect 25118 50482 25170 50494
rect 30606 50482 30658 50494
rect 26226 50430 26238 50482
rect 26290 50430 26302 50482
rect 25118 50418 25170 50430
rect 30606 50418 30658 50430
rect 47854 50482 47906 50494
rect 47854 50418 47906 50430
rect 13694 50370 13746 50382
rect 13694 50306 13746 50318
rect 14254 50370 14306 50382
rect 14254 50306 14306 50318
rect 19742 50370 19794 50382
rect 19742 50306 19794 50318
rect 45054 50370 45106 50382
rect 45054 50306 45106 50318
rect 46958 50370 47010 50382
rect 46958 50306 47010 50318
rect 47070 50370 47122 50382
rect 47070 50306 47122 50318
rect 54910 50370 54962 50382
rect 54910 50306 54962 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 4510 50034 4562 50046
rect 4510 49970 4562 49982
rect 9438 50034 9490 50046
rect 9438 49970 9490 49982
rect 28478 50034 28530 50046
rect 28478 49970 28530 49982
rect 29374 50034 29426 50046
rect 29374 49970 29426 49982
rect 29486 50034 29538 50046
rect 29486 49970 29538 49982
rect 29934 50034 29986 50046
rect 29934 49970 29986 49982
rect 30158 50034 30210 50046
rect 30158 49970 30210 49982
rect 30494 50034 30546 50046
rect 41022 50034 41074 50046
rect 35410 49982 35422 50034
rect 35474 49982 35486 50034
rect 30494 49970 30546 49982
rect 41022 49970 41074 49982
rect 50878 50034 50930 50046
rect 50878 49970 50930 49982
rect 51102 50034 51154 50046
rect 51102 49970 51154 49982
rect 4062 49922 4114 49934
rect 4062 49858 4114 49870
rect 9662 49922 9714 49934
rect 9662 49858 9714 49870
rect 10222 49922 10274 49934
rect 10222 49858 10274 49870
rect 19294 49922 19346 49934
rect 21534 49922 21586 49934
rect 20402 49870 20414 49922
rect 20466 49870 20478 49922
rect 19294 49858 19346 49870
rect 21534 49858 21586 49870
rect 28366 49922 28418 49934
rect 28366 49858 28418 49870
rect 34078 49922 34130 49934
rect 39342 49922 39394 49934
rect 37762 49870 37774 49922
rect 37826 49870 37838 49922
rect 34078 49858 34130 49870
rect 39342 49858 39394 49870
rect 41918 49922 41970 49934
rect 41918 49858 41970 49870
rect 47294 49922 47346 49934
rect 47294 49858 47346 49870
rect 50766 49922 50818 49934
rect 50766 49858 50818 49870
rect 52222 49922 52274 49934
rect 52222 49858 52274 49870
rect 3950 49810 4002 49822
rect 3378 49758 3390 49810
rect 3442 49758 3454 49810
rect 3950 49746 4002 49758
rect 4286 49810 4338 49822
rect 4286 49746 4338 49758
rect 4734 49810 4786 49822
rect 4734 49746 4786 49758
rect 4846 49810 4898 49822
rect 8878 49810 8930 49822
rect 8642 49758 8654 49810
rect 8706 49758 8718 49810
rect 4846 49746 4898 49758
rect 8878 49746 8930 49758
rect 9774 49810 9826 49822
rect 9774 49746 9826 49758
rect 9998 49810 10050 49822
rect 9998 49746 10050 49758
rect 10334 49810 10386 49822
rect 10334 49746 10386 49758
rect 12686 49810 12738 49822
rect 12686 49746 12738 49758
rect 13246 49810 13298 49822
rect 14814 49810 14866 49822
rect 14354 49758 14366 49810
rect 14418 49758 14430 49810
rect 13246 49746 13298 49758
rect 14814 49746 14866 49758
rect 19182 49810 19234 49822
rect 21422 49810 21474 49822
rect 28702 49810 28754 49822
rect 20290 49758 20302 49810
rect 20354 49758 20366 49810
rect 21186 49758 21198 49810
rect 21250 49758 21262 49810
rect 23762 49758 23774 49810
rect 23826 49758 23838 49810
rect 19182 49746 19234 49758
rect 21422 49746 21474 49758
rect 28702 49746 28754 49758
rect 28814 49810 28866 49822
rect 28814 49746 28866 49758
rect 29262 49810 29314 49822
rect 29262 49746 29314 49758
rect 29822 49810 29874 49822
rect 35086 49810 35138 49822
rect 41246 49810 41298 49822
rect 31490 49758 31502 49810
rect 31554 49758 31566 49810
rect 32050 49758 32062 49810
rect 32114 49758 32126 49810
rect 33394 49758 33406 49810
rect 33458 49758 33470 49810
rect 38658 49758 38670 49810
rect 38722 49758 38734 49810
rect 29822 49746 29874 49758
rect 35086 49746 35138 49758
rect 41246 49746 41298 49758
rect 41358 49810 41410 49822
rect 41358 49746 41410 49758
rect 41470 49810 41522 49822
rect 41470 49746 41522 49758
rect 51998 49810 52050 49822
rect 51998 49746 52050 49758
rect 52670 49810 52722 49822
rect 52670 49746 52722 49758
rect 5406 49698 5458 49710
rect 5406 49634 5458 49646
rect 7982 49698 8034 49710
rect 7982 49634 8034 49646
rect 12350 49698 12402 49710
rect 34862 49698 34914 49710
rect 42142 49698 42194 49710
rect 13906 49646 13918 49698
rect 13970 49646 13982 49698
rect 20514 49646 20526 49698
rect 20578 49646 20590 49698
rect 23650 49646 23662 49698
rect 23714 49646 23726 49698
rect 31154 49646 31166 49698
rect 31218 49646 31230 49698
rect 32386 49646 32398 49698
rect 32450 49646 32462 49698
rect 33730 49646 33742 49698
rect 33794 49646 33806 49698
rect 37202 49646 37214 49698
rect 37266 49646 37278 49698
rect 41794 49646 41806 49698
rect 41858 49646 41870 49698
rect 12350 49634 12402 49646
rect 34862 49634 34914 49646
rect 42142 49634 42194 49646
rect 49870 49698 49922 49710
rect 49870 49634 49922 49646
rect 50430 49698 50482 49710
rect 50430 49634 50482 49646
rect 51662 49698 51714 49710
rect 51662 49634 51714 49646
rect 52446 49698 52498 49710
rect 52446 49634 52498 49646
rect 19294 49586 19346 49598
rect 19294 49522 19346 49534
rect 21534 49586 21586 49598
rect 21534 49522 21586 49534
rect 23438 49586 23490 49598
rect 23438 49522 23490 49534
rect 47406 49586 47458 49598
rect 47406 49522 47458 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 33294 49250 33346 49262
rect 33294 49186 33346 49198
rect 53006 49250 53058 49262
rect 53006 49186 53058 49198
rect 10222 49138 10274 49150
rect 22542 49138 22594 49150
rect 32734 49138 32786 49150
rect 8866 49086 8878 49138
rect 8930 49086 8942 49138
rect 16258 49086 16270 49138
rect 16322 49086 16334 49138
rect 19506 49086 19518 49138
rect 19570 49086 19582 49138
rect 23650 49086 23662 49138
rect 23714 49086 23726 49138
rect 25778 49086 25790 49138
rect 25842 49086 25854 49138
rect 10222 49074 10274 49086
rect 22542 49074 22594 49086
rect 32734 49074 32786 49086
rect 32958 49138 33010 49150
rect 32958 49074 33010 49086
rect 33742 49138 33794 49150
rect 33742 49074 33794 49086
rect 42142 49138 42194 49150
rect 46722 49086 46734 49138
rect 46786 49086 46798 49138
rect 48850 49086 48862 49138
rect 48914 49086 48926 49138
rect 50754 49086 50766 49138
rect 50818 49086 50830 49138
rect 58146 49086 58158 49138
rect 58210 49086 58222 49138
rect 42142 49074 42194 49086
rect 9102 49026 9154 49038
rect 6066 48974 6078 49026
rect 6130 48974 6142 49026
rect 9102 48962 9154 48974
rect 9662 49026 9714 49038
rect 21982 49026 22034 49038
rect 32174 49026 32226 49038
rect 15026 48974 15038 49026
rect 15090 48974 15102 49026
rect 15586 48974 15598 49026
rect 15650 48974 15662 49026
rect 16706 48974 16718 49026
rect 16770 48974 16782 49026
rect 22978 48974 22990 49026
rect 23042 48974 23054 49026
rect 31490 48974 31502 49026
rect 31554 48974 31566 49026
rect 9662 48962 9714 48974
rect 21982 48962 22034 48974
rect 32174 48962 32226 48974
rect 32398 49026 32450 49038
rect 32398 48962 32450 48974
rect 41918 49026 41970 49038
rect 41918 48962 41970 48974
rect 42030 49026 42082 49038
rect 42030 48962 42082 48974
rect 42254 49026 42306 49038
rect 42254 48962 42306 48974
rect 42814 49026 42866 49038
rect 50654 49026 50706 49038
rect 49634 48974 49646 49026
rect 49698 48974 49710 49026
rect 42814 48962 42866 48974
rect 50654 48962 50706 48974
rect 51550 49026 51602 49038
rect 51550 48962 51602 48974
rect 52782 49026 52834 49038
rect 54910 49026 54962 49038
rect 53218 48974 53230 49026
rect 53282 48974 53294 49026
rect 54114 48974 54126 49026
rect 54178 48974 54190 49026
rect 54450 48974 54462 49026
rect 54514 48974 54526 49026
rect 55234 48974 55246 49026
rect 55298 48974 55310 49026
rect 52782 48962 52834 48974
rect 54910 48962 54962 48974
rect 9326 48914 9378 48926
rect 6738 48862 6750 48914
rect 6802 48862 6814 48914
rect 9326 48850 9378 48862
rect 9550 48914 9602 48926
rect 9550 48850 9602 48862
rect 11118 48914 11170 48926
rect 20078 48914 20130 48926
rect 17378 48862 17390 48914
rect 17442 48862 17454 48914
rect 11118 48850 11170 48862
rect 20078 48850 20130 48862
rect 20190 48914 20242 48926
rect 20190 48850 20242 48862
rect 20414 48914 20466 48926
rect 20414 48850 20466 48862
rect 20638 48914 20690 48926
rect 20638 48850 20690 48862
rect 21422 48914 21474 48926
rect 21422 48850 21474 48862
rect 43150 48914 43202 48926
rect 56018 48862 56030 48914
rect 56082 48862 56094 48914
rect 43150 48850 43202 48862
rect 11230 48802 11282 48814
rect 11230 48738 11282 48750
rect 11342 48802 11394 48814
rect 11342 48738 11394 48750
rect 21310 48802 21362 48814
rect 21310 48738 21362 48750
rect 21534 48802 21586 48814
rect 21534 48738 21586 48750
rect 42366 48802 42418 48814
rect 42366 48738 42418 48750
rect 43038 48802 43090 48814
rect 43038 48738 43090 48750
rect 50990 48802 51042 48814
rect 50990 48738 51042 48750
rect 52110 48802 52162 48814
rect 52110 48738 52162 48750
rect 53118 48802 53170 48814
rect 53118 48738 53170 48750
rect 53902 48802 53954 48814
rect 53902 48738 53954 48750
rect 54686 48802 54738 48814
rect 54686 48738 54738 48750
rect 54798 48802 54850 48814
rect 54798 48738 54850 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 8318 48466 8370 48478
rect 8318 48402 8370 48414
rect 8430 48466 8482 48478
rect 8430 48402 8482 48414
rect 8542 48466 8594 48478
rect 8542 48402 8594 48414
rect 19070 48466 19122 48478
rect 24446 48466 24498 48478
rect 22082 48414 22094 48466
rect 22146 48414 22158 48466
rect 19070 48402 19122 48414
rect 24446 48402 24498 48414
rect 27358 48466 27410 48478
rect 27358 48402 27410 48414
rect 32510 48466 32562 48478
rect 32510 48402 32562 48414
rect 41694 48466 41746 48478
rect 41694 48402 41746 48414
rect 42478 48466 42530 48478
rect 42478 48402 42530 48414
rect 55918 48466 55970 48478
rect 55918 48402 55970 48414
rect 6190 48354 6242 48366
rect 4834 48302 4846 48354
rect 4898 48302 4910 48354
rect 6190 48290 6242 48302
rect 8094 48354 8146 48366
rect 8094 48290 8146 48302
rect 8878 48354 8930 48366
rect 13582 48354 13634 48366
rect 20414 48354 20466 48366
rect 28366 48354 28418 48366
rect 42366 48354 42418 48366
rect 10546 48302 10558 48354
rect 10610 48302 10622 48354
rect 15250 48302 15262 48354
rect 15314 48302 15326 48354
rect 15698 48302 15710 48354
rect 15762 48302 15774 48354
rect 23650 48302 23662 48354
rect 23714 48302 23726 48354
rect 37202 48302 37214 48354
rect 37266 48302 37278 48354
rect 8878 48290 8930 48302
rect 13582 48290 13634 48302
rect 20414 48290 20466 48302
rect 28366 48290 28418 48302
rect 42366 48290 42418 48302
rect 43374 48354 43426 48366
rect 55470 48354 55522 48366
rect 52994 48302 53006 48354
rect 53058 48302 53070 48354
rect 43374 48290 43426 48302
rect 55470 48290 55522 48302
rect 55694 48354 55746 48366
rect 55694 48290 55746 48302
rect 5966 48242 6018 48254
rect 4722 48190 4734 48242
rect 4786 48190 4798 48242
rect 5730 48190 5742 48242
rect 5794 48190 5806 48242
rect 5966 48178 6018 48190
rect 6302 48242 6354 48254
rect 13358 48242 13410 48254
rect 27246 48242 27298 48254
rect 11106 48190 11118 48242
rect 11170 48190 11182 48242
rect 11778 48190 11790 48242
rect 11842 48190 11854 48242
rect 14802 48190 14814 48242
rect 14866 48190 14878 48242
rect 15922 48190 15934 48242
rect 15986 48190 15998 48242
rect 19954 48190 19966 48242
rect 20018 48190 20030 48242
rect 22418 48190 22430 48242
rect 22482 48190 22494 48242
rect 6302 48178 6354 48190
rect 13358 48178 13410 48190
rect 27246 48178 27298 48190
rect 27470 48242 27522 48254
rect 27470 48178 27522 48190
rect 27918 48242 27970 48254
rect 27918 48178 27970 48190
rect 28254 48242 28306 48254
rect 43262 48242 43314 48254
rect 35970 48190 35982 48242
rect 36034 48190 36046 48242
rect 37090 48190 37102 48242
rect 37154 48190 37166 48242
rect 28254 48178 28306 48190
rect 43262 48178 43314 48190
rect 43486 48242 43538 48254
rect 43486 48178 43538 48190
rect 43934 48242 43986 48254
rect 43934 48178 43986 48190
rect 49198 48242 49250 48254
rect 49198 48178 49250 48190
rect 50094 48242 50146 48254
rect 56142 48242 56194 48254
rect 53666 48190 53678 48242
rect 53730 48190 53742 48242
rect 50094 48178 50146 48190
rect 56142 48178 56194 48190
rect 8990 48130 9042 48142
rect 5170 48078 5182 48130
rect 5234 48078 5246 48130
rect 8990 48066 9042 48078
rect 12462 48130 12514 48142
rect 20974 48130 21026 48142
rect 13682 48078 13694 48130
rect 13746 48078 13758 48130
rect 15138 48078 15150 48130
rect 15202 48078 15214 48130
rect 19618 48078 19630 48130
rect 19682 48078 19694 48130
rect 12462 48066 12514 48078
rect 20974 48066 21026 48078
rect 23774 48130 23826 48142
rect 41582 48130 41634 48142
rect 36642 48078 36654 48130
rect 36706 48078 36718 48130
rect 23774 48066 23826 48078
rect 41582 48066 41634 48078
rect 48862 48130 48914 48142
rect 54238 48130 54290 48142
rect 49634 48078 49646 48130
rect 49698 48078 49710 48130
rect 50866 48078 50878 48130
rect 50930 48078 50942 48130
rect 48862 48066 48914 48078
rect 54238 48066 54290 48078
rect 54910 48130 54962 48142
rect 54910 48066 54962 48078
rect 24334 48018 24386 48030
rect 24334 47954 24386 47966
rect 24670 48018 24722 48030
rect 24670 47954 24722 47966
rect 28366 48018 28418 48030
rect 28366 47954 28418 47966
rect 42478 48018 42530 48030
rect 42478 47954 42530 47966
rect 50206 48018 50258 48030
rect 50206 47954 50258 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 5630 47682 5682 47694
rect 29374 47682 29426 47694
rect 11106 47630 11118 47682
rect 11170 47630 11182 47682
rect 22642 47630 22654 47682
rect 22706 47630 22718 47682
rect 35410 47630 35422 47682
rect 35474 47630 35486 47682
rect 5630 47618 5682 47630
rect 29374 47618 29426 47630
rect 5070 47570 5122 47582
rect 16270 47570 16322 47582
rect 44270 47570 44322 47582
rect 49758 47570 49810 47582
rect 4610 47518 4622 47570
rect 4674 47518 4686 47570
rect 11218 47518 11230 47570
rect 11282 47518 11294 47570
rect 19058 47518 19070 47570
rect 19122 47518 19134 47570
rect 23090 47518 23102 47570
rect 23154 47518 23166 47570
rect 25778 47518 25790 47570
rect 25842 47518 25854 47570
rect 28466 47518 28478 47570
rect 28530 47518 28542 47570
rect 34626 47518 34638 47570
rect 34690 47518 34702 47570
rect 37426 47518 37438 47570
rect 37490 47518 37502 47570
rect 47730 47518 47742 47570
rect 47794 47518 47806 47570
rect 5070 47506 5122 47518
rect 16270 47506 16322 47518
rect 44270 47506 44322 47518
rect 49758 47506 49810 47518
rect 13358 47458 13410 47470
rect 1810 47406 1822 47458
rect 1874 47406 1886 47458
rect 11106 47406 11118 47458
rect 11170 47406 11182 47458
rect 12226 47406 12238 47458
rect 12290 47406 12302 47458
rect 13358 47394 13410 47406
rect 13694 47458 13746 47470
rect 13694 47394 13746 47406
rect 14030 47458 14082 47470
rect 14030 47394 14082 47406
rect 15822 47458 15874 47470
rect 15822 47394 15874 47406
rect 16046 47458 16098 47470
rect 16046 47394 16098 47406
rect 16382 47458 16434 47470
rect 16382 47394 16434 47406
rect 16606 47458 16658 47470
rect 18174 47458 18226 47470
rect 24558 47458 24610 47470
rect 38110 47458 38162 47470
rect 56254 47458 56306 47470
rect 17602 47406 17614 47458
rect 17666 47406 17678 47458
rect 22866 47406 22878 47458
rect 22930 47406 22942 47458
rect 23650 47406 23662 47458
rect 23714 47406 23726 47458
rect 27458 47406 27470 47458
rect 27522 47406 27534 47458
rect 34738 47406 34750 47458
rect 34802 47406 34814 47458
rect 37650 47406 37662 47458
rect 37714 47406 37726 47458
rect 38434 47406 38446 47458
rect 38498 47406 38510 47458
rect 38994 47406 39006 47458
rect 39058 47406 39070 47458
rect 41682 47406 41694 47458
rect 41746 47406 41758 47458
rect 42466 47406 42478 47458
rect 42530 47406 42542 47458
rect 44818 47406 44830 47458
rect 44882 47406 44894 47458
rect 52658 47406 52670 47458
rect 52722 47406 52734 47458
rect 16606 47394 16658 47406
rect 18174 47394 18226 47406
rect 24558 47394 24610 47406
rect 38110 47394 38162 47406
rect 56254 47394 56306 47406
rect 5742 47346 5794 47358
rect 2482 47294 2494 47346
rect 2546 47294 2558 47346
rect 5742 47282 5794 47294
rect 5966 47346 6018 47358
rect 5966 47282 6018 47294
rect 12574 47346 12626 47358
rect 12574 47282 12626 47294
rect 12910 47346 12962 47358
rect 12910 47282 12962 47294
rect 13582 47346 13634 47358
rect 13582 47282 13634 47294
rect 15486 47346 15538 47358
rect 15486 47282 15538 47294
rect 18286 47346 18338 47358
rect 24894 47346 24946 47358
rect 23986 47294 23998 47346
rect 24050 47294 24062 47346
rect 26114 47294 26126 47346
rect 26178 47294 26190 47346
rect 39106 47294 39118 47346
rect 39170 47294 39182 47346
rect 42578 47294 42590 47346
rect 42642 47294 42654 47346
rect 45602 47294 45614 47346
rect 45666 47294 45678 47346
rect 53442 47294 53454 47346
rect 53506 47294 53518 47346
rect 18286 47282 18338 47294
rect 24894 47282 24946 47294
rect 14590 47234 14642 47246
rect 14590 47170 14642 47182
rect 18622 47234 18674 47246
rect 18622 47170 18674 47182
rect 24334 47234 24386 47246
rect 24334 47170 24386 47182
rect 24782 47234 24834 47246
rect 24782 47170 24834 47182
rect 25454 47234 25506 47246
rect 25454 47170 25506 47182
rect 29486 47234 29538 47246
rect 29486 47170 29538 47182
rect 29598 47234 29650 47246
rect 48526 47234 48578 47246
rect 38546 47182 38558 47234
rect 38610 47182 38622 47234
rect 41346 47182 41358 47234
rect 41410 47182 41422 47234
rect 55682 47182 55694 47234
rect 55746 47182 55758 47234
rect 29598 47170 29650 47182
rect 48526 47170 48578 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 2606 46898 2658 46910
rect 32510 46898 32562 46910
rect 36094 46898 36146 46910
rect 24546 46846 24558 46898
rect 24610 46846 24622 46898
rect 27234 46846 27246 46898
rect 27298 46846 27310 46898
rect 35298 46846 35310 46898
rect 35362 46846 35374 46898
rect 2606 46834 2658 46846
rect 32510 46834 32562 46846
rect 36094 46834 36146 46846
rect 36430 46898 36482 46910
rect 36430 46834 36482 46846
rect 45950 46898 46002 46910
rect 45950 46834 46002 46846
rect 53566 46898 53618 46910
rect 53566 46834 53618 46846
rect 2494 46786 2546 46798
rect 8878 46786 8930 46798
rect 5282 46734 5294 46786
rect 5346 46734 5358 46786
rect 2494 46722 2546 46734
rect 8878 46722 8930 46734
rect 12574 46786 12626 46798
rect 12574 46722 12626 46734
rect 12798 46786 12850 46798
rect 28590 46786 28642 46798
rect 23650 46734 23662 46786
rect 23714 46734 23726 46786
rect 12798 46722 12850 46734
rect 28590 46722 28642 46734
rect 28702 46786 28754 46798
rect 34750 46786 34802 46798
rect 29810 46734 29822 46786
rect 29874 46734 29886 46786
rect 31154 46734 31166 46786
rect 31218 46734 31230 46786
rect 28702 46722 28754 46734
rect 34750 46722 34802 46734
rect 35870 46786 35922 46798
rect 41022 46786 41074 46798
rect 37426 46734 37438 46786
rect 37490 46734 37502 46786
rect 39890 46734 39902 46786
rect 39954 46734 39966 46786
rect 35870 46722 35922 46734
rect 41022 46722 41074 46734
rect 41246 46786 41298 46798
rect 41246 46722 41298 46734
rect 46174 46786 46226 46798
rect 46174 46722 46226 46734
rect 48750 46786 48802 46798
rect 48750 46722 48802 46734
rect 8766 46674 8818 46686
rect 4162 46622 4174 46674
rect 4226 46622 4238 46674
rect 8766 46610 8818 46622
rect 9102 46674 9154 46686
rect 13470 46674 13522 46686
rect 28926 46674 28978 46686
rect 34974 46674 35026 46686
rect 11890 46622 11902 46674
rect 11954 46622 11966 46674
rect 13906 46622 13918 46674
rect 13970 46622 13982 46674
rect 14466 46622 14478 46674
rect 14530 46622 14542 46674
rect 14802 46622 14814 46674
rect 14866 46622 14878 46674
rect 17714 46622 17726 46674
rect 17778 46622 17790 46674
rect 19394 46622 19406 46674
rect 19458 46622 19470 46674
rect 23538 46622 23550 46674
rect 23602 46622 23614 46674
rect 24434 46622 24446 46674
rect 24498 46622 24510 46674
rect 26002 46622 26014 46674
rect 26066 46622 26078 46674
rect 27458 46622 27470 46674
rect 27522 46622 27534 46674
rect 32050 46622 32062 46674
rect 32114 46622 32126 46674
rect 9102 46610 9154 46622
rect 13470 46610 13522 46622
rect 28926 46610 28978 46622
rect 34974 46610 35026 46622
rect 35758 46674 35810 46686
rect 44494 46674 44546 46686
rect 45390 46674 45442 46686
rect 36642 46622 36654 46674
rect 36706 46622 36718 46674
rect 38882 46622 38894 46674
rect 38946 46622 38958 46674
rect 44818 46622 44830 46674
rect 44882 46622 44894 46674
rect 35758 46610 35810 46622
rect 44494 46610 44546 46622
rect 45390 46610 45442 46622
rect 45726 46674 45778 46686
rect 45726 46610 45778 46622
rect 47630 46674 47682 46686
rect 49310 46674 49362 46686
rect 50542 46674 50594 46686
rect 53678 46674 53730 46686
rect 48066 46622 48078 46674
rect 48130 46622 48142 46674
rect 49746 46622 49758 46674
rect 49810 46622 49822 46674
rect 53330 46622 53342 46674
rect 53394 46622 53406 46674
rect 47630 46610 47682 46622
rect 49310 46610 49362 46622
rect 50542 46610 50594 46622
rect 53678 46610 53730 46622
rect 54126 46674 54178 46686
rect 55010 46622 55022 46674
rect 55074 46622 55086 46674
rect 54126 46610 54178 46622
rect 2718 46562 2770 46574
rect 2718 46498 2770 46510
rect 3166 46562 3218 46574
rect 3166 46498 3218 46510
rect 3502 46562 3554 46574
rect 3502 46498 3554 46510
rect 5518 46562 5570 46574
rect 12686 46562 12738 46574
rect 26798 46562 26850 46574
rect 10098 46510 10110 46562
rect 10162 46510 10174 46562
rect 15922 46510 15934 46562
rect 15986 46510 15998 46562
rect 17938 46510 17950 46562
rect 18002 46510 18014 46562
rect 26226 46510 26238 46562
rect 26290 46510 26302 46562
rect 5518 46498 5570 46510
rect 12686 46498 12738 46510
rect 26798 46498 26850 46510
rect 29374 46562 29426 46574
rect 29374 46498 29426 46510
rect 31390 46562 31442 46574
rect 31390 46498 31442 46510
rect 31726 46562 31778 46574
rect 41694 46562 41746 46574
rect 37090 46510 37102 46562
rect 37154 46510 37166 46562
rect 31726 46498 31778 46510
rect 41694 46498 41746 46510
rect 45838 46562 45890 46574
rect 51102 46562 51154 46574
rect 50082 46510 50094 46562
rect 50146 46510 50158 46562
rect 45838 46498 45890 46510
rect 51102 46498 51154 46510
rect 53006 46562 53058 46574
rect 54898 46510 54910 46562
rect 54962 46510 54974 46562
rect 53006 46498 53058 46510
rect 32062 46450 32114 46462
rect 19730 46398 19742 46450
rect 19794 46398 19806 46450
rect 32062 46386 32114 46398
rect 36318 46450 36370 46462
rect 36318 46386 36370 46398
rect 40910 46450 40962 46462
rect 41458 46398 41470 46450
rect 41522 46447 41534 46450
rect 41794 46447 41806 46450
rect 41522 46401 41806 46447
rect 41522 46398 41534 46401
rect 41794 46398 41806 46401
rect 41858 46398 41870 46450
rect 40910 46386 40962 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 29262 46114 29314 46126
rect 9650 46062 9662 46114
rect 9714 46062 9726 46114
rect 18162 46062 18174 46114
rect 18226 46062 18238 46114
rect 27346 46062 27358 46114
rect 27410 46062 27422 46114
rect 29262 46050 29314 46062
rect 9102 46002 9154 46014
rect 14030 46002 14082 46014
rect 20190 46002 20242 46014
rect 37550 46002 37602 46014
rect 42142 46002 42194 46014
rect 9986 45950 9998 46002
rect 10050 45950 10062 46002
rect 12114 45950 12126 46002
rect 12178 45950 12190 46002
rect 17938 45950 17950 46002
rect 18002 45950 18014 46002
rect 29698 45950 29710 46002
rect 29762 45950 29774 46002
rect 31042 45950 31054 46002
rect 31106 45950 31118 46002
rect 39554 45950 39566 46002
rect 39618 45950 39630 46002
rect 41682 45950 41694 46002
rect 41746 45950 41758 46002
rect 9102 45938 9154 45950
rect 14030 45938 14082 45950
rect 20190 45938 20242 45950
rect 37550 45938 37602 45950
rect 42142 45938 42194 45950
rect 50654 46002 50706 46014
rect 50866 45950 50878 46002
rect 50930 45950 50942 46002
rect 55234 45950 55246 46002
rect 55298 45950 55310 46002
rect 50654 45938 50706 45950
rect 9326 45890 9378 45902
rect 15822 45890 15874 45902
rect 27246 45890 27298 45902
rect 45054 45890 45106 45902
rect 12786 45838 12798 45890
rect 12850 45838 12862 45890
rect 15026 45838 15038 45890
rect 15090 45838 15102 45890
rect 17042 45838 17054 45890
rect 17106 45838 17118 45890
rect 17826 45838 17838 45890
rect 17890 45838 17902 45890
rect 27906 45838 27918 45890
rect 27970 45838 27982 45890
rect 29026 45838 29038 45890
rect 29090 45838 29102 45890
rect 30146 45838 30158 45890
rect 30210 45838 30222 45890
rect 33954 45838 33966 45890
rect 34018 45838 34030 45890
rect 37986 45838 37998 45890
rect 38050 45838 38062 45890
rect 38882 45838 38894 45890
rect 38946 45838 38958 45890
rect 9326 45826 9378 45838
rect 15822 45826 15874 45838
rect 27246 45826 27298 45838
rect 45054 45826 45106 45838
rect 45278 45890 45330 45902
rect 45278 45826 45330 45838
rect 45502 45890 45554 45902
rect 45502 45826 45554 45838
rect 48414 45890 48466 45902
rect 49298 45838 49310 45890
rect 49362 45838 49374 45890
rect 58034 45838 58046 45890
rect 58098 45838 58110 45890
rect 48414 45826 48466 45838
rect 15486 45778 15538 45790
rect 49534 45778 49586 45790
rect 33170 45726 33182 45778
rect 33234 45726 33246 45778
rect 15486 45714 15538 45726
rect 49534 45714 49586 45726
rect 49982 45778 50034 45790
rect 49982 45714 50034 45726
rect 51214 45778 51266 45790
rect 57362 45726 57374 45778
rect 57426 45726 57438 45778
rect 51214 45714 51266 45726
rect 8094 45666 8146 45678
rect 8094 45602 8146 45614
rect 8206 45666 8258 45678
rect 8206 45602 8258 45614
rect 8318 45666 8370 45678
rect 8318 45602 8370 45614
rect 8542 45666 8594 45678
rect 8542 45602 8594 45614
rect 13582 45666 13634 45678
rect 15598 45666 15650 45678
rect 14802 45614 14814 45666
rect 14866 45614 14878 45666
rect 13582 45602 13634 45614
rect 15598 45602 15650 45614
rect 20750 45666 20802 45678
rect 20750 45602 20802 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 23102 45666 23154 45678
rect 23102 45602 23154 45614
rect 28590 45666 28642 45678
rect 28590 45602 28642 45614
rect 34414 45666 34466 45678
rect 34414 45602 34466 45614
rect 45390 45666 45442 45678
rect 45390 45602 45442 45614
rect 45950 45666 46002 45678
rect 50990 45666 51042 45678
rect 48066 45614 48078 45666
rect 48130 45614 48142 45666
rect 45950 45602 46002 45614
rect 50990 45602 51042 45614
rect 54910 45666 54962 45678
rect 54910 45602 54962 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 3054 45330 3106 45342
rect 3054 45266 3106 45278
rect 9662 45330 9714 45342
rect 9662 45266 9714 45278
rect 9774 45330 9826 45342
rect 9774 45266 9826 45278
rect 12462 45330 12514 45342
rect 22318 45330 22370 45342
rect 36654 45330 36706 45342
rect 14466 45278 14478 45330
rect 14530 45278 14542 45330
rect 23650 45278 23662 45330
rect 23714 45278 23726 45330
rect 24098 45278 24110 45330
rect 24162 45278 24174 45330
rect 28690 45278 28702 45330
rect 28754 45278 28766 45330
rect 12462 45266 12514 45278
rect 22318 45266 22370 45278
rect 36654 45266 36706 45278
rect 38446 45330 38498 45342
rect 38446 45266 38498 45278
rect 48302 45330 48354 45342
rect 48302 45266 48354 45278
rect 48750 45330 48802 45342
rect 48750 45266 48802 45278
rect 55918 45330 55970 45342
rect 55918 45266 55970 45278
rect 58158 45330 58210 45342
rect 58158 45266 58210 45278
rect 4958 45218 5010 45230
rect 21758 45218 21810 45230
rect 15362 45166 15374 45218
rect 15426 45166 15438 45218
rect 17490 45166 17502 45218
rect 17554 45166 17566 45218
rect 4958 45154 5010 45166
rect 21758 45154 21810 45166
rect 22206 45218 22258 45230
rect 55694 45218 55746 45230
rect 25218 45166 25230 45218
rect 25282 45166 25294 45218
rect 31826 45166 31838 45218
rect 31890 45166 31902 45218
rect 49074 45166 49086 45218
rect 49138 45166 49150 45218
rect 50754 45166 50766 45218
rect 50818 45166 50830 45218
rect 22206 45154 22258 45166
rect 55694 45154 55746 45166
rect 57150 45218 57202 45230
rect 57150 45154 57202 45166
rect 5070 45106 5122 45118
rect 9550 45106 9602 45118
rect 21646 45106 21698 45118
rect 6066 45054 6078 45106
rect 6130 45054 6142 45106
rect 10098 45054 10110 45106
rect 10162 45054 10174 45106
rect 14578 45054 14590 45106
rect 14642 45054 14654 45106
rect 15810 45054 15822 45106
rect 15874 45054 15886 45106
rect 18050 45054 18062 45106
rect 18114 45054 18126 45106
rect 18610 45054 18622 45106
rect 18674 45054 18686 45106
rect 5070 45042 5122 45054
rect 9550 45042 9602 45054
rect 21646 45042 21698 45054
rect 21982 45106 22034 45118
rect 21982 45042 22034 45054
rect 22430 45106 22482 45118
rect 22430 45042 22482 45054
rect 22878 45106 22930 45118
rect 22878 45042 22930 45054
rect 23326 45106 23378 45118
rect 43822 45106 43874 45118
rect 53342 45106 53394 45118
rect 25890 45054 25902 45106
rect 25954 45054 25966 45106
rect 26226 45054 26238 45106
rect 26290 45054 26302 45106
rect 28466 45054 28478 45106
rect 28530 45054 28542 45106
rect 31714 45054 31726 45106
rect 31778 45054 31790 45106
rect 32498 45054 32510 45106
rect 32562 45054 32574 45106
rect 36194 45054 36206 45106
rect 36258 45054 36270 45106
rect 49970 45054 49982 45106
rect 50034 45054 50046 45106
rect 23326 45042 23378 45054
rect 43822 45042 43874 45054
rect 53342 45042 53394 45054
rect 55470 45106 55522 45118
rect 55470 45042 55522 45054
rect 56030 45106 56082 45118
rect 56814 45106 56866 45118
rect 56578 45054 56590 45106
rect 56642 45054 56654 45106
rect 56030 45042 56082 45054
rect 56814 45042 56866 45054
rect 57038 45106 57090 45118
rect 57038 45042 57090 45054
rect 20974 44994 21026 45006
rect 6738 44942 6750 44994
rect 6802 44942 6814 44994
rect 8866 44942 8878 44994
rect 8930 44942 8942 44994
rect 15698 44942 15710 44994
rect 15762 44942 15774 44994
rect 17602 44942 17614 44994
rect 17666 44942 17678 44994
rect 20974 44930 21026 44942
rect 23102 44994 23154 45006
rect 23102 44930 23154 44942
rect 24670 44994 24722 45006
rect 24670 44930 24722 44942
rect 29150 44994 29202 45006
rect 55134 44994 55186 45006
rect 31938 44942 31950 44994
rect 32002 44942 32014 44994
rect 33282 44942 33294 44994
rect 33346 44942 33358 44994
rect 35410 44942 35422 44994
rect 35474 44942 35486 44994
rect 52882 44942 52894 44994
rect 52946 44942 52958 44994
rect 29150 44930 29202 44942
rect 55134 44930 55186 44942
rect 57598 44994 57650 45006
rect 57598 44930 57650 44942
rect 4958 44882 5010 44894
rect 4958 44818 5010 44830
rect 24446 44882 24498 44894
rect 24446 44818 24498 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 3502 44546 3554 44558
rect 3502 44482 3554 44494
rect 5966 44546 6018 44558
rect 5966 44482 6018 44494
rect 31726 44546 31778 44558
rect 54574 44546 54626 44558
rect 45378 44494 45390 44546
rect 45442 44494 45454 44546
rect 51202 44494 51214 44546
rect 51266 44494 51278 44546
rect 31726 44482 31778 44494
rect 54574 44482 54626 44494
rect 55246 44546 55298 44558
rect 56130 44494 56142 44546
rect 56194 44494 56206 44546
rect 57698 44494 57710 44546
rect 57762 44543 57774 44546
rect 58034 44543 58046 44546
rect 57762 44497 58046 44543
rect 57762 44494 57774 44497
rect 58034 44494 58046 44497
rect 58098 44494 58110 44546
rect 55246 44482 55298 44494
rect 5630 44434 5682 44446
rect 4162 44382 4174 44434
rect 4226 44382 4238 44434
rect 5630 44370 5682 44382
rect 7310 44434 7362 44446
rect 7310 44370 7362 44382
rect 8094 44434 8146 44446
rect 9550 44434 9602 44446
rect 35646 44434 35698 44446
rect 58270 44434 58322 44446
rect 8978 44382 8990 44434
rect 9042 44382 9054 44434
rect 16146 44382 16158 44434
rect 16210 44382 16222 44434
rect 19282 44382 19294 44434
rect 19346 44382 19358 44434
rect 43586 44382 43598 44434
rect 43650 44382 43662 44434
rect 45490 44382 45502 44434
rect 45554 44382 45566 44434
rect 51762 44382 51774 44434
rect 51826 44382 51838 44434
rect 54226 44382 54238 44434
rect 54290 44382 54302 44434
rect 8094 44370 8146 44382
rect 9550 44370 9602 44382
rect 35646 44370 35698 44382
rect 58270 44370 58322 44382
rect 6190 44322 6242 44334
rect 2482 44270 2494 44322
rect 2546 44270 2558 44322
rect 4498 44270 4510 44322
rect 4562 44270 4574 44322
rect 4946 44270 4958 44322
rect 5010 44270 5022 44322
rect 6190 44258 6242 44270
rect 7198 44322 7250 44334
rect 7198 44258 7250 44270
rect 7534 44322 7586 44334
rect 15150 44322 15202 44334
rect 23326 44322 23378 44334
rect 8754 44270 8766 44322
rect 8818 44270 8830 44322
rect 13682 44270 13694 44322
rect 13746 44270 13758 44322
rect 18722 44270 18734 44322
rect 18786 44270 18798 44322
rect 21746 44270 21758 44322
rect 21810 44270 21822 44322
rect 22082 44270 22094 44322
rect 22146 44270 22158 44322
rect 7534 44258 7586 44270
rect 15150 44258 15202 44270
rect 23326 44258 23378 44270
rect 24782 44322 24834 44334
rect 24782 44258 24834 44270
rect 31390 44322 31442 44334
rect 31390 44258 31442 44270
rect 32174 44322 32226 44334
rect 33630 44322 33682 44334
rect 32610 44270 32622 44322
rect 32674 44270 32686 44322
rect 32174 44258 32226 44270
rect 33630 44258 33682 44270
rect 34302 44322 34354 44334
rect 34302 44258 34354 44270
rect 34750 44322 34802 44334
rect 44270 44322 44322 44334
rect 46510 44322 46562 44334
rect 40786 44270 40798 44322
rect 40850 44270 40862 44322
rect 44706 44270 44718 44322
rect 44770 44270 44782 44322
rect 45602 44270 45614 44322
rect 45666 44270 45678 44322
rect 34750 44258 34802 44270
rect 44270 44258 44322 44270
rect 46510 44258 46562 44270
rect 46958 44322 47010 44334
rect 55470 44322 55522 44334
rect 51874 44270 51886 44322
rect 51938 44270 51950 44322
rect 46958 44258 47010 44270
rect 55470 44258 55522 44270
rect 56590 44322 56642 44334
rect 56914 44270 56926 44322
rect 56978 44270 56990 44322
rect 56590 44258 56642 44270
rect 2830 44210 2882 44222
rect 2830 44146 2882 44158
rect 3502 44210 3554 44222
rect 3502 44146 3554 44158
rect 3614 44210 3666 44222
rect 7758 44210 7810 44222
rect 15486 44210 15538 44222
rect 22318 44210 22370 44222
rect 3938 44158 3950 44210
rect 4002 44158 4014 44210
rect 13458 44158 13470 44210
rect 13522 44158 13534 44210
rect 17042 44158 17054 44210
rect 17106 44158 17118 44210
rect 3614 44146 3666 44158
rect 7758 44146 7810 44158
rect 15486 44146 15538 44158
rect 22318 44146 22370 44158
rect 22654 44210 22706 44222
rect 22654 44146 22706 44158
rect 24110 44210 24162 44222
rect 25566 44210 25618 44222
rect 24434 44158 24446 44210
rect 24498 44158 24510 44210
rect 24110 44146 24162 44158
rect 25566 44146 25618 44158
rect 25902 44210 25954 44222
rect 25902 44146 25954 44158
rect 31166 44210 31218 44222
rect 31166 44146 31218 44158
rect 33070 44210 33122 44222
rect 33070 44146 33122 44158
rect 34078 44210 34130 44222
rect 34078 44146 34130 44158
rect 35086 44210 35138 44222
rect 43934 44210 43986 44222
rect 41458 44158 41470 44210
rect 41522 44158 41534 44210
rect 35086 44146 35138 44158
rect 43934 44146 43986 44158
rect 44046 44210 44098 44222
rect 44046 44146 44098 44158
rect 46846 44210 46898 44222
rect 46846 44146 46898 44158
rect 56702 44210 56754 44222
rect 56702 44146 56754 44158
rect 57598 44210 57650 44222
rect 57598 44146 57650 44158
rect 2718 44098 2770 44110
rect 2718 44034 2770 44046
rect 15374 44098 15426 44110
rect 15374 44034 15426 44046
rect 22766 44098 22818 44110
rect 22766 44034 22818 44046
rect 22878 44098 22930 44110
rect 22878 44034 22930 44046
rect 23662 44098 23714 44110
rect 23662 44034 23714 44046
rect 33966 44098 34018 44110
rect 33966 44034 34018 44046
rect 34638 44098 34690 44110
rect 34638 44034 34690 44046
rect 34862 44098 34914 44110
rect 34862 44034 34914 44046
rect 37886 44098 37938 44110
rect 37886 44034 37938 44046
rect 46622 44098 46674 44110
rect 46622 44034 46674 44046
rect 54350 44098 54402 44110
rect 54898 44046 54910 44098
rect 54962 44046 54974 44098
rect 54350 44034 54402 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 4958 43762 5010 43774
rect 23214 43762 23266 43774
rect 14690 43710 14702 43762
rect 14754 43710 14766 43762
rect 32386 43710 32398 43762
rect 32450 43710 32462 43762
rect 37650 43710 37662 43762
rect 37714 43710 37726 43762
rect 4958 43698 5010 43710
rect 23214 43698 23266 43710
rect 5070 43650 5122 43662
rect 2482 43598 2494 43650
rect 2546 43598 2558 43650
rect 5070 43586 5122 43598
rect 5518 43650 5570 43662
rect 16382 43650 16434 43662
rect 22206 43650 22258 43662
rect 13906 43598 13918 43650
rect 13970 43598 13982 43650
rect 17714 43598 17726 43650
rect 17778 43598 17790 43650
rect 18386 43598 18398 43650
rect 18450 43598 18462 43650
rect 5518 43586 5570 43598
rect 16382 43586 16434 43598
rect 22206 43586 22258 43598
rect 22766 43650 22818 43662
rect 22766 43586 22818 43598
rect 29822 43650 29874 43662
rect 57374 43650 57426 43662
rect 36642 43598 36654 43650
rect 36706 43598 36718 43650
rect 38546 43598 38558 43650
rect 38610 43598 38622 43650
rect 46050 43598 46062 43650
rect 46114 43598 46126 43650
rect 29822 43586 29874 43598
rect 57374 43586 57426 43598
rect 57822 43650 57874 43662
rect 57822 43586 57874 43598
rect 17502 43538 17554 43550
rect 22542 43538 22594 43550
rect 1810 43486 1822 43538
rect 1874 43486 1886 43538
rect 13794 43486 13806 43538
rect 13858 43486 13870 43538
rect 14802 43486 14814 43538
rect 14866 43486 14878 43538
rect 15474 43486 15486 43538
rect 15538 43486 15550 43538
rect 19058 43486 19070 43538
rect 19122 43486 19134 43538
rect 17502 43474 17554 43486
rect 22542 43474 22594 43486
rect 29710 43538 29762 43550
rect 29710 43474 29762 43486
rect 29934 43538 29986 43550
rect 31838 43538 31890 43550
rect 30258 43486 30270 43538
rect 30322 43486 30334 43538
rect 29934 43474 29986 43486
rect 31838 43474 31890 43486
rect 32062 43538 32114 43550
rect 41022 43538 41074 43550
rect 52782 43538 52834 43550
rect 37090 43486 37102 43538
rect 37154 43486 37166 43538
rect 37762 43486 37774 43538
rect 37826 43486 37838 43538
rect 39666 43486 39678 43538
rect 39730 43486 39742 43538
rect 41458 43486 41470 43538
rect 41522 43486 41534 43538
rect 45266 43486 45278 43538
rect 45330 43486 45342 43538
rect 53218 43486 53230 43538
rect 53282 43486 53294 43538
rect 32062 43474 32114 43486
rect 41022 43474 41074 43486
rect 52782 43474 52834 43486
rect 17390 43426 17442 43438
rect 22318 43426 22370 43438
rect 40350 43426 40402 43438
rect 44942 43426 44994 43438
rect 4610 43374 4622 43426
rect 4674 43374 4686 43426
rect 16146 43374 16158 43426
rect 16210 43374 16222 43426
rect 19730 43374 19742 43426
rect 19794 43374 19806 43426
rect 21858 43374 21870 43426
rect 21922 43374 21934 43426
rect 38210 43374 38222 43426
rect 38274 43374 38286 43426
rect 42466 43374 42478 43426
rect 42530 43374 42542 43426
rect 48178 43374 48190 43426
rect 48242 43374 48254 43426
rect 54786 43374 54798 43426
rect 54850 43374 54862 43426
rect 57138 43374 57150 43426
rect 57202 43374 57214 43426
rect 17390 43362 17442 43374
rect 22318 43362 22370 43374
rect 40350 43362 40402 43374
rect 44942 43362 44994 43374
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 15934 42978 15986 42990
rect 10098 42926 10110 42978
rect 10162 42926 10174 42978
rect 15934 42914 15986 42926
rect 20190 42978 20242 42990
rect 20190 42914 20242 42926
rect 30942 42978 30994 42990
rect 30942 42914 30994 42926
rect 37102 42978 37154 42990
rect 37102 42914 37154 42926
rect 41358 42978 41410 42990
rect 41358 42914 41410 42926
rect 45614 42978 45666 42990
rect 45614 42914 45666 42926
rect 50094 42978 50146 42990
rect 50094 42914 50146 42926
rect 53566 42978 53618 42990
rect 53566 42914 53618 42926
rect 53678 42978 53730 42990
rect 53678 42914 53730 42926
rect 2942 42866 2994 42878
rect 8430 42866 8482 42878
rect 22094 42866 22146 42878
rect 31278 42866 31330 42878
rect 3714 42814 3726 42866
rect 3778 42814 3790 42866
rect 16370 42814 16382 42866
rect 16434 42814 16446 42866
rect 25330 42814 25342 42866
rect 25394 42814 25406 42866
rect 2942 42802 2994 42814
rect 8430 42802 8482 42814
rect 22094 42802 22146 42814
rect 31278 42802 31330 42814
rect 33518 42866 33570 42878
rect 33518 42802 33570 42814
rect 36430 42866 36482 42878
rect 36430 42802 36482 42814
rect 40238 42866 40290 42878
rect 46734 42866 46786 42878
rect 44146 42814 44158 42866
rect 44210 42814 44222 42866
rect 40238 42802 40290 42814
rect 46734 42802 46786 42814
rect 51662 42866 51714 42878
rect 57026 42814 57038 42866
rect 57090 42814 57102 42866
rect 51662 42802 51714 42814
rect 8878 42754 8930 42766
rect 27470 42754 27522 42766
rect 3602 42702 3614 42754
rect 3666 42702 3678 42754
rect 9650 42702 9662 42754
rect 9714 42702 9726 42754
rect 10098 42702 10110 42754
rect 10162 42702 10174 42754
rect 10546 42702 10558 42754
rect 10610 42702 10622 42754
rect 12562 42702 12574 42754
rect 12626 42702 12638 42754
rect 16482 42702 16494 42754
rect 16546 42702 16558 42754
rect 18162 42702 18174 42754
rect 18226 42702 18238 42754
rect 19618 42702 19630 42754
rect 19682 42702 19694 42754
rect 24770 42702 24782 42754
rect 24834 42702 24846 42754
rect 26002 42702 26014 42754
rect 26066 42702 26078 42754
rect 26226 42702 26238 42754
rect 26290 42702 26302 42754
rect 27122 42702 27134 42754
rect 27186 42702 27198 42754
rect 8878 42690 8930 42702
rect 27470 42690 27522 42702
rect 27694 42754 27746 42766
rect 27694 42690 27746 42702
rect 28366 42754 28418 42766
rect 39342 42754 39394 42766
rect 46622 42754 46674 42766
rect 53902 42754 53954 42766
rect 56478 42754 56530 42766
rect 29138 42702 29150 42754
rect 29202 42702 29214 42754
rect 30034 42702 30046 42754
rect 30098 42702 30110 42754
rect 30930 42702 30942 42754
rect 30994 42702 31006 42754
rect 37762 42702 37774 42754
rect 37826 42702 37838 42754
rect 38098 42702 38110 42754
rect 38162 42702 38174 42754
rect 39778 42702 39790 42754
rect 39842 42702 39854 42754
rect 40786 42702 40798 42754
rect 40850 42702 40862 42754
rect 51538 42702 51550 42754
rect 51602 42702 51614 42754
rect 51762 42702 51774 42754
rect 51826 42702 51838 42754
rect 55906 42702 55918 42754
rect 55970 42702 55982 42754
rect 28366 42690 28418 42702
rect 39342 42690 39394 42702
rect 46622 42690 46674 42702
rect 53902 42690 53954 42702
rect 56478 42690 56530 42702
rect 8766 42642 8818 42654
rect 15598 42642 15650 42654
rect 20302 42642 20354 42654
rect 14130 42590 14142 42642
rect 14194 42590 14206 42642
rect 16818 42590 16830 42642
rect 16882 42590 16894 42642
rect 8766 42578 8818 42590
rect 15598 42578 15650 42590
rect 20302 42578 20354 42590
rect 20750 42642 20802 42654
rect 20750 42578 20802 42590
rect 21310 42642 21362 42654
rect 21310 42578 21362 42590
rect 21646 42642 21698 42654
rect 37214 42642 37266 42654
rect 40574 42642 40626 42654
rect 24994 42590 25006 42642
rect 25058 42590 25070 42642
rect 30594 42590 30606 42642
rect 30658 42590 30670 42642
rect 38546 42590 38558 42642
rect 38610 42590 38622 42642
rect 21646 42578 21698 42590
rect 37214 42578 37266 42590
rect 40574 42578 40626 42590
rect 41694 42642 41746 42654
rect 41694 42578 41746 42590
rect 42030 42642 42082 42654
rect 45614 42642 45666 42654
rect 42242 42590 42254 42642
rect 42306 42590 42318 42642
rect 43922 42590 43934 42642
rect 43986 42590 43998 42642
rect 42030 42578 42082 42590
rect 45614 42578 45666 42590
rect 45726 42642 45778 42654
rect 45726 42578 45778 42590
rect 50206 42642 50258 42654
rect 50206 42578 50258 42590
rect 54014 42642 54066 42654
rect 54014 42578 54066 42590
rect 55470 42642 55522 42654
rect 55470 42578 55522 42590
rect 56926 42642 56978 42654
rect 56926 42578 56978 42590
rect 8990 42530 9042 42542
rect 8990 42466 9042 42478
rect 12350 42530 12402 42542
rect 12350 42466 12402 42478
rect 13806 42530 13858 42542
rect 13806 42466 13858 42478
rect 15822 42530 15874 42542
rect 15822 42466 15874 42478
rect 20526 42530 20578 42542
rect 20526 42466 20578 42478
rect 28478 42530 28530 42542
rect 28478 42466 28530 42478
rect 28702 42530 28754 42542
rect 33182 42530 33234 42542
rect 29250 42478 29262 42530
rect 29314 42478 29326 42530
rect 29474 42478 29486 42530
rect 29538 42478 29550 42530
rect 28702 42466 28754 42478
rect 33182 42466 33234 42478
rect 34078 42530 34130 42542
rect 34078 42466 34130 42478
rect 37102 42530 37154 42542
rect 41470 42530 41522 42542
rect 37650 42478 37662 42530
rect 37714 42478 37726 42530
rect 37102 42466 37154 42478
rect 41470 42466 41522 42478
rect 45166 42530 45218 42542
rect 45166 42466 45218 42478
rect 46398 42530 46450 42542
rect 46398 42466 46450 42478
rect 46846 42530 46898 42542
rect 46846 42466 46898 42478
rect 49646 42530 49698 42542
rect 49646 42466 49698 42478
rect 50094 42530 50146 42542
rect 50094 42466 50146 42478
rect 51998 42530 52050 42542
rect 51998 42466 52050 42478
rect 53118 42530 53170 42542
rect 53118 42466 53170 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 9662 42194 9714 42206
rect 9662 42130 9714 42142
rect 28030 42194 28082 42206
rect 28030 42130 28082 42142
rect 28478 42194 28530 42206
rect 28478 42130 28530 42142
rect 32622 42194 32674 42206
rect 32622 42130 32674 42142
rect 33630 42194 33682 42206
rect 33630 42130 33682 42142
rect 15038 42082 15090 42094
rect 23662 42082 23714 42094
rect 11554 42030 11566 42082
rect 11618 42030 11630 42082
rect 13570 42030 13582 42082
rect 13634 42030 13646 42082
rect 15586 42030 15598 42082
rect 15650 42030 15662 42082
rect 19506 42030 19518 42082
rect 19570 42030 19582 42082
rect 21186 42030 21198 42082
rect 21250 42030 21262 42082
rect 21634 42030 21646 42082
rect 21698 42030 21710 42082
rect 15038 42018 15090 42030
rect 23662 42018 23714 42030
rect 23774 42082 23826 42094
rect 34078 42082 34130 42094
rect 27234 42030 27246 42082
rect 27298 42030 27310 42082
rect 23774 42018 23826 42030
rect 34078 42018 34130 42030
rect 35534 42082 35586 42094
rect 57038 42082 57090 42094
rect 53778 42030 53790 42082
rect 53842 42030 53854 42082
rect 35534 42018 35586 42030
rect 57038 42018 57090 42030
rect 9550 41970 9602 41982
rect 5394 41918 5406 41970
rect 5458 41918 5470 41970
rect 8978 41918 8990 41970
rect 9042 41918 9054 41970
rect 9550 41906 9602 41918
rect 9886 41970 9938 41982
rect 14702 41970 14754 41982
rect 11666 41918 11678 41970
rect 11730 41918 11742 41970
rect 12786 41918 12798 41970
rect 12850 41918 12862 41970
rect 9886 41906 9938 41918
rect 14702 41906 14754 41918
rect 15374 41970 15426 41982
rect 26910 41970 26962 41982
rect 16034 41918 16046 41970
rect 16098 41918 16110 41970
rect 16706 41918 16718 41970
rect 16770 41918 16782 41970
rect 18274 41918 18286 41970
rect 18338 41918 18350 41970
rect 18722 41918 18734 41970
rect 18786 41918 18798 41970
rect 20402 41918 20414 41970
rect 20466 41918 20478 41970
rect 20738 41918 20750 41970
rect 20802 41918 20814 41970
rect 21522 41918 21534 41970
rect 21586 41918 21598 41970
rect 25106 41918 25118 41970
rect 25170 41918 25182 41970
rect 25890 41918 25902 41970
rect 25954 41918 25966 41970
rect 15374 41906 15426 41918
rect 26910 41906 26962 41918
rect 27918 41970 27970 41982
rect 28590 41970 28642 41982
rect 28130 41918 28142 41970
rect 28194 41918 28206 41970
rect 27918 41906 27970 41918
rect 28590 41906 28642 41918
rect 28702 41970 28754 41982
rect 29486 41970 29538 41982
rect 30382 41970 30434 41982
rect 41134 41970 41186 41982
rect 29026 41918 29038 41970
rect 29090 41918 29102 41970
rect 29698 41918 29710 41970
rect 29762 41918 29774 41970
rect 35858 41918 35870 41970
rect 35922 41918 35934 41970
rect 36866 41918 36878 41970
rect 36930 41918 36942 41970
rect 38770 41918 38782 41970
rect 38834 41918 38846 41970
rect 28702 41906 28754 41918
rect 29486 41906 29538 41918
rect 30382 41906 30434 41918
rect 41134 41906 41186 41918
rect 41358 41970 41410 41982
rect 52446 41970 52498 41982
rect 57374 41970 57426 41982
rect 41682 41918 41694 41970
rect 41746 41918 41758 41970
rect 43810 41918 43822 41970
rect 43874 41918 43886 41970
rect 49186 41918 49198 41970
rect 49250 41918 49262 41970
rect 53106 41918 53118 41970
rect 53170 41918 53182 41970
rect 41358 41906 41410 41918
rect 52446 41906 52498 41918
rect 57374 41906 57426 41918
rect 57710 41970 57762 41982
rect 57710 41906 57762 41918
rect 58158 41970 58210 41982
rect 58158 41906 58210 41918
rect 3278 41858 3330 41870
rect 8766 41858 8818 41870
rect 6066 41806 6078 41858
rect 6130 41806 6142 41858
rect 8194 41806 8206 41858
rect 8258 41806 8270 41858
rect 3278 41794 3330 41806
rect 8766 41794 8818 41806
rect 10334 41858 10386 41870
rect 22542 41858 22594 41870
rect 14578 41806 14590 41858
rect 14642 41806 14654 41858
rect 19954 41806 19966 41858
rect 20018 41806 20030 41858
rect 10334 41794 10386 41806
rect 22542 41794 22594 41806
rect 22878 41858 22930 41870
rect 40350 41858 40402 41870
rect 25778 41806 25790 41858
rect 25842 41806 25854 41858
rect 33730 41806 33742 41858
rect 33794 41806 33806 41858
rect 34402 41806 34414 41858
rect 34466 41806 34478 41858
rect 37202 41806 37214 41858
rect 37266 41806 37278 41858
rect 38098 41806 38110 41858
rect 38162 41806 38174 41858
rect 38882 41806 38894 41858
rect 38946 41806 38958 41858
rect 22878 41794 22930 41806
rect 40350 41794 40402 41806
rect 41246 41858 41298 41870
rect 41246 41794 41298 41806
rect 42142 41858 42194 41870
rect 42142 41794 42194 41806
rect 43486 41858 43538 41870
rect 43486 41794 43538 41806
rect 44494 41858 44546 41870
rect 56702 41858 56754 41870
rect 49858 41806 49870 41858
rect 49922 41806 49934 41858
rect 51986 41806 51998 41858
rect 52050 41806 52062 41858
rect 55906 41806 55918 41858
rect 55970 41806 55982 41858
rect 44494 41794 44546 41806
rect 56702 41794 56754 41806
rect 57486 41858 57538 41870
rect 57486 41794 57538 41806
rect 8654 41746 8706 41758
rect 8654 41682 8706 41694
rect 15262 41746 15314 41758
rect 23662 41746 23714 41758
rect 22530 41694 22542 41746
rect 22594 41743 22606 41746
rect 22866 41743 22878 41746
rect 22594 41697 22878 41743
rect 22594 41694 22606 41697
rect 22866 41694 22878 41697
rect 22930 41694 22942 41746
rect 15262 41682 15314 41694
rect 23662 41682 23714 41694
rect 25678 41746 25730 41758
rect 25678 41682 25730 41694
rect 27694 41746 27746 41758
rect 27694 41682 27746 41694
rect 33406 41746 33458 41758
rect 43822 41746 43874 41758
rect 34626 41694 34638 41746
rect 34690 41694 34702 41746
rect 38994 41694 39006 41746
rect 39058 41694 39070 41746
rect 33406 41682 33458 41694
rect 43822 41682 43874 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 44158 41410 44210 41422
rect 27122 41358 27134 41410
rect 27186 41358 27198 41410
rect 32274 41358 32286 41410
rect 32338 41358 32350 41410
rect 44158 41346 44210 41358
rect 45166 41410 45218 41422
rect 45166 41346 45218 41358
rect 50318 41410 50370 41422
rect 50318 41346 50370 41358
rect 52894 41410 52946 41422
rect 52894 41346 52946 41358
rect 21310 41298 21362 41310
rect 2706 41246 2718 41298
rect 2770 41246 2782 41298
rect 4162 41246 4174 41298
rect 4226 41246 4238 41298
rect 21310 41234 21362 41246
rect 22318 41298 22370 41310
rect 23774 41298 23826 41310
rect 33630 41298 33682 41310
rect 23314 41246 23326 41298
rect 23378 41246 23390 41298
rect 24882 41246 24894 41298
rect 24946 41246 24958 41298
rect 27458 41246 27470 41298
rect 27522 41246 27534 41298
rect 32498 41246 32510 41298
rect 32562 41246 32574 41298
rect 22318 41234 22370 41246
rect 23774 41234 23826 41246
rect 33630 41234 33682 41246
rect 34862 41298 34914 41310
rect 34862 41234 34914 41246
rect 36990 41298 37042 41310
rect 36990 41234 37042 41246
rect 38558 41298 38610 41310
rect 43486 41298 43538 41310
rect 52670 41298 52722 41310
rect 40114 41246 40126 41298
rect 40178 41246 40190 41298
rect 45490 41246 45502 41298
rect 45554 41246 45566 41298
rect 50530 41246 50542 41298
rect 50594 41246 50606 41298
rect 38558 41234 38610 41246
rect 43486 41234 43538 41246
rect 52670 41234 52722 41246
rect 5518 41186 5570 41198
rect 20526 41186 20578 41198
rect 4050 41134 4062 41186
rect 4114 41134 4126 41186
rect 5170 41134 5182 41186
rect 5234 41134 5246 41186
rect 8530 41134 8542 41186
rect 8594 41134 8606 41186
rect 9538 41134 9550 41186
rect 9602 41134 9614 41186
rect 15138 41134 15150 41186
rect 15202 41134 15214 41186
rect 15698 41134 15710 41186
rect 15762 41134 15774 41186
rect 17826 41134 17838 41186
rect 17890 41134 17902 41186
rect 19506 41134 19518 41186
rect 19570 41134 19582 41186
rect 5518 41122 5570 41134
rect 20526 41122 20578 41134
rect 21870 41186 21922 41198
rect 21870 41122 21922 41134
rect 23438 41186 23490 41198
rect 25566 41186 25618 41198
rect 25106 41134 25118 41186
rect 25170 41134 25182 41186
rect 23438 41122 23490 41134
rect 25566 41122 25618 41134
rect 25902 41186 25954 41198
rect 25902 41122 25954 41134
rect 28030 41186 28082 41198
rect 28030 41122 28082 41134
rect 29038 41186 29090 41198
rect 34638 41186 34690 41198
rect 32050 41134 32062 41186
rect 32114 41134 32126 41186
rect 33170 41134 33182 41186
rect 33234 41134 33246 41186
rect 33954 41134 33966 41186
rect 34018 41134 34030 41186
rect 29038 41122 29090 41134
rect 34638 41122 34690 41134
rect 34750 41186 34802 41198
rect 34750 41122 34802 41134
rect 35534 41186 35586 41198
rect 35534 41122 35586 41134
rect 35758 41186 35810 41198
rect 37102 41186 37154 41198
rect 51886 41186 51938 41198
rect 36082 41134 36094 41186
rect 36146 41134 36158 41186
rect 37426 41134 37438 41186
rect 37490 41134 37502 41186
rect 43026 41134 43038 41186
rect 43090 41134 43102 41186
rect 35758 41122 35810 41134
rect 37102 41122 37154 41134
rect 51886 41122 51938 41134
rect 51998 41186 52050 41198
rect 51998 41122 52050 41134
rect 53118 41186 53170 41198
rect 55682 41134 55694 41186
rect 55746 41134 55758 41186
rect 57586 41134 57598 41186
rect 57650 41134 57662 41186
rect 53118 41122 53170 41134
rect 2830 41074 2882 41086
rect 2830 41010 2882 41022
rect 3054 41074 3106 41086
rect 5854 41074 5906 41086
rect 12686 41074 12738 41086
rect 19966 41074 20018 41086
rect 3714 41022 3726 41074
rect 3778 41022 3790 41074
rect 9650 41022 9662 41074
rect 9714 41022 9726 41074
rect 16370 41022 16382 41074
rect 16434 41022 16446 41074
rect 17154 41022 17166 41074
rect 17218 41022 17230 41074
rect 18722 41022 18734 41074
rect 18786 41022 18798 41074
rect 3054 41010 3106 41022
rect 5854 41010 5906 41022
rect 12686 41010 12738 41022
rect 19966 41010 20018 41022
rect 20190 41074 20242 41086
rect 20190 41010 20242 41022
rect 26462 41074 26514 41086
rect 26462 41010 26514 41022
rect 26574 41074 26626 41086
rect 26574 41010 26626 41022
rect 26686 41074 26738 41086
rect 26686 41010 26738 41022
rect 29374 41074 29426 41086
rect 44270 41074 44322 41086
rect 42242 41022 42254 41074
rect 42306 41022 42318 41074
rect 29374 41010 29426 41022
rect 44270 41010 44322 41022
rect 51550 41074 51602 41086
rect 55346 41022 55358 41074
rect 55410 41022 55422 41074
rect 57250 41022 57262 41074
rect 57314 41022 57326 41074
rect 51550 41010 51602 41022
rect 5742 40962 5794 40974
rect 12350 40962 12402 40974
rect 8306 40910 8318 40962
rect 8370 40910 8382 40962
rect 5742 40898 5794 40910
rect 12350 40898 12402 40910
rect 14590 40962 14642 40974
rect 14590 40898 14642 40910
rect 20302 40962 20354 40974
rect 20302 40898 20354 40910
rect 27470 40962 27522 40974
rect 27470 40898 27522 40910
rect 27694 40962 27746 40974
rect 27694 40898 27746 40910
rect 29262 40962 29314 40974
rect 29262 40898 29314 40910
rect 34078 40962 34130 40974
rect 34078 40898 34130 40910
rect 34974 40962 35026 40974
rect 34974 40898 35026 40910
rect 35086 40962 35138 40974
rect 35086 40898 35138 40910
rect 44158 40962 44210 40974
rect 44158 40898 44210 40910
rect 45390 40962 45442 40974
rect 45390 40898 45442 40910
rect 50542 40962 50594 40974
rect 50542 40898 50594 40910
rect 51662 40962 51714 40974
rect 51662 40898 51714 40910
rect 53566 40962 53618 40974
rect 56018 40910 56030 40962
rect 56082 40910 56094 40962
rect 53566 40898 53618 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 5070 40626 5122 40638
rect 12238 40626 12290 40638
rect 8082 40574 8094 40626
rect 8146 40574 8158 40626
rect 5070 40562 5122 40574
rect 12238 40562 12290 40574
rect 13582 40626 13634 40638
rect 13582 40562 13634 40574
rect 14590 40626 14642 40638
rect 14590 40562 14642 40574
rect 19742 40626 19794 40638
rect 19742 40562 19794 40574
rect 22542 40626 22594 40638
rect 22542 40562 22594 40574
rect 24334 40626 24386 40638
rect 24334 40562 24386 40574
rect 41134 40626 41186 40638
rect 41134 40562 41186 40574
rect 55694 40626 55746 40638
rect 55694 40562 55746 40574
rect 58158 40626 58210 40638
rect 58158 40562 58210 40574
rect 6190 40514 6242 40526
rect 2482 40462 2494 40514
rect 2546 40462 2558 40514
rect 6190 40450 6242 40462
rect 6526 40514 6578 40526
rect 6526 40450 6578 40462
rect 12462 40514 12514 40526
rect 12462 40450 12514 40462
rect 13358 40514 13410 40526
rect 13358 40450 13410 40462
rect 14366 40514 14418 40526
rect 17950 40514 18002 40526
rect 16706 40462 16718 40514
rect 16770 40462 16782 40514
rect 14366 40450 14418 40462
rect 17950 40450 18002 40462
rect 21198 40514 21250 40526
rect 21198 40450 21250 40462
rect 21310 40514 21362 40526
rect 21310 40450 21362 40462
rect 24110 40514 24162 40526
rect 38782 40514 38834 40526
rect 34850 40462 34862 40514
rect 34914 40462 34926 40514
rect 35634 40462 35646 40514
rect 35698 40462 35710 40514
rect 24110 40450 24162 40462
rect 38782 40450 38834 40462
rect 40238 40514 40290 40526
rect 40238 40450 40290 40462
rect 40350 40514 40402 40526
rect 55918 40514 55970 40526
rect 43474 40462 43486 40514
rect 43538 40462 43550 40514
rect 45938 40462 45950 40514
rect 46002 40462 46014 40514
rect 56690 40462 56702 40514
rect 56754 40462 56766 40514
rect 40350 40450 40402 40462
rect 55918 40450 55970 40462
rect 12574 40402 12626 40414
rect 14254 40402 14306 40414
rect 1810 40350 1822 40402
rect 1874 40350 1886 40402
rect 7858 40350 7870 40402
rect 7922 40350 7934 40402
rect 13794 40350 13806 40402
rect 13858 40350 13870 40402
rect 12574 40338 12626 40350
rect 14254 40338 14306 40350
rect 14814 40402 14866 40414
rect 15710 40402 15762 40414
rect 15138 40350 15150 40402
rect 15202 40350 15214 40402
rect 14814 40338 14866 40350
rect 15710 40338 15762 40350
rect 17502 40402 17554 40414
rect 17502 40338 17554 40350
rect 20302 40402 20354 40414
rect 20302 40338 20354 40350
rect 20862 40402 20914 40414
rect 20862 40338 20914 40350
rect 21870 40402 21922 40414
rect 21870 40338 21922 40350
rect 22990 40402 23042 40414
rect 22990 40338 23042 40350
rect 23774 40402 23826 40414
rect 28926 40402 28978 40414
rect 27122 40350 27134 40402
rect 27186 40350 27198 40402
rect 27794 40350 27806 40402
rect 27858 40350 27870 40402
rect 23774 40338 23826 40350
rect 28926 40338 28978 40350
rect 29262 40402 29314 40414
rect 40798 40402 40850 40414
rect 31378 40350 31390 40402
rect 31442 40350 31454 40402
rect 34514 40350 34526 40402
rect 34578 40350 34590 40402
rect 35746 40350 35758 40402
rect 35810 40350 35822 40402
rect 37986 40350 37998 40402
rect 38050 40350 38062 40402
rect 29262 40338 29314 40350
rect 40798 40338 40850 40350
rect 41246 40402 41298 40414
rect 41246 40338 41298 40350
rect 41358 40402 41410 40414
rect 48750 40402 48802 40414
rect 43810 40350 43822 40402
rect 43874 40350 43886 40402
rect 44706 40350 44718 40402
rect 44770 40350 44782 40402
rect 45154 40350 45166 40402
rect 45218 40350 45230 40402
rect 41358 40338 41410 40350
rect 48750 40338 48802 40350
rect 49310 40402 49362 40414
rect 56030 40402 56082 40414
rect 51650 40350 51662 40402
rect 51714 40350 51726 40402
rect 57026 40350 57038 40402
rect 57090 40350 57102 40402
rect 57474 40350 57486 40402
rect 57538 40350 57550 40402
rect 49310 40338 49362 40350
rect 56030 40338 56082 40350
rect 8542 40290 8594 40302
rect 4610 40238 4622 40290
rect 4674 40238 4686 40290
rect 8542 40226 8594 40238
rect 13694 40290 13746 40302
rect 13694 40226 13746 40238
rect 15374 40290 15426 40302
rect 15374 40226 15426 40238
rect 19182 40290 19234 40302
rect 24446 40290 24498 40302
rect 29374 40290 29426 40302
rect 22642 40238 22654 40290
rect 22706 40238 22718 40290
rect 23426 40238 23438 40290
rect 23490 40238 23502 40290
rect 27570 40238 27582 40290
rect 27634 40238 27646 40290
rect 28018 40238 28030 40290
rect 28082 40238 28094 40290
rect 19182 40226 19234 40238
rect 24446 40226 24498 40238
rect 29374 40226 29426 40238
rect 31166 40290 31218 40302
rect 43710 40290 43762 40302
rect 50990 40290 51042 40302
rect 35858 40238 35870 40290
rect 35922 40238 35934 40290
rect 38098 40238 38110 40290
rect 38162 40238 38174 40290
rect 48066 40238 48078 40290
rect 48130 40238 48142 40290
rect 51762 40238 51774 40290
rect 51826 40238 51838 40290
rect 56914 40238 56926 40290
rect 56978 40238 56990 40290
rect 31166 40226 31218 40238
rect 43710 40226 43762 40238
rect 50990 40226 51042 40238
rect 21310 40178 21362 40190
rect 16594 40126 16606 40178
rect 16658 40126 16670 40178
rect 21310 40114 21362 40126
rect 22318 40178 22370 40190
rect 22318 40114 22370 40126
rect 40238 40178 40290 40190
rect 40238 40114 40290 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 5630 39842 5682 39854
rect 5630 39778 5682 39790
rect 5966 39842 6018 39854
rect 45838 39842 45890 39854
rect 26002 39790 26014 39842
rect 26066 39790 26078 39842
rect 5966 39778 6018 39790
rect 45838 39778 45890 39790
rect 47406 39842 47458 39854
rect 47406 39778 47458 39790
rect 51326 39842 51378 39854
rect 51326 39778 51378 39790
rect 57486 39842 57538 39854
rect 57486 39778 57538 39790
rect 57822 39842 57874 39854
rect 57822 39778 57874 39790
rect 6862 39730 6914 39742
rect 17726 39730 17778 39742
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 12786 39678 12798 39730
rect 12850 39678 12862 39730
rect 14578 39678 14590 39730
rect 14642 39678 14654 39730
rect 14802 39678 14814 39730
rect 14866 39678 14878 39730
rect 6862 39666 6914 39678
rect 17726 39666 17778 39678
rect 17838 39730 17890 39742
rect 17838 39666 17890 39678
rect 22654 39730 22706 39742
rect 22654 39666 22706 39678
rect 23774 39730 23826 39742
rect 32174 39730 32226 39742
rect 26114 39678 26126 39730
rect 26178 39678 26190 39730
rect 27906 39678 27918 39730
rect 27970 39678 27982 39730
rect 23774 39666 23826 39678
rect 32174 39666 32226 39678
rect 32510 39730 32562 39742
rect 47518 39730 47570 39742
rect 35186 39678 35198 39730
rect 35250 39678 35262 39730
rect 45266 39678 45278 39730
rect 45330 39678 45342 39730
rect 32510 39666 32562 39678
rect 47518 39666 47570 39678
rect 50654 39730 50706 39742
rect 50978 39678 50990 39730
rect 51042 39678 51054 39730
rect 56466 39678 56478 39730
rect 56530 39678 56542 39730
rect 50654 39666 50706 39678
rect 18734 39618 18786 39630
rect 31278 39618 31330 39630
rect 34638 39618 34690 39630
rect 3154 39566 3166 39618
rect 3218 39566 3230 39618
rect 11442 39566 11454 39618
rect 11506 39566 11518 39618
rect 12338 39566 12350 39618
rect 12402 39566 12414 39618
rect 14130 39566 14142 39618
rect 14194 39566 14206 39618
rect 14914 39566 14926 39618
rect 14978 39566 14990 39618
rect 15922 39566 15934 39618
rect 15986 39566 15998 39618
rect 20178 39566 20190 39618
rect 20242 39566 20254 39618
rect 22194 39566 22206 39618
rect 22258 39566 22270 39618
rect 25554 39566 25566 39618
rect 25618 39566 25630 39618
rect 26226 39566 26238 39618
rect 26290 39566 26302 39618
rect 26450 39566 26462 39618
rect 26514 39566 26526 39618
rect 31490 39566 31502 39618
rect 31554 39566 31566 39618
rect 18734 39554 18786 39566
rect 31278 39554 31330 39566
rect 34638 39554 34690 39566
rect 34862 39618 34914 39630
rect 34862 39554 34914 39566
rect 41694 39618 41746 39630
rect 41694 39554 41746 39566
rect 43374 39618 43426 39630
rect 43810 39566 43822 39618
rect 43874 39566 43886 39618
rect 45378 39566 45390 39618
rect 45442 39566 45454 39618
rect 49186 39566 49198 39618
rect 49250 39566 49262 39618
rect 53666 39566 53678 39618
rect 53730 39566 53742 39618
rect 57026 39566 57038 39618
rect 57090 39566 57102 39618
rect 43374 39554 43426 39566
rect 5742 39506 5794 39518
rect 16494 39506 16546 39518
rect 21310 39506 21362 39518
rect 4274 39454 4286 39506
rect 4338 39454 4350 39506
rect 12786 39454 12798 39506
rect 12850 39454 12862 39506
rect 13794 39454 13806 39506
rect 13858 39454 13870 39506
rect 20402 39454 20414 39506
rect 20466 39454 20478 39506
rect 5742 39442 5794 39454
rect 16494 39442 16546 39454
rect 21310 39442 21362 39454
rect 21646 39506 21698 39518
rect 21646 39442 21698 39454
rect 25006 39506 25058 39518
rect 25006 39442 25058 39454
rect 44270 39506 44322 39518
rect 44270 39442 44322 39454
rect 45054 39506 45106 39518
rect 45054 39442 45106 39454
rect 45726 39506 45778 39518
rect 45726 39442 45778 39454
rect 51102 39506 51154 39518
rect 57598 39506 57650 39518
rect 54338 39454 54350 39506
rect 54402 39454 54414 39506
rect 56802 39454 56814 39506
rect 56866 39454 56878 39506
rect 51102 39442 51154 39454
rect 57598 39442 57650 39454
rect 13470 39394 13522 39406
rect 2818 39342 2830 39394
rect 2882 39342 2894 39394
rect 11554 39342 11566 39394
rect 11618 39342 11630 39394
rect 13470 39330 13522 39342
rect 23998 39394 24050 39406
rect 23998 39330 24050 39342
rect 27470 39394 27522 39406
rect 27470 39330 27522 39342
rect 33070 39394 33122 39406
rect 33070 39330 33122 39342
rect 42254 39394 42306 39406
rect 42254 39330 42306 39342
rect 45838 39394 45890 39406
rect 45838 39330 45890 39342
rect 48974 39394 49026 39406
rect 48974 39330 49026 39342
rect 49758 39394 49810 39406
rect 49758 39330 49810 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 6190 39058 6242 39070
rect 6190 38994 6242 39006
rect 8206 39058 8258 39070
rect 8206 38994 8258 39006
rect 8542 39058 8594 39070
rect 19630 39058 19682 39070
rect 13122 39006 13134 39058
rect 13186 39006 13198 39058
rect 18834 39006 18846 39058
rect 18898 39006 18910 39058
rect 8542 38994 8594 39006
rect 19630 38994 19682 39006
rect 27694 39058 27746 39070
rect 27694 38994 27746 39006
rect 27918 39058 27970 39070
rect 27918 38994 27970 39006
rect 44830 39058 44882 39070
rect 44830 38994 44882 39006
rect 48862 39058 48914 39070
rect 48862 38994 48914 39006
rect 53566 39058 53618 39070
rect 53566 38994 53618 39006
rect 54126 39058 54178 39070
rect 54126 38994 54178 39006
rect 7982 38946 8034 38958
rect 7982 38882 8034 38894
rect 12126 38946 12178 38958
rect 12126 38882 12178 38894
rect 12350 38946 12402 38958
rect 12350 38882 12402 38894
rect 17838 38946 17890 38958
rect 17838 38882 17890 38894
rect 20526 38946 20578 38958
rect 20526 38882 20578 38894
rect 30382 38946 30434 38958
rect 30382 38882 30434 38894
rect 37550 38946 37602 38958
rect 37550 38882 37602 38894
rect 37886 38946 37938 38958
rect 39442 38894 39454 38946
rect 39506 38894 39518 38946
rect 50978 38894 50990 38946
rect 51042 38894 51054 38946
rect 57810 38894 57822 38946
rect 57874 38894 57886 38946
rect 37886 38882 37938 38894
rect 6414 38834 6466 38846
rect 6414 38770 6466 38782
rect 6638 38834 6690 38846
rect 7870 38834 7922 38846
rect 7074 38782 7086 38834
rect 7138 38782 7150 38834
rect 6638 38770 6690 38782
rect 7870 38770 7922 38782
rect 11342 38834 11394 38846
rect 11342 38770 11394 38782
rect 12462 38834 12514 38846
rect 12462 38770 12514 38782
rect 12686 38834 12738 38846
rect 20974 38834 21026 38846
rect 15698 38782 15710 38834
rect 15762 38782 15774 38834
rect 16034 38782 16046 38834
rect 16098 38782 16110 38834
rect 12686 38770 12738 38782
rect 20974 38770 21026 38782
rect 21310 38834 21362 38846
rect 21310 38770 21362 38782
rect 23438 38834 23490 38846
rect 23438 38770 23490 38782
rect 23662 38834 23714 38846
rect 23662 38770 23714 38782
rect 24110 38834 24162 38846
rect 28030 38834 28082 38846
rect 25666 38782 25678 38834
rect 25730 38782 25742 38834
rect 27010 38782 27022 38834
rect 27074 38782 27086 38834
rect 27234 38782 27246 38834
rect 27298 38782 27310 38834
rect 24110 38770 24162 38782
rect 28030 38770 28082 38782
rect 30046 38834 30098 38846
rect 30046 38770 30098 38782
rect 30606 38834 30658 38846
rect 30606 38770 30658 38782
rect 32510 38834 32562 38846
rect 58158 38834 58210 38846
rect 34066 38782 34078 38834
rect 34130 38782 34142 38834
rect 34738 38782 34750 38834
rect 34802 38782 34814 38834
rect 39666 38782 39678 38834
rect 39730 38782 39742 38834
rect 40002 38782 40014 38834
rect 40066 38782 40078 38834
rect 50306 38782 50318 38834
rect 50370 38782 50382 38834
rect 32510 38770 32562 38782
rect 58158 38770 58210 38782
rect 6526 38722 6578 38734
rect 11566 38722 11618 38734
rect 22654 38722 22706 38734
rect 29934 38722 29986 38734
rect 39230 38722 39282 38734
rect 7410 38670 7422 38722
rect 7474 38670 7486 38722
rect 15810 38670 15822 38722
rect 15874 38670 15886 38722
rect 23874 38670 23886 38722
rect 23938 38670 23950 38722
rect 25554 38670 25566 38722
rect 25618 38670 25630 38722
rect 26898 38670 26910 38722
rect 26962 38670 26974 38722
rect 32162 38670 32174 38722
rect 32226 38670 32238 38722
rect 34290 38670 34302 38722
rect 34354 38670 34366 38722
rect 34962 38670 34974 38722
rect 35026 38670 35038 38722
rect 6526 38658 6578 38670
rect 11566 38658 11618 38670
rect 22654 38658 22706 38670
rect 29934 38658 29986 38670
rect 39230 38658 39282 38670
rect 45950 38722 46002 38734
rect 45950 38658 46002 38670
rect 46174 38722 46226 38734
rect 46174 38658 46226 38670
rect 49422 38722 49474 38734
rect 53902 38722 53954 38734
rect 56702 38722 56754 38734
rect 53106 38670 53118 38722
rect 53170 38670 53182 38722
rect 54226 38670 54238 38722
rect 54290 38670 54302 38722
rect 49422 38658 49474 38670
rect 53902 38658 53954 38670
rect 56702 38658 56754 38670
rect 57598 38722 57650 38734
rect 57598 38658 57650 38670
rect 24222 38610 24274 38622
rect 30270 38610 30322 38622
rect 10994 38558 11006 38610
rect 11058 38558 11070 38610
rect 15362 38558 15374 38610
rect 15426 38558 15438 38610
rect 26562 38558 26574 38610
rect 26626 38558 26638 38610
rect 24222 38546 24274 38558
rect 30270 38546 30322 38558
rect 30830 38610 30882 38622
rect 31938 38558 31950 38610
rect 32002 38558 32014 38610
rect 46498 38558 46510 38610
rect 46562 38558 46574 38610
rect 30830 38546 30882 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 3950 38274 4002 38286
rect 3950 38210 4002 38222
rect 9774 38274 9826 38286
rect 9774 38210 9826 38222
rect 11790 38274 11842 38286
rect 12574 38274 12626 38286
rect 12226 38222 12238 38274
rect 12290 38222 12302 38274
rect 11790 38210 11842 38222
rect 12574 38210 12626 38222
rect 13694 38274 13746 38286
rect 13694 38210 13746 38222
rect 24558 38274 24610 38286
rect 24558 38210 24610 38222
rect 26014 38274 26066 38286
rect 26014 38210 26066 38222
rect 29262 38274 29314 38286
rect 29262 38210 29314 38222
rect 30494 38274 30546 38286
rect 30494 38210 30546 38222
rect 4510 38162 4562 38174
rect 7758 38162 7810 38174
rect 6850 38110 6862 38162
rect 6914 38110 6926 38162
rect 4510 38098 4562 38110
rect 7758 38098 7810 38110
rect 12798 38162 12850 38174
rect 17950 38162 18002 38174
rect 16594 38110 16606 38162
rect 16658 38110 16670 38162
rect 12798 38098 12850 38110
rect 17950 38098 18002 38110
rect 19742 38162 19794 38174
rect 19742 38098 19794 38110
rect 21198 38162 21250 38174
rect 36318 38162 36370 38174
rect 27010 38110 27022 38162
rect 27074 38110 27086 38162
rect 27570 38110 27582 38162
rect 27634 38110 27646 38162
rect 28130 38110 28142 38162
rect 28194 38110 28206 38162
rect 21198 38098 21250 38110
rect 36318 38098 36370 38110
rect 38334 38162 38386 38174
rect 58146 38166 58158 38218
rect 58210 38166 58222 38218
rect 38770 38110 38782 38162
rect 38834 38110 38846 38162
rect 46386 38110 46398 38162
rect 46450 38110 46462 38162
rect 38334 38098 38386 38110
rect 4062 38050 4114 38062
rect 4062 37986 4114 37998
rect 5854 38050 5906 38062
rect 5854 37986 5906 37998
rect 6190 38050 6242 38062
rect 6190 37986 6242 37998
rect 6414 38050 6466 38062
rect 9438 38050 9490 38062
rect 7186 37998 7198 38050
rect 7250 37998 7262 38050
rect 8754 37998 8766 38050
rect 8818 37998 8830 38050
rect 6414 37986 6466 37998
rect 9438 37986 9490 37998
rect 11454 38050 11506 38062
rect 11454 37986 11506 37998
rect 14030 38050 14082 38062
rect 17614 38050 17666 38062
rect 21310 38050 21362 38062
rect 24222 38050 24274 38062
rect 14802 37998 14814 38050
rect 14866 37998 14878 38050
rect 17042 37998 17054 38050
rect 17106 37998 17118 38050
rect 20178 37998 20190 38050
rect 20242 37998 20254 38050
rect 22978 37998 22990 38050
rect 23042 37998 23054 38050
rect 14030 37986 14082 37998
rect 17614 37986 17666 37998
rect 21310 37986 21362 37998
rect 24222 37986 24274 37998
rect 26126 38050 26178 38062
rect 35310 38050 35362 38062
rect 27122 37998 27134 38050
rect 27186 37998 27198 38050
rect 27458 37998 27470 38050
rect 27522 37998 27534 38050
rect 28578 37998 28590 38050
rect 28642 37998 28654 38050
rect 31266 37998 31278 38050
rect 31330 37998 31342 38050
rect 32946 37998 32958 38050
rect 33010 37998 33022 38050
rect 34402 37998 34414 38050
rect 34466 37998 34478 38050
rect 26126 37986 26178 37998
rect 35310 37986 35362 37998
rect 36542 38050 36594 38062
rect 41582 38050 41634 38062
rect 37090 37998 37102 38050
rect 37154 37998 37166 38050
rect 40226 37998 40238 38050
rect 40290 37998 40302 38050
rect 36542 37986 36594 37998
rect 41582 37986 41634 37998
rect 42142 38050 42194 38062
rect 42142 37986 42194 37998
rect 45390 38050 45442 38062
rect 45390 37986 45442 37998
rect 45838 38050 45890 38062
rect 54910 38050 54962 38062
rect 49298 37998 49310 38050
rect 49362 37998 49374 38050
rect 55346 37998 55358 38050
rect 55410 37998 55422 38050
rect 45838 37986 45890 37998
rect 54910 37986 54962 37998
rect 23998 37938 24050 37950
rect 8642 37886 8654 37938
rect 8706 37886 8718 37938
rect 10658 37886 10670 37938
rect 10722 37886 10734 37938
rect 11218 37886 11230 37938
rect 11282 37886 11294 37938
rect 14690 37886 14702 37938
rect 14754 37886 14766 37938
rect 21522 37886 21534 37938
rect 21586 37886 21598 37938
rect 22082 37886 22094 37938
rect 22146 37886 22158 37938
rect 22754 37886 22766 37938
rect 22818 37886 22830 37938
rect 23998 37874 24050 37886
rect 28142 37938 28194 37950
rect 28142 37874 28194 37886
rect 29262 37938 29314 37950
rect 29262 37874 29314 37886
rect 29374 37938 29426 37950
rect 29374 37874 29426 37886
rect 30606 37938 30658 37950
rect 35646 37938 35698 37950
rect 31826 37886 31838 37938
rect 31890 37886 31902 37938
rect 35074 37886 35086 37938
rect 35138 37886 35150 37938
rect 30606 37874 30658 37886
rect 35646 37874 35698 37886
rect 35982 37938 36034 37950
rect 46062 37938 46114 37950
rect 37314 37886 37326 37938
rect 37378 37886 37390 37938
rect 37650 37886 37662 37938
rect 37714 37886 37726 37938
rect 38994 37886 39006 37938
rect 39058 37886 39070 37938
rect 48514 37886 48526 37938
rect 48578 37886 48590 37938
rect 56018 37886 56030 37938
rect 56082 37886 56094 37938
rect 35982 37874 36034 37886
rect 46062 37874 46114 37886
rect 3950 37826 4002 37838
rect 3950 37762 4002 37774
rect 5966 37826 6018 37838
rect 5966 37762 6018 37774
rect 16158 37826 16210 37838
rect 16158 37762 16210 37774
rect 26014 37826 26066 37838
rect 26014 37762 26066 37774
rect 28366 37826 28418 37838
rect 28366 37762 28418 37774
rect 30494 37826 30546 37838
rect 35534 37826 35586 37838
rect 34850 37774 34862 37826
rect 34914 37774 34926 37826
rect 30494 37762 30546 37774
rect 35534 37762 35586 37774
rect 36206 37826 36258 37838
rect 45278 37826 45330 37838
rect 40786 37774 40798 37826
rect 40850 37774 40862 37826
rect 36206 37762 36258 37774
rect 45278 37762 45330 37774
rect 45950 37826 46002 37838
rect 45950 37762 46002 37774
rect 49758 37826 49810 37838
rect 49758 37762 49810 37774
rect 53566 37826 53618 37838
rect 53566 37762 53618 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 3614 37490 3666 37502
rect 3614 37426 3666 37438
rect 7870 37490 7922 37502
rect 7870 37426 7922 37438
rect 8990 37490 9042 37502
rect 14142 37490 14194 37502
rect 12562 37438 12574 37490
rect 12626 37438 12638 37490
rect 8990 37426 9042 37438
rect 14142 37426 14194 37438
rect 17502 37490 17554 37502
rect 17502 37426 17554 37438
rect 24558 37490 24610 37502
rect 24558 37426 24610 37438
rect 25342 37490 25394 37502
rect 39006 37490 39058 37502
rect 30706 37438 30718 37490
rect 30770 37438 30782 37490
rect 37090 37438 37102 37490
rect 37154 37438 37166 37490
rect 25342 37426 25394 37438
rect 39006 37426 39058 37438
rect 39902 37490 39954 37502
rect 39902 37426 39954 37438
rect 44270 37490 44322 37502
rect 44270 37426 44322 37438
rect 46510 37490 46562 37502
rect 46510 37426 46562 37438
rect 46622 37490 46674 37502
rect 46622 37426 46674 37438
rect 2718 37378 2770 37390
rect 2718 37314 2770 37326
rect 3054 37378 3106 37390
rect 8654 37378 8706 37390
rect 5282 37326 5294 37378
rect 5346 37326 5358 37378
rect 8418 37326 8430 37378
rect 8482 37326 8494 37378
rect 3054 37314 3106 37326
rect 8654 37314 8706 37326
rect 8766 37378 8818 37390
rect 8766 37314 8818 37326
rect 11342 37378 11394 37390
rect 14366 37378 14418 37390
rect 12226 37326 12238 37378
rect 12290 37326 12302 37378
rect 12450 37326 12462 37378
rect 12514 37326 12526 37378
rect 11342 37314 11394 37326
rect 14366 37314 14418 37326
rect 14478 37378 14530 37390
rect 14478 37314 14530 37326
rect 14814 37378 14866 37390
rect 23662 37378 23714 37390
rect 16818 37326 16830 37378
rect 16882 37326 16894 37378
rect 14814 37314 14866 37326
rect 23662 37314 23714 37326
rect 26014 37378 26066 37390
rect 26014 37314 26066 37326
rect 26126 37378 26178 37390
rect 35758 37378 35810 37390
rect 39566 37378 39618 37390
rect 26786 37326 26798 37378
rect 26850 37326 26862 37378
rect 37202 37326 37214 37378
rect 37266 37326 37278 37378
rect 37762 37326 37774 37378
rect 37826 37326 37838 37378
rect 26126 37314 26178 37326
rect 35758 37314 35810 37326
rect 39566 37314 39618 37326
rect 39678 37378 39730 37390
rect 39678 37314 39730 37326
rect 46398 37378 46450 37390
rect 46398 37314 46450 37326
rect 3166 37266 3218 37278
rect 3166 37202 3218 37214
rect 3726 37266 3778 37278
rect 3726 37202 3778 37214
rect 3838 37266 3890 37278
rect 3838 37202 3890 37214
rect 4286 37266 4338 37278
rect 9438 37266 9490 37278
rect 4610 37214 4622 37266
rect 4674 37214 4686 37266
rect 4286 37202 4338 37214
rect 9438 37202 9490 37214
rect 10222 37266 10274 37278
rect 14926 37266 14978 37278
rect 24558 37266 24610 37278
rect 27134 37266 27186 37278
rect 31278 37266 31330 37278
rect 33630 37266 33682 37278
rect 37102 37266 37154 37278
rect 11890 37214 11902 37266
rect 11954 37214 11966 37266
rect 15362 37214 15374 37266
rect 15426 37214 15438 37266
rect 15922 37214 15934 37266
rect 15986 37214 15998 37266
rect 16482 37214 16494 37266
rect 16546 37214 16558 37266
rect 18834 37214 18846 37266
rect 18898 37214 18910 37266
rect 20290 37214 20302 37266
rect 20354 37214 20366 37266
rect 21410 37214 21422 37266
rect 21474 37214 21486 37266
rect 26562 37214 26574 37266
rect 26626 37214 26638 37266
rect 27570 37214 27582 37266
rect 27634 37214 27646 37266
rect 29138 37214 29150 37266
rect 29202 37214 29214 37266
rect 33394 37214 33406 37266
rect 33458 37214 33470 37266
rect 36642 37214 36654 37266
rect 36706 37214 36718 37266
rect 39218 37214 39230 37266
rect 39282 37214 39294 37266
rect 43810 37214 43822 37266
rect 43874 37214 43886 37266
rect 10222 37202 10274 37214
rect 14926 37202 14978 37214
rect 24558 37202 24610 37214
rect 27134 37202 27186 37214
rect 31278 37202 31330 37214
rect 33630 37202 33682 37214
rect 37102 37202 37154 37214
rect 2830 37154 2882 37166
rect 8878 37154 8930 37166
rect 22878 37154 22930 37166
rect 7410 37102 7422 37154
rect 7474 37102 7486 37154
rect 16706 37102 16718 37154
rect 16770 37102 16782 37154
rect 20402 37102 20414 37154
rect 20466 37102 20478 37154
rect 21186 37102 21198 37154
rect 21250 37102 21262 37154
rect 2830 37090 2882 37102
rect 8878 37090 8930 37102
rect 22878 37090 22930 37102
rect 25230 37154 25282 37166
rect 34066 37102 34078 37154
rect 34130 37102 34142 37154
rect 40898 37102 40910 37154
rect 40962 37102 40974 37154
rect 43026 37102 43038 37154
rect 43090 37102 43102 37154
rect 25230 37090 25282 37102
rect 9662 37042 9714 37054
rect 15150 37042 15202 37054
rect 31054 37042 31106 37054
rect 11106 36990 11118 37042
rect 11170 36990 11182 37042
rect 20626 36990 20638 37042
rect 20690 36990 20702 37042
rect 27234 36990 27246 37042
rect 27298 36990 27310 37042
rect 9662 36978 9714 36990
rect 15150 36978 15202 36990
rect 31054 36978 31106 36990
rect 38894 37042 38946 37054
rect 38894 36978 38946 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 23102 36706 23154 36718
rect 23102 36642 23154 36654
rect 24558 36706 24610 36718
rect 35646 36706 35698 36718
rect 27346 36654 27358 36706
rect 27410 36654 27422 36706
rect 24558 36642 24610 36654
rect 35646 36642 35698 36654
rect 36878 36706 36930 36718
rect 36878 36642 36930 36654
rect 40910 36706 40962 36718
rect 40910 36642 40962 36654
rect 41246 36706 41298 36718
rect 41246 36642 41298 36654
rect 5182 36594 5234 36606
rect 16270 36594 16322 36606
rect 2482 36542 2494 36594
rect 2546 36542 2558 36594
rect 4610 36542 4622 36594
rect 4674 36542 4686 36594
rect 9314 36542 9326 36594
rect 9378 36542 9390 36594
rect 11890 36542 11902 36594
rect 11954 36542 11966 36594
rect 15810 36542 15822 36594
rect 15874 36542 15886 36594
rect 5182 36530 5234 36542
rect 16270 36530 16322 36542
rect 17278 36594 17330 36606
rect 17278 36530 17330 36542
rect 22542 36594 22594 36606
rect 22542 36530 22594 36542
rect 24110 36594 24162 36606
rect 28366 36594 28418 36606
rect 33294 36594 33346 36606
rect 37886 36594 37938 36606
rect 52894 36594 52946 36606
rect 56702 36594 56754 36606
rect 27010 36542 27022 36594
rect 27074 36542 27086 36594
rect 30706 36542 30718 36594
rect 30770 36542 30782 36594
rect 35522 36542 35534 36594
rect 35586 36542 35598 36594
rect 52098 36542 52110 36594
rect 52162 36542 52174 36594
rect 56130 36542 56142 36594
rect 56194 36542 56206 36594
rect 24110 36530 24162 36542
rect 28366 36530 28418 36542
rect 33294 36530 33346 36542
rect 37886 36530 37938 36542
rect 52894 36530 52946 36542
rect 56702 36530 56754 36542
rect 8542 36482 8594 36494
rect 13470 36482 13522 36494
rect 22766 36482 22818 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 11442 36430 11454 36482
rect 11506 36430 11518 36482
rect 12786 36430 12798 36482
rect 12850 36430 12862 36482
rect 15698 36430 15710 36482
rect 15762 36430 15774 36482
rect 16818 36430 16830 36482
rect 16882 36430 16894 36482
rect 17714 36430 17726 36482
rect 17778 36430 17790 36482
rect 18274 36430 18286 36482
rect 18338 36430 18350 36482
rect 18834 36430 18846 36482
rect 18898 36430 18910 36482
rect 19394 36430 19406 36482
rect 19458 36430 19470 36482
rect 8542 36418 8594 36430
rect 13470 36418 13522 36430
rect 22766 36418 22818 36430
rect 23662 36482 23714 36494
rect 23662 36418 23714 36430
rect 23998 36482 24050 36494
rect 23998 36418 24050 36430
rect 24334 36482 24386 36494
rect 24334 36418 24386 36430
rect 24670 36482 24722 36494
rect 37102 36482 37154 36494
rect 26898 36430 26910 36482
rect 26962 36430 26974 36482
rect 33058 36430 33070 36482
rect 33122 36430 33134 36482
rect 35410 36430 35422 36482
rect 35474 36430 35486 36482
rect 36194 36430 36206 36482
rect 36258 36430 36270 36482
rect 24670 36418 24722 36430
rect 37102 36418 37154 36430
rect 37662 36482 37714 36494
rect 49298 36430 49310 36482
rect 49362 36430 49374 36482
rect 53330 36430 53342 36482
rect 53394 36430 53406 36482
rect 37662 36418 37714 36430
rect 8878 36370 8930 36382
rect 8878 36306 8930 36318
rect 11118 36370 11170 36382
rect 19630 36370 19682 36382
rect 11554 36318 11566 36370
rect 11618 36318 11630 36370
rect 17602 36318 17614 36370
rect 17666 36318 17678 36370
rect 11118 36306 11170 36318
rect 19630 36306 19682 36318
rect 32062 36370 32114 36382
rect 44046 36370 44098 36382
rect 37426 36318 37438 36370
rect 37490 36318 37502 36370
rect 49970 36318 49982 36370
rect 50034 36318 50046 36370
rect 54002 36318 54014 36370
rect 54066 36318 54078 36370
rect 32062 36306 32114 36318
rect 44046 36306 44098 36318
rect 8766 36258 8818 36270
rect 8766 36194 8818 36206
rect 9774 36258 9826 36270
rect 9774 36194 9826 36206
rect 10782 36258 10834 36270
rect 10782 36194 10834 36206
rect 11006 36258 11058 36270
rect 11006 36194 11058 36206
rect 12686 36258 12738 36270
rect 12686 36194 12738 36206
rect 13582 36258 13634 36270
rect 13582 36194 13634 36206
rect 13806 36258 13858 36270
rect 13806 36194 13858 36206
rect 20750 36258 20802 36270
rect 20750 36194 20802 36206
rect 21310 36258 21362 36270
rect 27806 36258 27858 36270
rect 21634 36206 21646 36258
rect 21698 36206 21710 36258
rect 21310 36194 21362 36206
rect 27806 36194 27858 36206
rect 31166 36258 31218 36270
rect 31166 36194 31218 36206
rect 32958 36258 33010 36270
rect 32958 36194 33010 36206
rect 41134 36258 41186 36270
rect 41134 36194 41186 36206
rect 41694 36258 41746 36270
rect 41694 36194 41746 36206
rect 43822 36258 43874 36270
rect 43822 36194 43874 36206
rect 43934 36258 43986 36270
rect 43934 36194 43986 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 11678 35922 11730 35934
rect 11678 35858 11730 35870
rect 12910 35922 12962 35934
rect 12910 35858 12962 35870
rect 23326 35922 23378 35934
rect 27246 35922 27298 35934
rect 24210 35870 24222 35922
rect 24274 35870 24286 35922
rect 23326 35858 23378 35870
rect 27246 35858 27298 35870
rect 28366 35922 28418 35934
rect 37326 35922 37378 35934
rect 31378 35870 31390 35922
rect 31442 35870 31454 35922
rect 28366 35858 28418 35870
rect 37326 35858 37378 35870
rect 38334 35922 38386 35934
rect 38334 35858 38386 35870
rect 38782 35922 38834 35934
rect 38782 35858 38834 35870
rect 39006 35922 39058 35934
rect 39006 35858 39058 35870
rect 50430 35922 50482 35934
rect 51214 35922 51266 35934
rect 50978 35919 50990 35922
rect 50430 35858 50482 35870
rect 50769 35873 50990 35919
rect 2270 35810 2322 35822
rect 2270 35746 2322 35758
rect 10334 35810 10386 35822
rect 10334 35746 10386 35758
rect 12798 35810 12850 35822
rect 27358 35810 27410 35822
rect 32398 35810 32450 35822
rect 15026 35758 15038 35810
rect 15090 35758 15102 35810
rect 18834 35758 18846 35810
rect 18898 35758 18910 35810
rect 30930 35758 30942 35810
rect 30994 35758 31006 35810
rect 12798 35746 12850 35758
rect 27358 35746 27410 35758
rect 32398 35746 32450 35758
rect 34974 35810 35026 35822
rect 34974 35746 35026 35758
rect 36318 35810 36370 35822
rect 36318 35746 36370 35758
rect 37438 35810 37490 35822
rect 50769 35810 50815 35873
rect 50978 35870 50990 35873
rect 51042 35870 51054 35922
rect 51214 35858 51266 35870
rect 55134 35922 55186 35934
rect 55134 35858 55186 35870
rect 56814 35922 56866 35934
rect 56814 35858 56866 35870
rect 57710 35922 57762 35934
rect 57710 35858 57762 35870
rect 44818 35758 44830 35810
rect 44882 35758 44894 35810
rect 50754 35758 50766 35810
rect 50818 35758 50830 35810
rect 37438 35746 37490 35758
rect 11342 35698 11394 35710
rect 1810 35646 1822 35698
rect 1874 35646 1886 35698
rect 10098 35646 10110 35698
rect 10162 35646 10174 35698
rect 11342 35634 11394 35646
rect 11678 35698 11730 35710
rect 11678 35634 11730 35646
rect 12014 35698 12066 35710
rect 32510 35698 32562 35710
rect 36654 35698 36706 35710
rect 37998 35698 38050 35710
rect 12338 35646 12350 35698
rect 12402 35646 12414 35698
rect 12562 35646 12574 35698
rect 12626 35646 12638 35698
rect 13906 35646 13918 35698
rect 13970 35646 13982 35698
rect 15810 35646 15822 35698
rect 15874 35646 15886 35698
rect 18498 35646 18510 35698
rect 18562 35646 18574 35698
rect 20290 35646 20302 35698
rect 20354 35646 20366 35698
rect 21074 35646 21086 35698
rect 21138 35646 21150 35698
rect 23986 35646 23998 35698
rect 24050 35646 24062 35698
rect 25330 35646 25342 35698
rect 25394 35646 25406 35698
rect 30482 35646 30494 35698
rect 30546 35646 30558 35698
rect 31378 35646 31390 35698
rect 31442 35646 31454 35698
rect 35970 35646 35982 35698
rect 36034 35646 36046 35698
rect 36418 35646 36430 35698
rect 36482 35646 36494 35698
rect 37650 35646 37662 35698
rect 37714 35646 37726 35698
rect 12014 35634 12066 35646
rect 32510 35634 32562 35646
rect 36654 35634 36706 35646
rect 37998 35634 38050 35646
rect 39118 35698 39170 35710
rect 39118 35634 39170 35646
rect 42478 35698 42530 35710
rect 52894 35698 52946 35710
rect 45490 35646 45502 35698
rect 45554 35646 45566 35698
rect 50642 35646 50654 35698
rect 50706 35646 50718 35698
rect 52098 35646 52110 35698
rect 52162 35646 52174 35698
rect 42478 35634 42530 35646
rect 52894 35634 52946 35646
rect 54910 35698 54962 35710
rect 54910 35634 54962 35646
rect 55358 35698 55410 35710
rect 55358 35634 55410 35646
rect 55582 35698 55634 35710
rect 55582 35634 55634 35646
rect 56590 35698 56642 35710
rect 56590 35634 56642 35646
rect 57038 35698 57090 35710
rect 57038 35634 57090 35646
rect 57150 35698 57202 35710
rect 57150 35634 57202 35646
rect 57598 35698 57650 35710
rect 57598 35634 57650 35646
rect 57934 35698 57986 35710
rect 57934 35634 57986 35646
rect 33630 35586 33682 35598
rect 13570 35534 13582 35586
rect 13634 35534 13646 35586
rect 16034 35534 16046 35586
rect 16098 35534 16110 35586
rect 18610 35534 18622 35586
rect 18674 35534 18686 35586
rect 22866 35534 22878 35586
rect 22930 35534 22942 35586
rect 25666 35534 25678 35586
rect 25730 35534 25742 35586
rect 33630 35522 33682 35534
rect 34190 35586 34242 35598
rect 34190 35522 34242 35534
rect 38222 35586 38274 35598
rect 42690 35534 42702 35586
rect 42754 35534 42766 35586
rect 51986 35534 51998 35586
rect 52050 35534 52062 35586
rect 38222 35522 38274 35534
rect 21646 35474 21698 35486
rect 21646 35410 21698 35422
rect 32398 35474 32450 35486
rect 32398 35410 32450 35422
rect 50318 35474 50370 35486
rect 50318 35410 50370 35422
rect 51774 35474 51826 35486
rect 51774 35410 51826 35422
rect 53118 35474 53170 35486
rect 53118 35410 53170 35422
rect 53454 35474 53506 35486
rect 53454 35410 53506 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 37550 35138 37602 35150
rect 10658 35086 10670 35138
rect 10722 35086 10734 35138
rect 37550 35074 37602 35086
rect 38110 35138 38162 35150
rect 38110 35074 38162 35086
rect 44942 35138 44994 35150
rect 44942 35074 44994 35086
rect 1822 35026 1874 35038
rect 17054 35026 17106 35038
rect 10322 34974 10334 35026
rect 10386 34974 10398 35026
rect 1822 34962 1874 34974
rect 17054 34962 17106 34974
rect 20078 35026 20130 35038
rect 28366 35026 28418 35038
rect 24210 34974 24222 35026
rect 24274 34974 24286 35026
rect 20078 34962 20130 34974
rect 28366 34962 28418 34974
rect 29710 35026 29762 35038
rect 29710 34962 29762 34974
rect 35758 35026 35810 35038
rect 40798 35026 40850 35038
rect 37874 34974 37886 35026
rect 37938 34974 37950 35026
rect 35758 34962 35810 34974
rect 40798 34962 40850 34974
rect 44046 35026 44098 35038
rect 44046 34962 44098 34974
rect 45502 35026 45554 35038
rect 49982 35026 50034 35038
rect 46050 34974 46062 35026
rect 46114 34974 46126 35026
rect 45502 34962 45554 34974
rect 49982 34962 50034 34974
rect 15374 34914 15426 34926
rect 43934 34914 43986 34926
rect 55470 34914 55522 34926
rect 7298 34862 7310 34914
rect 7362 34862 7374 34914
rect 7970 34862 7982 34914
rect 8034 34862 8046 34914
rect 9874 34862 9886 34914
rect 9938 34862 9950 34914
rect 10546 34862 10558 34914
rect 10610 34862 10622 34914
rect 12786 34862 12798 34914
rect 12850 34862 12862 34914
rect 21298 34862 21310 34914
rect 21362 34862 21374 34914
rect 27906 34862 27918 34914
rect 27970 34862 27982 34914
rect 30258 34862 30270 34914
rect 30322 34862 30334 34914
rect 36194 34862 36206 34914
rect 36258 34862 36270 34914
rect 48850 34862 48862 34914
rect 48914 34862 48926 34914
rect 53218 34862 53230 34914
rect 53282 34862 53294 34914
rect 15374 34850 15426 34862
rect 43934 34850 43986 34862
rect 55470 34850 55522 34862
rect 56590 34914 56642 34926
rect 56590 34850 56642 34862
rect 12574 34802 12626 34814
rect 7522 34750 7534 34802
rect 7586 34750 7598 34802
rect 12574 34738 12626 34750
rect 16270 34802 16322 34814
rect 16270 34738 16322 34750
rect 20862 34802 20914 34814
rect 29822 34802 29874 34814
rect 36990 34802 37042 34814
rect 22082 34750 22094 34802
rect 22146 34750 22158 34802
rect 34962 34750 34974 34802
rect 35026 34750 35038 34802
rect 20862 34738 20914 34750
rect 29822 34738 29874 34750
rect 36990 34738 37042 34750
rect 43598 34802 43650 34814
rect 43598 34738 43650 34750
rect 44158 34802 44210 34814
rect 44158 34738 44210 34750
rect 44942 34802 44994 34814
rect 44942 34738 44994 34750
rect 45054 34802 45106 34814
rect 49422 34802 49474 34814
rect 48178 34750 48190 34802
rect 48242 34750 48254 34802
rect 45054 34738 45106 34750
rect 49422 34738 49474 34750
rect 49534 34802 49586 34814
rect 49534 34738 49586 34750
rect 55806 34802 55858 34814
rect 55806 34738 55858 34750
rect 56254 34802 56306 34814
rect 56254 34738 56306 34750
rect 56366 34802 56418 34814
rect 56366 34738 56418 34750
rect 56926 34802 56978 34814
rect 56926 34738 56978 34750
rect 57038 34802 57090 34814
rect 57038 34738 57090 34750
rect 16718 34690 16770 34702
rect 8082 34638 8094 34690
rect 8146 34638 8158 34690
rect 16718 34626 16770 34638
rect 19518 34690 19570 34702
rect 19518 34626 19570 34638
rect 27582 34690 27634 34702
rect 27582 34626 27634 34638
rect 29374 34690 29426 34702
rect 29374 34626 29426 34638
rect 29598 34690 29650 34702
rect 29598 34626 29650 34638
rect 37214 34690 37266 34702
rect 37214 34626 37266 34638
rect 37438 34690 37490 34702
rect 37438 34626 37490 34638
rect 37886 34690 37938 34702
rect 37886 34626 37938 34638
rect 38670 34690 38722 34702
rect 38670 34626 38722 34638
rect 39342 34690 39394 34702
rect 55694 34690 55746 34702
rect 53442 34638 53454 34690
rect 53506 34638 53518 34690
rect 39342 34626 39394 34638
rect 55694 34626 55746 34638
rect 56702 34690 56754 34702
rect 56702 34626 56754 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 7870 34354 7922 34366
rect 7870 34290 7922 34302
rect 8094 34354 8146 34366
rect 8094 34290 8146 34302
rect 9662 34354 9714 34366
rect 9662 34290 9714 34302
rect 15150 34354 15202 34366
rect 29150 34354 29202 34366
rect 19282 34302 19294 34354
rect 19346 34302 19358 34354
rect 20290 34302 20302 34354
rect 20354 34302 20366 34354
rect 15150 34290 15202 34302
rect 29150 34290 29202 34302
rect 29822 34354 29874 34366
rect 29822 34290 29874 34302
rect 34078 34354 34130 34366
rect 34078 34290 34130 34302
rect 41246 34354 41298 34366
rect 41246 34290 41298 34302
rect 41470 34354 41522 34366
rect 44270 34354 44322 34366
rect 42354 34302 42366 34354
rect 42418 34302 42430 34354
rect 41470 34290 41522 34302
rect 44270 34290 44322 34302
rect 44494 34354 44546 34366
rect 44494 34290 44546 34302
rect 54686 34354 54738 34366
rect 54686 34290 54738 34302
rect 8430 34242 8482 34254
rect 17950 34242 18002 34254
rect 10434 34190 10446 34242
rect 10498 34190 10510 34242
rect 10770 34190 10782 34242
rect 10834 34190 10846 34242
rect 8430 34178 8482 34190
rect 17950 34178 18002 34190
rect 30270 34242 30322 34254
rect 34638 34242 34690 34254
rect 30930 34190 30942 34242
rect 30994 34190 31006 34242
rect 31378 34190 31390 34242
rect 31442 34190 31454 34242
rect 30270 34178 30322 34190
rect 34638 34178 34690 34190
rect 47182 34242 47234 34254
rect 47182 34178 47234 34190
rect 54910 34242 54962 34254
rect 54910 34178 54962 34190
rect 56702 34242 56754 34254
rect 56702 34178 56754 34190
rect 7758 34130 7810 34142
rect 7758 34066 7810 34078
rect 8990 34130 9042 34142
rect 28702 34130 28754 34142
rect 10210 34078 10222 34130
rect 10274 34078 10286 34130
rect 16146 34078 16158 34130
rect 16210 34078 16222 34130
rect 17378 34078 17390 34130
rect 17442 34078 17454 34130
rect 20738 34078 20750 34130
rect 20802 34078 20814 34130
rect 23874 34078 23886 34130
rect 23938 34078 23950 34130
rect 28354 34078 28366 34130
rect 28418 34078 28430 34130
rect 8990 34066 9042 34078
rect 28702 34066 28754 34078
rect 28926 34130 28978 34142
rect 28926 34066 28978 34078
rect 30046 34130 30098 34142
rect 30046 34066 30098 34078
rect 30382 34130 30434 34142
rect 36318 34130 36370 34142
rect 39230 34130 39282 34142
rect 40126 34130 40178 34142
rect 30706 34078 30718 34130
rect 30770 34078 30782 34130
rect 31826 34078 31838 34130
rect 31890 34078 31902 34130
rect 34066 34078 34078 34130
rect 34130 34078 34142 34130
rect 36082 34078 36094 34130
rect 36146 34078 36158 34130
rect 37090 34078 37102 34130
rect 37154 34078 37166 34130
rect 39666 34078 39678 34130
rect 39730 34078 39742 34130
rect 30382 34066 30434 34078
rect 36318 34066 36370 34078
rect 39230 34066 39282 34078
rect 40126 34066 40178 34078
rect 41694 34130 41746 34142
rect 41694 34066 41746 34078
rect 42030 34130 42082 34142
rect 42030 34066 42082 34078
rect 43934 34130 43986 34142
rect 43934 34066 43986 34078
rect 44606 34130 44658 34142
rect 44606 34066 44658 34078
rect 45726 34130 45778 34142
rect 55022 34130 55074 34142
rect 45938 34078 45950 34130
rect 46002 34078 46014 34130
rect 45726 34066 45778 34078
rect 55022 34066 55074 34078
rect 57038 34130 57090 34142
rect 57038 34066 57090 34078
rect 57150 34130 57202 34142
rect 57150 34066 57202 34078
rect 11454 34018 11506 34030
rect 9538 33966 9550 34018
rect 9602 33966 9614 34018
rect 11454 33954 11506 33966
rect 16718 34018 16770 34030
rect 16718 33954 16770 33966
rect 19182 34018 19234 34030
rect 19182 33954 19234 33966
rect 21310 34018 21362 34030
rect 28814 34018 28866 34030
rect 33854 34018 33906 34030
rect 23538 33966 23550 34018
rect 23602 33966 23614 34018
rect 25442 33966 25454 34018
rect 25506 33966 25518 34018
rect 27570 33966 27582 34018
rect 27634 33966 27646 34018
rect 31602 33966 31614 34018
rect 31666 33966 31678 34018
rect 21310 33954 21362 33966
rect 28814 33954 28866 33966
rect 33854 33954 33906 33966
rect 37662 34018 37714 34030
rect 41582 34018 41634 34030
rect 38770 33966 38782 34018
rect 38834 33966 38846 34018
rect 37662 33954 37714 33966
rect 41582 33954 41634 33966
rect 46622 34018 46674 34030
rect 46622 33954 46674 33966
rect 46958 34018 47010 34030
rect 47742 34018 47794 34030
rect 47282 33966 47294 34018
rect 47346 33966 47358 34018
rect 46958 33954 47010 33966
rect 47742 33954 47794 33966
rect 56814 34018 56866 34030
rect 56814 33954 56866 33966
rect 9886 33906 9938 33918
rect 36082 33854 36094 33906
rect 36146 33854 36158 33906
rect 9886 33842 9938 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 57038 33570 57090 33582
rect 37538 33518 37550 33570
rect 37602 33518 37614 33570
rect 57038 33506 57090 33518
rect 57598 33570 57650 33582
rect 57598 33506 57650 33518
rect 14590 33458 14642 33470
rect 27918 33458 27970 33470
rect 10882 33406 10894 33458
rect 10946 33406 10958 33458
rect 12674 33406 12686 33458
rect 12738 33406 12750 33458
rect 14130 33406 14142 33458
rect 14194 33406 14206 33458
rect 19394 33406 19406 33458
rect 19458 33406 19470 33458
rect 24210 33406 24222 33458
rect 24274 33406 24286 33458
rect 14590 33394 14642 33406
rect 27918 33394 27970 33406
rect 38110 33458 38162 33470
rect 51202 33406 51214 33458
rect 51266 33406 51278 33458
rect 55570 33406 55582 33458
rect 55634 33406 55646 33458
rect 38110 33394 38162 33406
rect 20190 33346 20242 33358
rect 11218 33294 11230 33346
rect 11282 33294 11294 33346
rect 11666 33294 11678 33346
rect 11730 33294 11742 33346
rect 12226 33294 12238 33346
rect 12290 33294 12302 33346
rect 13010 33294 13022 33346
rect 13074 33294 13086 33346
rect 13794 33294 13806 33346
rect 13858 33294 13870 33346
rect 14802 33294 14814 33346
rect 14866 33294 14878 33346
rect 15810 33294 15822 33346
rect 15874 33294 15886 33346
rect 20190 33282 20242 33294
rect 20638 33346 20690 33358
rect 28142 33346 28194 33358
rect 21410 33294 21422 33346
rect 21474 33294 21486 33346
rect 20638 33282 20690 33294
rect 28142 33282 28194 33294
rect 28366 33346 28418 33358
rect 34302 33346 34354 33358
rect 39790 33346 39842 33358
rect 41694 33346 41746 33358
rect 31826 33294 31838 33346
rect 31890 33294 31902 33346
rect 33618 33294 33630 33346
rect 33682 33294 33694 33346
rect 35074 33294 35086 33346
rect 35138 33294 35150 33346
rect 36978 33294 36990 33346
rect 37042 33294 37054 33346
rect 38434 33294 38446 33346
rect 38498 33294 38510 33346
rect 38882 33294 38894 33346
rect 38946 33294 38958 33346
rect 40226 33294 40238 33346
rect 40290 33294 40302 33346
rect 41234 33294 41246 33346
rect 41298 33294 41310 33346
rect 28366 33282 28418 33294
rect 34302 33282 34354 33294
rect 39790 33282 39842 33294
rect 41694 33282 41746 33294
rect 42030 33346 42082 33358
rect 42030 33282 42082 33294
rect 42366 33346 42418 33358
rect 51886 33346 51938 33358
rect 57150 33346 57202 33358
rect 43922 33294 43934 33346
rect 43986 33294 43998 33346
rect 48290 33294 48302 33346
rect 48354 33294 48366 33346
rect 52770 33294 52782 33346
rect 52834 33294 52846 33346
rect 42366 33282 42418 33294
rect 51886 33282 51938 33294
rect 57150 33282 57202 33294
rect 57486 33346 57538 33358
rect 57486 33282 57538 33294
rect 27806 33234 27858 33246
rect 51550 33234 51602 33246
rect 14242 33182 14254 33234
rect 14306 33182 14318 33234
rect 16706 33182 16718 33234
rect 16770 33182 16782 33234
rect 22082 33182 22094 33234
rect 22146 33182 22158 33234
rect 25778 33182 25790 33234
rect 25842 33182 25854 33234
rect 32386 33182 32398 33234
rect 32450 33182 32462 33234
rect 39106 33182 39118 33234
rect 39170 33182 39182 33234
rect 43698 33182 43710 33234
rect 43762 33182 43774 33234
rect 49074 33182 49086 33234
rect 49138 33182 49150 33234
rect 27806 33170 27858 33182
rect 51550 33170 51602 33182
rect 51998 33234 52050 33246
rect 51998 33170 52050 33182
rect 52110 33234 52162 33246
rect 53442 33182 53454 33234
rect 53506 33182 53518 33234
rect 52110 33170 52162 33182
rect 19966 33122 20018 33134
rect 19966 33058 20018 33070
rect 20078 33122 20130 33134
rect 20078 33058 20130 33070
rect 24670 33122 24722 33134
rect 24670 33058 24722 33070
rect 25118 33122 25170 33134
rect 25118 33058 25170 33070
rect 25454 33122 25506 33134
rect 25454 33058 25506 33070
rect 27582 33122 27634 33134
rect 27582 33058 27634 33070
rect 29486 33122 29538 33134
rect 31278 33122 31330 33134
rect 30930 33070 30942 33122
rect 30994 33070 31006 33122
rect 29486 33058 29538 33070
rect 31278 33058 31330 33070
rect 31502 33122 31554 33134
rect 31502 33058 31554 33070
rect 36206 33122 36258 33134
rect 36206 33058 36258 33070
rect 42030 33122 42082 33134
rect 42030 33058 42082 33070
rect 56030 33122 56082 33134
rect 56030 33058 56082 33070
rect 57038 33122 57090 33134
rect 57038 33058 57090 33070
rect 57598 33122 57650 33134
rect 57598 33058 57650 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 10670 32786 10722 32798
rect 8978 32734 8990 32786
rect 9042 32734 9054 32786
rect 10670 32722 10722 32734
rect 11902 32786 11954 32798
rect 11902 32722 11954 32734
rect 15150 32786 15202 32798
rect 18622 32786 18674 32798
rect 17602 32734 17614 32786
rect 17666 32734 17678 32786
rect 15150 32722 15202 32734
rect 18622 32722 18674 32734
rect 19406 32786 19458 32798
rect 19406 32722 19458 32734
rect 20414 32786 20466 32798
rect 20414 32722 20466 32734
rect 24110 32786 24162 32798
rect 33182 32786 33234 32798
rect 24434 32734 24446 32786
rect 24498 32734 24510 32786
rect 32050 32734 32062 32786
rect 32114 32734 32126 32786
rect 24110 32722 24162 32734
rect 33182 32722 33234 32734
rect 39006 32786 39058 32798
rect 39006 32722 39058 32734
rect 43374 32786 43426 32798
rect 43374 32722 43426 32734
rect 49086 32786 49138 32798
rect 49086 32722 49138 32734
rect 51774 32786 51826 32798
rect 51774 32722 51826 32734
rect 53902 32786 53954 32798
rect 55122 32734 55134 32786
rect 55186 32734 55198 32786
rect 53902 32722 53954 32734
rect 14926 32674 14978 32686
rect 14578 32622 14590 32674
rect 14642 32622 14654 32674
rect 14926 32610 14978 32622
rect 16046 32674 16098 32686
rect 16046 32610 16098 32622
rect 18846 32674 18898 32686
rect 18846 32610 18898 32622
rect 19070 32674 19122 32686
rect 19070 32610 19122 32622
rect 40462 32674 40514 32686
rect 40462 32610 40514 32622
rect 41806 32674 41858 32686
rect 41806 32610 41858 32622
rect 50654 32674 50706 32686
rect 50654 32610 50706 32622
rect 51998 32674 52050 32686
rect 51998 32610 52050 32622
rect 52110 32674 52162 32686
rect 52110 32610 52162 32622
rect 52894 32674 52946 32686
rect 52894 32610 52946 32622
rect 53230 32674 53282 32686
rect 53230 32610 53282 32622
rect 54014 32674 54066 32686
rect 54014 32610 54066 32622
rect 54798 32674 54850 32686
rect 54798 32610 54850 32622
rect 10334 32562 10386 32574
rect 8754 32510 8766 32562
rect 8818 32510 8830 32562
rect 10334 32498 10386 32510
rect 11566 32562 11618 32574
rect 16382 32562 16434 32574
rect 12786 32510 12798 32562
rect 12850 32510 12862 32562
rect 13570 32510 13582 32562
rect 13634 32510 13646 32562
rect 15362 32510 15374 32562
rect 15426 32510 15438 32562
rect 11566 32498 11618 32510
rect 16382 32498 16434 32510
rect 16830 32562 16882 32574
rect 18510 32562 18562 32574
rect 18162 32510 18174 32562
rect 18226 32510 18238 32562
rect 16830 32498 16882 32510
rect 18510 32498 18562 32510
rect 19966 32562 20018 32574
rect 34526 32562 34578 32574
rect 40910 32562 40962 32574
rect 31602 32510 31614 32562
rect 31666 32510 31678 32562
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 34850 32510 34862 32562
rect 34914 32510 34926 32562
rect 37202 32510 37214 32562
rect 37266 32510 37278 32562
rect 37986 32510 37998 32562
rect 38050 32510 38062 32562
rect 38434 32510 38446 32562
rect 38498 32510 38510 32562
rect 19966 32498 20018 32510
rect 34526 32498 34578 32510
rect 40910 32498 40962 32510
rect 41470 32562 41522 32574
rect 41470 32498 41522 32510
rect 43934 32562 43986 32574
rect 43934 32498 43986 32510
rect 44158 32562 44210 32574
rect 44942 32562 44994 32574
rect 47406 32562 47458 32574
rect 44482 32510 44494 32562
rect 44546 32510 44558 32562
rect 46722 32510 46734 32562
rect 46786 32510 46798 32562
rect 44158 32498 44210 32510
rect 44942 32498 44994 32510
rect 47406 32498 47458 32510
rect 48974 32562 49026 32574
rect 48974 32498 49026 32510
rect 49198 32562 49250 32574
rect 49198 32498 49250 32510
rect 49646 32562 49698 32574
rect 49646 32498 49698 32510
rect 50318 32562 50370 32574
rect 50318 32498 50370 32510
rect 50430 32562 50482 32574
rect 50430 32498 50482 32510
rect 50878 32562 50930 32574
rect 50878 32498 50930 32510
rect 20302 32450 20354 32462
rect 10546 32398 10558 32450
rect 10610 32398 10622 32450
rect 13122 32398 13134 32450
rect 13186 32398 13198 32450
rect 20302 32386 20354 32398
rect 21086 32450 21138 32462
rect 21086 32386 21138 32398
rect 28590 32450 28642 32462
rect 43598 32450 43650 32462
rect 32162 32398 32174 32450
rect 32226 32398 32238 32450
rect 36306 32398 36318 32450
rect 36370 32398 36382 32450
rect 37650 32398 37662 32450
rect 37714 32398 37726 32450
rect 42242 32398 42254 32450
rect 42306 32398 42318 32450
rect 28590 32386 28642 32398
rect 43598 32386 43650 32398
rect 44046 32450 44098 32462
rect 51438 32450 51490 32462
rect 46498 32398 46510 32450
rect 46562 32398 46574 32450
rect 44046 32386 44098 32398
rect 51438 32386 51490 32398
rect 58158 32450 58210 32462
rect 58158 32386 58210 32398
rect 14814 32338 14866 32350
rect 14814 32274 14866 32286
rect 43262 32338 43314 32350
rect 43262 32274 43314 32286
rect 53902 32338 53954 32350
rect 53902 32274 53954 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 35758 32002 35810 32014
rect 44046 32002 44098 32014
rect 43698 31950 43710 32002
rect 43762 31950 43774 32002
rect 49858 31950 49870 32002
rect 49922 31950 49934 32002
rect 35758 31938 35810 31950
rect 44046 31938 44098 31950
rect 8654 31890 8706 31902
rect 7298 31838 7310 31890
rect 7362 31838 7374 31890
rect 8654 31826 8706 31838
rect 12462 31890 12514 31902
rect 19854 31890 19906 31902
rect 42142 31890 42194 31902
rect 14242 31838 14254 31890
rect 14306 31838 14318 31890
rect 18274 31838 18286 31890
rect 18338 31838 18350 31890
rect 18610 31838 18622 31890
rect 18674 31838 18686 31890
rect 26786 31838 26798 31890
rect 26850 31838 26862 31890
rect 30818 31838 30830 31890
rect 30882 31838 30894 31890
rect 32610 31838 32622 31890
rect 32674 31838 32686 31890
rect 34738 31838 34750 31890
rect 34802 31838 34814 31890
rect 37090 31838 37102 31890
rect 37154 31838 37166 31890
rect 39554 31838 39566 31890
rect 39618 31838 39630 31890
rect 41682 31838 41694 31890
rect 41746 31838 41758 31890
rect 45378 31838 45390 31890
rect 45442 31838 45454 31890
rect 56018 31838 56030 31890
rect 56082 31838 56094 31890
rect 58146 31838 58158 31890
rect 58210 31838 58222 31890
rect 12462 31826 12514 31838
rect 19854 31826 19906 31838
rect 42142 31826 42194 31838
rect 12126 31778 12178 31790
rect 13694 31778 13746 31790
rect 7186 31726 7198 31778
rect 7250 31726 7262 31778
rect 8082 31726 8094 31778
rect 8146 31726 8158 31778
rect 8866 31726 8878 31778
rect 8930 31726 8942 31778
rect 10658 31726 10670 31778
rect 10722 31726 10734 31778
rect 11330 31726 11342 31778
rect 11394 31726 11406 31778
rect 12338 31726 12350 31778
rect 12402 31726 12414 31778
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 12126 31714 12178 31726
rect 13694 31714 13746 31726
rect 13806 31778 13858 31790
rect 19406 31778 19458 31790
rect 33294 31778 33346 31790
rect 15474 31726 15486 31778
rect 15538 31726 15550 31778
rect 23874 31726 23886 31778
rect 23938 31726 23950 31778
rect 31154 31726 31166 31778
rect 31218 31726 31230 31778
rect 32946 31726 32958 31778
rect 33010 31726 33022 31778
rect 13806 31714 13858 31726
rect 19406 31714 19458 31726
rect 33294 31714 33346 31726
rect 34526 31778 34578 31790
rect 34526 31714 34578 31726
rect 35198 31778 35250 31790
rect 35198 31714 35250 31726
rect 35422 31778 35474 31790
rect 37886 31778 37938 31790
rect 44270 31778 44322 31790
rect 49310 31778 49362 31790
rect 37426 31726 37438 31778
rect 37490 31726 37502 31778
rect 38210 31726 38222 31778
rect 38274 31726 38286 31778
rect 38770 31726 38782 31778
rect 38834 31726 38846 31778
rect 48290 31726 48302 31778
rect 48354 31726 48366 31778
rect 50082 31726 50094 31778
rect 50146 31726 50158 31778
rect 55234 31726 55246 31778
rect 55298 31726 55310 31778
rect 35422 31714 35474 31726
rect 37886 31714 37938 31726
rect 44270 31714 44322 31726
rect 49310 31714 49362 31726
rect 49422 31666 49474 31678
rect 16146 31614 16158 31666
rect 16210 31614 16222 31666
rect 24658 31614 24670 31666
rect 24722 31614 24734 31666
rect 47506 31614 47518 31666
rect 47570 31614 47582 31666
rect 49522 31614 49534 31666
rect 49586 31614 49598 31666
rect 49422 31602 49474 31614
rect 15038 31554 15090 31566
rect 15038 31490 15090 31502
rect 27246 31554 27298 31566
rect 27246 31490 27298 31502
rect 48750 31554 48802 31566
rect 50766 31554 50818 31566
rect 50418 31502 50430 31554
rect 50482 31502 50494 31554
rect 48750 31490 48802 31502
rect 50766 31490 50818 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 14030 31218 14082 31230
rect 14030 31154 14082 31166
rect 22542 31218 22594 31230
rect 22542 31154 22594 31166
rect 22766 31218 22818 31230
rect 22766 31154 22818 31166
rect 23326 31218 23378 31230
rect 23326 31154 23378 31166
rect 24110 31218 24162 31230
rect 34526 31218 34578 31230
rect 31042 31166 31054 31218
rect 31106 31166 31118 31218
rect 24110 31154 24162 31166
rect 34526 31154 34578 31166
rect 48974 31218 49026 31230
rect 48974 31154 49026 31166
rect 56926 31218 56978 31230
rect 56926 31154 56978 31166
rect 14478 31106 14530 31118
rect 14478 31042 14530 31054
rect 21982 31106 22034 31118
rect 21982 31042 22034 31054
rect 22094 31106 22146 31118
rect 49982 31106 50034 31118
rect 57822 31106 57874 31118
rect 43026 31054 43038 31106
rect 43090 31054 43102 31106
rect 55346 31054 55358 31106
rect 55410 31054 55422 31106
rect 22094 31042 22146 31054
rect 49982 31042 50034 31054
rect 57822 31042 57874 31054
rect 58158 31106 58210 31118
rect 58158 31042 58210 31054
rect 22318 30994 22370 31006
rect 7186 30942 7198 30994
rect 7250 30942 7262 30994
rect 9986 30942 9998 30994
rect 10050 30942 10062 30994
rect 11778 30942 11790 30994
rect 11842 30942 11854 30994
rect 13906 30942 13918 30994
rect 13970 30942 13982 30994
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 22318 30930 22370 30942
rect 22878 30994 22930 31006
rect 22878 30930 22930 30942
rect 23102 30994 23154 31006
rect 23102 30930 23154 30942
rect 23438 30994 23490 31006
rect 23438 30930 23490 30942
rect 23998 30994 24050 31006
rect 23998 30930 24050 30942
rect 24334 30994 24386 31006
rect 56590 30994 56642 31006
rect 28130 30942 28142 30994
rect 28194 30942 28206 30994
rect 42354 30942 42366 30994
rect 42418 30942 42430 30994
rect 55122 30942 55134 30994
rect 55186 30942 55198 30994
rect 24334 30930 24386 30942
rect 56590 30930 56642 30942
rect 56814 30994 56866 31006
rect 56814 30930 56866 30942
rect 57262 30994 57314 31006
rect 57262 30930 57314 30942
rect 15710 30882 15762 30894
rect 12226 30830 12238 30882
rect 12290 30830 12302 30882
rect 15710 30818 15762 30830
rect 21198 30882 21250 30894
rect 25454 30882 25506 30894
rect 22082 30830 22094 30882
rect 22146 30830 22158 30882
rect 21198 30818 21250 30830
rect 25454 30818 25506 30830
rect 27694 30882 27746 30894
rect 45614 30882 45666 30894
rect 28802 30830 28814 30882
rect 28866 30830 28878 30882
rect 45154 30830 45166 30882
rect 45218 30830 45230 30882
rect 49858 30830 49870 30882
rect 49922 30830 49934 30882
rect 27694 30818 27746 30830
rect 45614 30818 45666 30830
rect 7758 30770 7810 30782
rect 50206 30770 50258 30782
rect 11554 30718 11566 30770
rect 11618 30718 11630 30770
rect 7758 30706 7810 30718
rect 50206 30706 50258 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 46510 30434 46562 30446
rect 46510 30370 46562 30382
rect 11342 30322 11394 30334
rect 31950 30322 32002 30334
rect 16034 30270 16046 30322
rect 16098 30270 16110 30322
rect 21522 30270 21534 30322
rect 21586 30270 21598 30322
rect 24994 30270 25006 30322
rect 25058 30270 25070 30322
rect 28578 30270 28590 30322
rect 28642 30270 28654 30322
rect 29138 30270 29150 30322
rect 29202 30270 29214 30322
rect 11342 30258 11394 30270
rect 31950 30258 32002 30270
rect 32510 30322 32562 30334
rect 35074 30270 35086 30322
rect 35138 30270 35150 30322
rect 39890 30270 39902 30322
rect 39954 30270 39966 30322
rect 46946 30270 46958 30322
rect 47010 30270 47022 30322
rect 56018 30270 56030 30322
rect 56082 30270 56094 30322
rect 58146 30270 58158 30322
rect 58210 30270 58222 30322
rect 32510 30258 32562 30270
rect 9662 30210 9714 30222
rect 19070 30210 19122 30222
rect 8194 30158 8206 30210
rect 8258 30158 8270 30210
rect 13570 30158 13582 30210
rect 13634 30158 13646 30210
rect 13794 30158 13806 30210
rect 13858 30158 13870 30210
rect 14130 30158 14142 30210
rect 14194 30158 14206 30210
rect 9662 30146 9714 30158
rect 19070 30146 19122 30158
rect 19630 30210 19682 30222
rect 19630 30146 19682 30158
rect 22318 30210 22370 30222
rect 30158 30210 30210 30222
rect 34638 30210 34690 30222
rect 46622 30210 46674 30222
rect 50206 30210 50258 30222
rect 25778 30158 25790 30210
rect 25842 30158 25854 30210
rect 34290 30158 34302 30210
rect 34354 30158 34366 30210
rect 35746 30158 35758 30210
rect 35810 30158 35822 30210
rect 37090 30158 37102 30210
rect 37154 30158 37166 30210
rect 49858 30158 49870 30210
rect 49922 30158 49934 30210
rect 22318 30146 22370 30158
rect 30158 30146 30210 30158
rect 34638 30146 34690 30158
rect 46622 30146 46674 30158
rect 50206 30146 50258 30158
rect 50878 30210 50930 30222
rect 52670 30210 52722 30222
rect 51538 30158 51550 30210
rect 51602 30158 51614 30210
rect 55346 30158 55358 30210
rect 55410 30158 55422 30210
rect 50878 30146 50930 30158
rect 52670 30146 52722 30158
rect 10110 30098 10162 30110
rect 16494 30098 16546 30110
rect 16370 30046 16382 30098
rect 16434 30046 16446 30098
rect 10110 30034 10162 30046
rect 16494 30034 16546 30046
rect 17054 30098 17106 30110
rect 17054 30034 17106 30046
rect 17278 30098 17330 30110
rect 17278 30034 17330 30046
rect 17390 30098 17442 30110
rect 21982 30098 22034 30110
rect 21746 30046 21758 30098
rect 21810 30046 21822 30098
rect 17390 30034 17442 30046
rect 21982 30034 22034 30046
rect 22094 30098 22146 30110
rect 22094 30034 22146 30046
rect 24222 30098 24274 30110
rect 24222 30034 24274 30046
rect 24558 30098 24610 30110
rect 29598 30098 29650 30110
rect 24770 30046 24782 30098
rect 24834 30046 24846 30098
rect 26450 30046 26462 30098
rect 26514 30046 26526 30098
rect 29474 30046 29486 30098
rect 29538 30046 29550 30098
rect 24558 30034 24610 30046
rect 29598 30034 29650 30046
rect 30382 30098 30434 30110
rect 30382 30034 30434 30046
rect 30494 30098 30546 30110
rect 30494 30034 30546 30046
rect 31166 30098 31218 30110
rect 31166 30034 31218 30046
rect 31278 30098 31330 30110
rect 31278 30034 31330 30046
rect 33294 30098 33346 30110
rect 51774 30098 51826 30110
rect 37762 30046 37774 30098
rect 37826 30046 37838 30098
rect 49074 30046 49086 30098
rect 49138 30046 49150 30098
rect 33294 30034 33346 30046
rect 51774 30034 51826 30046
rect 7758 29986 7810 29998
rect 7758 29922 7810 29934
rect 9662 29986 9714 29998
rect 9662 29922 9714 29934
rect 14814 29986 14866 29998
rect 14814 29922 14866 29934
rect 16606 29986 16658 29998
rect 16606 29922 16658 29934
rect 16830 29986 16882 29998
rect 16830 29922 16882 29934
rect 17838 29986 17890 29998
rect 17838 29922 17890 29934
rect 22878 29986 22930 29998
rect 22878 29922 22930 29934
rect 24446 29986 24498 29998
rect 24446 29922 24498 29934
rect 29710 29986 29762 29998
rect 29710 29922 29762 29934
rect 29934 29986 29986 29998
rect 29934 29922 29986 29934
rect 31502 29986 31554 29998
rect 31502 29922 31554 29934
rect 35534 29986 35586 29998
rect 35534 29922 35586 29934
rect 36542 29986 36594 29998
rect 36542 29922 36594 29934
rect 40350 29986 40402 29998
rect 40350 29922 40402 29934
rect 46510 29986 46562 29998
rect 46510 29922 46562 29934
rect 50318 29986 50370 29998
rect 50318 29922 50370 29934
rect 50542 29986 50594 29998
rect 50542 29922 50594 29934
rect 53006 29986 53058 29998
rect 53006 29922 53058 29934
rect 54574 29986 54626 29998
rect 54898 29934 54910 29986
rect 54962 29934 54974 29986
rect 54574 29922 54626 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 21870 29650 21922 29662
rect 10434 29598 10446 29650
rect 10498 29598 10510 29650
rect 20402 29598 20414 29650
rect 20466 29598 20478 29650
rect 21870 29586 21922 29598
rect 22318 29650 22370 29662
rect 22318 29586 22370 29598
rect 23214 29650 23266 29662
rect 25566 29650 25618 29662
rect 24322 29598 24334 29650
rect 24386 29598 24398 29650
rect 23214 29586 23266 29598
rect 25566 29586 25618 29598
rect 26910 29650 26962 29662
rect 26910 29586 26962 29598
rect 27806 29650 27858 29662
rect 27806 29586 27858 29598
rect 28030 29650 28082 29662
rect 28030 29586 28082 29598
rect 28702 29650 28754 29662
rect 28702 29586 28754 29598
rect 34414 29650 34466 29662
rect 35310 29650 35362 29662
rect 34738 29598 34750 29650
rect 34802 29598 34814 29650
rect 34414 29586 34466 29598
rect 35310 29586 35362 29598
rect 37214 29650 37266 29662
rect 37214 29586 37266 29598
rect 42926 29650 42978 29662
rect 51102 29650 51154 29662
rect 43474 29598 43486 29650
rect 43538 29598 43550 29650
rect 42926 29586 42978 29598
rect 51102 29586 51154 29598
rect 53118 29650 53170 29662
rect 53118 29586 53170 29598
rect 56702 29650 56754 29662
rect 56702 29586 56754 29598
rect 56926 29650 56978 29662
rect 56926 29586 56978 29598
rect 57822 29650 57874 29662
rect 57822 29586 57874 29598
rect 12350 29538 12402 29550
rect 9762 29486 9774 29538
rect 9826 29486 9838 29538
rect 11330 29486 11342 29538
rect 11394 29486 11406 29538
rect 12350 29474 12402 29486
rect 21534 29538 21586 29550
rect 21534 29474 21586 29486
rect 21646 29538 21698 29550
rect 21646 29474 21698 29486
rect 22094 29538 22146 29550
rect 22094 29474 22146 29486
rect 22430 29538 22482 29550
rect 23662 29538 23714 29550
rect 27694 29538 27746 29550
rect 22866 29486 22878 29538
rect 22930 29486 22942 29538
rect 25218 29486 25230 29538
rect 25282 29486 25294 29538
rect 27570 29486 27582 29538
rect 27634 29486 27646 29538
rect 22430 29474 22482 29486
rect 23662 29474 23714 29486
rect 27694 29474 27746 29486
rect 28478 29538 28530 29550
rect 28478 29474 28530 29486
rect 30718 29538 30770 29550
rect 30718 29474 30770 29486
rect 30942 29538 30994 29550
rect 51550 29538 51602 29550
rect 57038 29538 57090 29550
rect 31266 29486 31278 29538
rect 31330 29486 31342 29538
rect 53442 29486 53454 29538
rect 53506 29486 53518 29538
rect 30942 29474 30994 29486
rect 51550 29474 51602 29486
rect 57038 29474 57090 29486
rect 23998 29426 24050 29438
rect 28814 29426 28866 29438
rect 36878 29426 36930 29438
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 7746 29374 7758 29426
rect 7810 29374 7822 29426
rect 9538 29374 9550 29426
rect 9602 29374 9614 29426
rect 10546 29374 10558 29426
rect 10610 29374 10622 29426
rect 13458 29374 13470 29426
rect 13522 29374 13534 29426
rect 14242 29374 14254 29426
rect 14306 29374 14318 29426
rect 15138 29374 15150 29426
rect 15202 29374 15214 29426
rect 15586 29374 15598 29426
rect 15650 29374 15662 29426
rect 17378 29374 17390 29426
rect 17442 29374 17454 29426
rect 21074 29374 21086 29426
rect 21138 29374 21150 29426
rect 24546 29374 24558 29426
rect 24610 29374 24622 29426
rect 31154 29374 31166 29426
rect 31218 29374 31230 29426
rect 35634 29374 35646 29426
rect 35698 29374 35710 29426
rect 23998 29362 24050 29374
rect 28814 29362 28866 29374
rect 36878 29362 36930 29374
rect 36990 29426 37042 29438
rect 36990 29362 37042 29374
rect 37438 29426 37490 29438
rect 37438 29362 37490 29374
rect 50990 29426 51042 29438
rect 50990 29362 51042 29374
rect 51214 29426 51266 29438
rect 51214 29362 51266 29374
rect 11006 29314 11058 29326
rect 29262 29314 29314 29326
rect 5058 29262 5070 29314
rect 5122 29262 5134 29314
rect 7186 29262 7198 29314
rect 7250 29262 7262 29314
rect 8530 29262 8542 29314
rect 8594 29262 8606 29314
rect 18162 29262 18174 29314
rect 18226 29262 18238 29314
rect 21522 29262 21534 29314
rect 21586 29262 21598 29314
rect 27682 29262 27694 29314
rect 27746 29262 27758 29314
rect 11006 29250 11058 29262
rect 29262 29250 29314 29262
rect 29710 29314 29762 29326
rect 31950 29314 32002 29326
rect 40238 29314 40290 29326
rect 31490 29262 31502 29314
rect 31554 29262 31566 29314
rect 35970 29262 35982 29314
rect 36034 29262 36046 29314
rect 29710 29250 29762 29262
rect 31950 29250 32002 29262
rect 40238 29250 40290 29262
rect 44046 29314 44098 29326
rect 44046 29250 44098 29262
rect 53902 29314 53954 29326
rect 53902 29250 53954 29262
rect 58158 29314 58210 29326
rect 58158 29250 58210 29262
rect 40126 29202 40178 29214
rect 13458 29150 13470 29202
rect 13522 29150 13534 29202
rect 40126 29138 40178 29150
rect 42814 29202 42866 29214
rect 42814 29138 42866 29150
rect 43150 29202 43202 29214
rect 43150 29138 43202 29150
rect 43822 29202 43874 29214
rect 43822 29138 43874 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 18174 28866 18226 28878
rect 18174 28802 18226 28814
rect 9102 28754 9154 28766
rect 9102 28690 9154 28702
rect 11118 28754 11170 28766
rect 15822 28754 15874 28766
rect 13458 28702 13470 28754
rect 13522 28702 13534 28754
rect 14914 28702 14926 28754
rect 14978 28702 14990 28754
rect 11118 28690 11170 28702
rect 15822 28690 15874 28702
rect 19630 28754 19682 28766
rect 37886 28754 37938 28766
rect 41918 28754 41970 28766
rect 31938 28702 31950 28754
rect 32002 28702 32014 28754
rect 34066 28702 34078 28754
rect 34130 28702 34142 28754
rect 41458 28702 41470 28754
rect 41522 28702 41534 28754
rect 19630 28690 19682 28702
rect 37886 28690 37938 28702
rect 41918 28690 41970 28702
rect 43486 28754 43538 28766
rect 43486 28690 43538 28702
rect 45278 28754 45330 28766
rect 49534 28754 49586 28766
rect 48514 28702 48526 28754
rect 48578 28702 48590 28754
rect 45278 28690 45330 28702
rect 49534 28690 49586 28702
rect 49758 28754 49810 28766
rect 49758 28690 49810 28702
rect 50654 28754 50706 28766
rect 56578 28702 56590 28754
rect 56642 28702 56654 28754
rect 50654 28690 50706 28702
rect 6974 28642 7026 28654
rect 16606 28642 16658 28654
rect 18062 28642 18114 28654
rect 7298 28590 7310 28642
rect 7362 28590 7374 28642
rect 12898 28590 12910 28642
rect 12962 28590 12974 28642
rect 15362 28590 15374 28642
rect 15426 28590 15438 28642
rect 17378 28590 17390 28642
rect 17442 28590 17454 28642
rect 6974 28578 7026 28590
rect 16606 28578 16658 28590
rect 18062 28578 18114 28590
rect 19182 28642 19234 28654
rect 19182 28578 19234 28590
rect 30270 28642 30322 28654
rect 30270 28578 30322 28590
rect 30606 28642 30658 28654
rect 30606 28578 30658 28590
rect 30942 28642 30994 28654
rect 34862 28642 34914 28654
rect 37326 28642 37378 28654
rect 42702 28642 42754 28654
rect 53230 28642 53282 28654
rect 31154 28590 31166 28642
rect 31218 28590 31230 28642
rect 35298 28590 35310 28642
rect 35362 28590 35374 28642
rect 35858 28590 35870 28642
rect 35922 28590 35934 28642
rect 38658 28590 38670 28642
rect 38722 28590 38734 28642
rect 43026 28590 43038 28642
rect 43090 28590 43102 28642
rect 45602 28590 45614 28642
rect 45666 28590 45678 28642
rect 52770 28590 52782 28642
rect 52834 28590 52846 28642
rect 54226 28590 54238 28642
rect 54290 28590 54302 28642
rect 30942 28578 30994 28590
rect 34862 28578 34914 28590
rect 37326 28578 37378 28590
rect 42702 28578 42754 28590
rect 53230 28578 53282 28590
rect 7870 28530 7922 28542
rect 7870 28466 7922 28478
rect 12350 28530 12402 28542
rect 13918 28530 13970 28542
rect 13682 28478 13694 28530
rect 13746 28478 13758 28530
rect 12350 28466 12402 28478
rect 13918 28466 13970 28478
rect 14814 28530 14866 28542
rect 14814 28466 14866 28478
rect 14926 28530 14978 28542
rect 18174 28530 18226 28542
rect 30718 28530 30770 28542
rect 37774 28530 37826 28542
rect 17490 28478 17502 28530
rect 17554 28478 17566 28530
rect 18834 28478 18846 28530
rect 18898 28478 18910 28530
rect 36082 28478 36094 28530
rect 36146 28478 36158 28530
rect 14926 28466 14978 28478
rect 18174 28466 18226 28478
rect 30718 28466 30770 28478
rect 37774 28466 37826 28478
rect 37998 28530 38050 28542
rect 53566 28530 53618 28542
rect 39330 28478 39342 28530
rect 39394 28478 39406 28530
rect 46386 28478 46398 28530
rect 46450 28478 46462 28530
rect 37998 28466 38050 28478
rect 53566 28466 53618 28478
rect 7422 28418 7474 28430
rect 7422 28354 7474 28366
rect 12798 28418 12850 28430
rect 12798 28354 12850 28366
rect 14030 28418 14082 28430
rect 14030 28354 14082 28366
rect 14254 28418 14306 28430
rect 14254 28354 14306 28366
rect 14590 28418 14642 28430
rect 14590 28354 14642 28366
rect 16942 28418 16994 28430
rect 16942 28354 16994 28366
rect 17054 28418 17106 28430
rect 17054 28354 17106 28366
rect 17166 28418 17218 28430
rect 17166 28354 17218 28366
rect 20750 28418 20802 28430
rect 20750 28354 20802 28366
rect 43374 28418 43426 28430
rect 43374 28354 43426 28366
rect 43598 28418 43650 28430
rect 53454 28418 53506 28430
rect 50082 28366 50094 28418
rect 50146 28366 50158 28418
rect 52994 28366 53006 28418
rect 53058 28366 53070 28418
rect 43598 28354 43650 28366
rect 53454 28354 53506 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 8654 28082 8706 28094
rect 8654 28018 8706 28030
rect 13246 28082 13298 28094
rect 13246 28018 13298 28030
rect 14478 28082 14530 28094
rect 14478 28018 14530 28030
rect 15038 28082 15090 28094
rect 15038 28018 15090 28030
rect 15822 28082 15874 28094
rect 15822 28018 15874 28030
rect 18174 28082 18226 28094
rect 18174 28018 18226 28030
rect 28254 28082 28306 28094
rect 30830 28082 30882 28094
rect 29026 28030 29038 28082
rect 29090 28030 29102 28082
rect 28254 28018 28306 28030
rect 30830 28018 30882 28030
rect 35086 28082 35138 28094
rect 35086 28018 35138 28030
rect 35758 28082 35810 28094
rect 35758 28018 35810 28030
rect 38894 28082 38946 28094
rect 38894 28018 38946 28030
rect 44382 28082 44434 28094
rect 44382 28018 44434 28030
rect 54686 28082 54738 28094
rect 54686 28018 54738 28030
rect 56590 28082 56642 28094
rect 56590 28018 56642 28030
rect 57374 28082 57426 28094
rect 57374 28018 57426 28030
rect 14702 27970 14754 27982
rect 11442 27918 11454 27970
rect 11506 27918 11518 27970
rect 14702 27906 14754 27918
rect 15262 27970 15314 27982
rect 31054 27970 31106 27982
rect 20290 27918 20302 27970
rect 20354 27918 20366 27970
rect 15262 27906 15314 27918
rect 31054 27906 31106 27918
rect 32062 27970 32114 27982
rect 32062 27906 32114 27918
rect 38110 27970 38162 27982
rect 38110 27906 38162 27918
rect 38222 27970 38274 27982
rect 38222 27906 38274 27918
rect 38446 27970 38498 27982
rect 38446 27906 38498 27918
rect 39006 27970 39058 27982
rect 57262 27970 57314 27982
rect 39106 27918 39118 27970
rect 39170 27918 39182 27970
rect 41794 27918 41806 27970
rect 41858 27918 41870 27970
rect 55458 27918 55470 27970
rect 55522 27918 55534 27970
rect 56914 27918 56926 27970
rect 56978 27918 56990 27970
rect 39006 27906 39058 27918
rect 57262 27906 57314 27918
rect 57934 27970 57986 27982
rect 57934 27906 57986 27918
rect 13134 27858 13186 27870
rect 14814 27858 14866 27870
rect 4722 27806 4734 27858
rect 4786 27806 4798 27858
rect 7970 27806 7982 27858
rect 8034 27806 8046 27858
rect 12114 27806 12126 27858
rect 12178 27806 12190 27858
rect 13458 27806 13470 27858
rect 13522 27806 13534 27858
rect 13134 27794 13186 27806
rect 14814 27794 14866 27806
rect 15374 27858 15426 27870
rect 22878 27858 22930 27870
rect 28702 27858 28754 27870
rect 32510 27858 32562 27870
rect 19618 27806 19630 27858
rect 19682 27806 19694 27858
rect 25778 27806 25790 27858
rect 25842 27806 25854 27858
rect 31266 27806 31278 27858
rect 31330 27806 31342 27858
rect 31490 27806 31502 27858
rect 31554 27806 31566 27858
rect 15374 27794 15426 27806
rect 22878 27794 22930 27806
rect 28702 27794 28754 27806
rect 32510 27794 32562 27806
rect 34526 27858 34578 27870
rect 34526 27794 34578 27806
rect 38670 27858 38722 27870
rect 55134 27858 55186 27870
rect 41122 27806 41134 27858
rect 41186 27806 41198 27858
rect 51426 27806 51438 27858
rect 51490 27806 51502 27858
rect 38670 27794 38722 27806
rect 55134 27794 55186 27806
rect 57822 27858 57874 27870
rect 57822 27794 57874 27806
rect 9662 27746 9714 27758
rect 18622 27746 18674 27758
rect 37774 27746 37826 27758
rect 5394 27694 5406 27746
rect 5458 27694 5470 27746
rect 7522 27694 7534 27746
rect 7586 27694 7598 27746
rect 12338 27694 12350 27746
rect 12402 27694 12414 27746
rect 22418 27694 22430 27746
rect 22482 27694 22494 27746
rect 26338 27694 26350 27746
rect 26402 27694 26414 27746
rect 31602 27694 31614 27746
rect 31666 27694 31678 27746
rect 39442 27694 39454 27746
rect 39506 27694 39518 27746
rect 43922 27694 43934 27746
rect 43986 27694 43998 27746
rect 52098 27694 52110 27746
rect 52162 27694 52174 27746
rect 54226 27694 54238 27746
rect 54290 27694 54302 27746
rect 9662 27682 9714 27694
rect 18622 27682 18674 27694
rect 37774 27682 37826 27694
rect 57374 27634 57426 27646
rect 57374 27570 57426 27582
rect 57934 27634 57986 27646
rect 57934 27570 57986 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 24558 27298 24610 27310
rect 7858 27246 7870 27298
rect 7922 27246 7934 27298
rect 8530 27246 8542 27298
rect 8594 27246 8606 27298
rect 24558 27234 24610 27246
rect 15710 27186 15762 27198
rect 12226 27134 12238 27186
rect 12290 27134 12302 27186
rect 13906 27134 13918 27186
rect 13970 27134 13982 27186
rect 15710 27122 15762 27134
rect 18510 27186 18562 27198
rect 18510 27122 18562 27134
rect 29374 27186 29426 27198
rect 38670 27186 38722 27198
rect 31714 27134 31726 27186
rect 31778 27134 31790 27186
rect 33842 27134 33854 27186
rect 33906 27134 33918 27186
rect 29374 27122 29426 27134
rect 38670 27122 38722 27134
rect 40014 27186 40066 27198
rect 41906 27134 41918 27186
rect 41970 27134 41982 27186
rect 58146 27134 58158 27186
rect 58210 27134 58222 27186
rect 40014 27122 40066 27134
rect 14702 27074 14754 27086
rect 6738 27022 6750 27074
rect 6802 27022 6814 27074
rect 7410 27022 7422 27074
rect 7474 27022 7486 27074
rect 9314 27022 9326 27074
rect 9378 27022 9390 27074
rect 10994 27022 11006 27074
rect 11058 27022 11070 27074
rect 11554 27022 11566 27074
rect 11618 27022 11630 27074
rect 14702 27010 14754 27022
rect 15262 27074 15314 27086
rect 15262 27010 15314 27022
rect 25902 27074 25954 27086
rect 25902 27010 25954 27022
rect 26126 27074 26178 27086
rect 26126 27010 26178 27022
rect 26798 27074 26850 27086
rect 26798 27010 26850 27022
rect 28030 27074 28082 27086
rect 28030 27010 28082 27022
rect 30606 27074 30658 27086
rect 45054 27074 45106 27086
rect 30930 27022 30942 27074
rect 30994 27022 31006 27074
rect 37986 27022 37998 27074
rect 38050 27022 38062 27074
rect 40898 27022 40910 27074
rect 40962 27022 40974 27074
rect 30606 27010 30658 27022
rect 45054 27010 45106 27022
rect 52558 27074 52610 27086
rect 52558 27010 52610 27022
rect 53230 27074 53282 27086
rect 53230 27010 53282 27022
rect 53790 27074 53842 27086
rect 55346 27022 55358 27074
rect 55410 27022 55422 27074
rect 53790 27010 53842 27022
rect 13470 26962 13522 26974
rect 15150 26962 15202 26974
rect 6962 26910 6974 26962
rect 7026 26910 7038 26962
rect 10098 26910 10110 26962
rect 10162 26910 10174 26962
rect 14354 26910 14366 26962
rect 14418 26910 14430 26962
rect 13470 26898 13522 26910
rect 15150 26898 15202 26910
rect 24670 26962 24722 26974
rect 24670 26898 24722 26910
rect 25678 26962 25730 26974
rect 25678 26898 25730 26910
rect 26462 26962 26514 26974
rect 44270 26962 44322 26974
rect 38210 26910 38222 26962
rect 38274 26910 38286 26962
rect 26462 26898 26514 26910
rect 44270 26898 44322 26910
rect 44830 26962 44882 26974
rect 44830 26898 44882 26910
rect 45390 26962 45442 26974
rect 45390 26898 45442 26910
rect 52782 26962 52834 26974
rect 52782 26898 52834 26910
rect 53006 26962 53058 26974
rect 53006 26898 53058 26910
rect 53454 26962 53506 26974
rect 56018 26910 56030 26962
rect 56082 26910 56094 26962
rect 53454 26898 53506 26910
rect 14926 26850 14978 26862
rect 24558 26850 24610 26862
rect 18162 26798 18174 26850
rect 18226 26847 18238 26850
rect 18386 26847 18398 26850
rect 18226 26801 18398 26847
rect 18226 26798 18238 26801
rect 18386 26798 18398 26801
rect 18450 26798 18462 26850
rect 14926 26786 14978 26798
rect 24558 26786 24610 26798
rect 25454 26850 25506 26862
rect 25454 26786 25506 26798
rect 25566 26850 25618 26862
rect 25566 26786 25618 26798
rect 26574 26850 26626 26862
rect 26574 26786 26626 26798
rect 27806 26850 27858 26862
rect 29822 26850 29874 26862
rect 28354 26798 28366 26850
rect 28418 26798 28430 26850
rect 27806 26786 27858 26798
rect 29822 26786 29874 26798
rect 43934 26850 43986 26862
rect 43934 26786 43986 26798
rect 44158 26850 44210 26862
rect 44158 26786 44210 26798
rect 44942 26850 44994 26862
rect 44942 26786 44994 26798
rect 53678 26850 53730 26862
rect 53678 26786 53730 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 9550 26514 9602 26526
rect 9550 26450 9602 26462
rect 10670 26514 10722 26526
rect 10670 26450 10722 26462
rect 11566 26514 11618 26526
rect 11566 26450 11618 26462
rect 11790 26514 11842 26526
rect 15934 26514 15986 26526
rect 15586 26462 15598 26514
rect 15650 26462 15662 26514
rect 11790 26450 11842 26462
rect 15934 26450 15986 26462
rect 18174 26514 18226 26526
rect 18174 26450 18226 26462
rect 25118 26514 25170 26526
rect 25118 26450 25170 26462
rect 25342 26514 25394 26526
rect 25342 26450 25394 26462
rect 26462 26514 26514 26526
rect 26462 26450 26514 26462
rect 27358 26514 27410 26526
rect 27358 26450 27410 26462
rect 28478 26514 28530 26526
rect 28478 26450 28530 26462
rect 29038 26514 29090 26526
rect 29038 26450 29090 26462
rect 30270 26514 30322 26526
rect 30270 26450 30322 26462
rect 30830 26514 30882 26526
rect 30830 26450 30882 26462
rect 34414 26514 34466 26526
rect 34414 26450 34466 26462
rect 37662 26514 37714 26526
rect 37662 26450 37714 26462
rect 39230 26514 39282 26526
rect 39230 26450 39282 26462
rect 40126 26514 40178 26526
rect 40126 26450 40178 26462
rect 41918 26514 41970 26526
rect 41918 26450 41970 26462
rect 52334 26514 52386 26526
rect 52334 26450 52386 26462
rect 57038 26514 57090 26526
rect 57038 26450 57090 26462
rect 12350 26402 12402 26414
rect 18062 26402 18114 26414
rect 16482 26350 16494 26402
rect 16546 26350 16558 26402
rect 17378 26350 17390 26402
rect 17442 26350 17454 26402
rect 12350 26338 12402 26350
rect 18062 26338 18114 26350
rect 18622 26402 18674 26414
rect 18622 26338 18674 26350
rect 25454 26402 25506 26414
rect 25454 26338 25506 26350
rect 28814 26402 28866 26414
rect 28814 26338 28866 26350
rect 29598 26402 29650 26414
rect 29598 26338 29650 26350
rect 33966 26402 34018 26414
rect 41470 26402 41522 26414
rect 39778 26350 39790 26402
rect 39842 26350 39854 26402
rect 33966 26338 34018 26350
rect 41470 26338 41522 26350
rect 52558 26402 52610 26414
rect 52558 26338 52610 26350
rect 52670 26402 52722 26414
rect 52670 26338 52722 26350
rect 10446 26290 10498 26302
rect 8754 26238 8766 26290
rect 8818 26238 8830 26290
rect 10446 26226 10498 26238
rect 11118 26290 11170 26302
rect 16830 26290 16882 26302
rect 13234 26238 13246 26290
rect 13298 26238 13310 26290
rect 11118 26226 11170 26238
rect 16830 26226 16882 26238
rect 17726 26290 17778 26302
rect 17726 26226 17778 26238
rect 19182 26290 19234 26302
rect 26126 26290 26178 26302
rect 22754 26238 22766 26290
rect 22818 26238 22830 26290
rect 23762 26238 23774 26290
rect 23826 26238 23838 26290
rect 19182 26226 19234 26238
rect 26126 26226 26178 26238
rect 26350 26290 26402 26302
rect 26350 26226 26402 26238
rect 26574 26290 26626 26302
rect 26574 26226 26626 26238
rect 27134 26290 27186 26302
rect 28254 26290 28306 26302
rect 27458 26238 27470 26290
rect 27522 26238 27534 26290
rect 27134 26226 27186 26238
rect 28254 26226 28306 26238
rect 28590 26290 28642 26302
rect 28590 26226 28642 26238
rect 29150 26290 29202 26302
rect 29150 26226 29202 26238
rect 30158 26290 30210 26302
rect 41134 26290 41186 26302
rect 48190 26290 48242 26302
rect 39442 26238 39454 26290
rect 39506 26238 39518 26290
rect 42578 26238 42590 26290
rect 42642 26238 42654 26290
rect 47618 26238 47630 26290
rect 47682 26238 47694 26290
rect 30158 26226 30210 26238
rect 41134 26226 41186 26238
rect 48190 26226 48242 26238
rect 56590 26290 56642 26302
rect 56590 26226 56642 26238
rect 56926 26290 56978 26302
rect 56926 26226 56978 26238
rect 57262 26290 57314 26302
rect 57262 26226 57314 26238
rect 10558 26178 10610 26190
rect 22318 26178 22370 26190
rect 5618 26126 5630 26178
rect 5682 26126 5694 26178
rect 7858 26126 7870 26178
rect 7922 26126 7934 26178
rect 9986 26126 9998 26178
rect 10050 26126 10062 26178
rect 15026 26126 15038 26178
rect 15090 26126 15102 26178
rect 10558 26114 10610 26126
rect 22318 26114 22370 26126
rect 23214 26178 23266 26190
rect 23214 26114 23266 26126
rect 24110 26178 24162 26190
rect 24110 26114 24162 26126
rect 24334 26178 24386 26190
rect 24334 26114 24386 26126
rect 27246 26178 27298 26190
rect 27246 26114 27298 26126
rect 36766 26178 36818 26190
rect 58158 26178 58210 26190
rect 43250 26126 43262 26178
rect 43314 26126 43326 26178
rect 45378 26126 45390 26178
rect 45442 26126 45454 26178
rect 36766 26114 36818 26126
rect 58158 26114 58210 26126
rect 18174 26066 18226 26078
rect 18174 26002 18226 26014
rect 25902 26066 25954 26078
rect 25902 26002 25954 26014
rect 27806 26066 27858 26078
rect 27806 26002 27858 26014
rect 29486 26066 29538 26078
rect 29486 26002 29538 26014
rect 30270 26066 30322 26078
rect 30270 26002 30322 26014
rect 33854 26066 33906 26078
rect 33854 26002 33906 26014
rect 39118 26066 39170 26078
rect 39118 26002 39170 26014
rect 41022 26066 41074 26078
rect 41022 26002 41074 26014
rect 41358 26066 41410 26078
rect 41358 26002 41410 26014
rect 47294 26066 47346 26078
rect 47294 26002 47346 26014
rect 47630 26066 47682 26078
rect 47630 26002 47682 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 24110 25730 24162 25742
rect 24110 25666 24162 25678
rect 33182 25730 33234 25742
rect 33182 25666 33234 25678
rect 39790 25730 39842 25742
rect 39790 25666 39842 25678
rect 39902 25730 39954 25742
rect 39902 25666 39954 25678
rect 40686 25730 40738 25742
rect 40686 25666 40738 25678
rect 43598 25730 43650 25742
rect 43598 25666 43650 25678
rect 43934 25730 43986 25742
rect 43934 25666 43986 25678
rect 44046 25730 44098 25742
rect 44046 25666 44098 25678
rect 23326 25618 23378 25630
rect 11554 25566 11566 25618
rect 11618 25566 11630 25618
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 15810 25566 15822 25618
rect 15874 25566 15886 25618
rect 19954 25566 19966 25618
rect 20018 25566 20030 25618
rect 23326 25554 23378 25566
rect 26126 25618 26178 25630
rect 27694 25618 27746 25630
rect 26674 25566 26686 25618
rect 26738 25566 26750 25618
rect 26126 25554 26178 25566
rect 27694 25554 27746 25566
rect 28590 25618 28642 25630
rect 28590 25554 28642 25566
rect 33854 25618 33906 25630
rect 33854 25554 33906 25566
rect 34190 25618 34242 25630
rect 34190 25554 34242 25566
rect 36206 25618 36258 25630
rect 36206 25554 36258 25566
rect 39006 25618 39058 25630
rect 39006 25554 39058 25566
rect 39342 25618 39394 25630
rect 50318 25618 50370 25630
rect 45154 25566 45166 25618
rect 45218 25566 45230 25618
rect 46946 25566 46958 25618
rect 47010 25566 47022 25618
rect 49074 25566 49086 25618
rect 49138 25566 49150 25618
rect 39342 25554 39394 25566
rect 50318 25554 50370 25566
rect 7646 25506 7698 25518
rect 7646 25442 7698 25454
rect 7982 25506 8034 25518
rect 7982 25442 8034 25454
rect 8206 25506 8258 25518
rect 12126 25506 12178 25518
rect 14702 25506 14754 25518
rect 8642 25454 8654 25506
rect 8706 25454 8718 25506
rect 14018 25454 14030 25506
rect 14082 25454 14094 25506
rect 8206 25442 8258 25454
rect 12126 25442 12178 25454
rect 14702 25442 14754 25454
rect 16606 25506 16658 25518
rect 24222 25506 24274 25518
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 16606 25442 16658 25454
rect 24222 25442 24274 25454
rect 24558 25506 24610 25518
rect 24558 25442 24610 25454
rect 25566 25506 25618 25518
rect 26014 25506 26066 25518
rect 25890 25454 25902 25506
rect 25954 25454 25966 25506
rect 25566 25442 25618 25454
rect 26014 25442 26066 25454
rect 26238 25506 26290 25518
rect 27806 25506 27858 25518
rect 32398 25506 32450 25518
rect 26898 25454 26910 25506
rect 26962 25454 26974 25506
rect 29698 25454 29710 25506
rect 29762 25454 29774 25506
rect 26238 25442 26290 25454
rect 27806 25442 27858 25454
rect 32398 25442 32450 25454
rect 32734 25506 32786 25518
rect 32734 25442 32786 25454
rect 33294 25506 33346 25518
rect 33294 25442 33346 25454
rect 34974 25506 35026 25518
rect 34974 25442 35026 25454
rect 35758 25506 35810 25518
rect 35758 25442 35810 25454
rect 36990 25506 37042 25518
rect 36990 25442 37042 25454
rect 38446 25506 38498 25518
rect 38446 25442 38498 25454
rect 40126 25506 40178 25518
rect 43710 25506 43762 25518
rect 45726 25506 45778 25518
rect 46622 25506 46674 25518
rect 52558 25506 52610 25518
rect 41906 25454 41918 25506
rect 41970 25454 41982 25506
rect 45042 25454 45054 25506
rect 45106 25454 45118 25506
rect 45938 25454 45950 25506
rect 46002 25454 46014 25506
rect 49858 25454 49870 25506
rect 49922 25454 49934 25506
rect 40126 25442 40178 25454
rect 43710 25442 43762 25454
rect 45726 25442 45778 25454
rect 46622 25442 46674 25454
rect 52558 25442 52610 25454
rect 53006 25506 53058 25518
rect 53006 25442 53058 25454
rect 53454 25506 53506 25518
rect 53454 25442 53506 25454
rect 53790 25506 53842 25518
rect 53790 25442 53842 25454
rect 56702 25506 56754 25518
rect 56702 25442 56754 25454
rect 14366 25394 14418 25406
rect 16270 25394 16322 25406
rect 21422 25394 21474 25406
rect 9314 25342 9326 25394
rect 9378 25342 9390 25394
rect 16034 25342 16046 25394
rect 16098 25342 16110 25394
rect 17714 25342 17726 25394
rect 17778 25342 17790 25394
rect 14366 25330 14418 25342
rect 16270 25330 16322 25342
rect 21422 25330 21474 25342
rect 21758 25394 21810 25406
rect 21758 25330 21810 25342
rect 21982 25394 22034 25406
rect 21982 25330 22034 25342
rect 24110 25394 24162 25406
rect 24110 25330 24162 25342
rect 24670 25394 24722 25406
rect 32622 25394 32674 25406
rect 37326 25394 37378 25406
rect 27346 25342 27358 25394
rect 27410 25342 27422 25394
rect 29474 25342 29486 25394
rect 29538 25342 29550 25394
rect 29810 25342 29822 25394
rect 29874 25342 29886 25394
rect 30930 25342 30942 25394
rect 30994 25342 31006 25394
rect 34626 25342 34638 25394
rect 34690 25342 34702 25394
rect 35410 25342 35422 25394
rect 35474 25342 35486 25394
rect 24670 25330 24722 25342
rect 32622 25330 32674 25342
rect 37326 25330 37378 25342
rect 37550 25394 37602 25406
rect 37550 25330 37602 25342
rect 38334 25394 38386 25406
rect 38334 25330 38386 25342
rect 39230 25394 39282 25406
rect 39230 25330 39282 25342
rect 40238 25394 40290 25406
rect 40238 25330 40290 25342
rect 40574 25394 40626 25406
rect 40574 25330 40626 25342
rect 40686 25394 40738 25406
rect 40686 25330 40738 25342
rect 42478 25394 42530 25406
rect 42478 25330 42530 25342
rect 44830 25394 44882 25406
rect 44830 25330 44882 25342
rect 45278 25394 45330 25406
rect 45278 25330 45330 25342
rect 53230 25394 53282 25406
rect 53230 25330 53282 25342
rect 53678 25394 53730 25406
rect 53678 25330 53730 25342
rect 56590 25394 56642 25406
rect 56590 25330 56642 25342
rect 58158 25394 58210 25406
rect 58158 25330 58210 25342
rect 7870 25282 7922 25294
rect 7870 25218 7922 25230
rect 12238 25282 12290 25294
rect 12238 25218 12290 25230
rect 12462 25282 12514 25294
rect 12462 25218 12514 25230
rect 12798 25282 12850 25294
rect 12798 25218 12850 25230
rect 13582 25282 13634 25294
rect 13582 25218 13634 25230
rect 14478 25282 14530 25294
rect 14478 25218 14530 25230
rect 15598 25282 15650 25294
rect 15598 25218 15650 25230
rect 16382 25282 16434 25294
rect 16382 25218 16434 25230
rect 21534 25282 21586 25294
rect 21534 25218 21586 25230
rect 22542 25282 22594 25294
rect 22542 25218 22594 25230
rect 31278 25282 31330 25294
rect 31278 25218 31330 25230
rect 33182 25282 33234 25294
rect 33182 25218 33234 25230
rect 34078 25282 34130 25294
rect 34078 25218 34130 25230
rect 37102 25282 37154 25294
rect 37102 25218 37154 25230
rect 37998 25282 38050 25294
rect 37998 25218 38050 25230
rect 38222 25282 38274 25294
rect 38222 25218 38274 25230
rect 41470 25282 41522 25294
rect 42926 25282 42978 25294
rect 41682 25230 41694 25282
rect 41746 25230 41758 25282
rect 41470 25218 41522 25230
rect 42926 25218 42978 25230
rect 52782 25282 52834 25294
rect 52782 25218 52834 25230
rect 56366 25282 56418 25294
rect 56366 25218 56418 25230
rect 57598 25282 57650 25294
rect 57598 25218 57650 25230
rect 57822 25282 57874 25294
rect 57822 25218 57874 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 8430 24946 8482 24958
rect 8430 24882 8482 24894
rect 8878 24946 8930 24958
rect 8878 24882 8930 24894
rect 13470 24946 13522 24958
rect 13470 24882 13522 24894
rect 14702 24946 14754 24958
rect 14702 24882 14754 24894
rect 15150 24946 15202 24958
rect 15150 24882 15202 24894
rect 16158 24946 16210 24958
rect 16158 24882 16210 24894
rect 16270 24946 16322 24958
rect 16270 24882 16322 24894
rect 17390 24946 17442 24958
rect 17390 24882 17442 24894
rect 19182 24946 19234 24958
rect 19182 24882 19234 24894
rect 25566 24946 25618 24958
rect 25566 24882 25618 24894
rect 26126 24946 26178 24958
rect 26126 24882 26178 24894
rect 27134 24946 27186 24958
rect 27134 24882 27186 24894
rect 28142 24946 28194 24958
rect 28142 24882 28194 24894
rect 29934 24946 29986 24958
rect 29934 24882 29986 24894
rect 31390 24946 31442 24958
rect 31390 24882 31442 24894
rect 39230 24946 39282 24958
rect 39230 24882 39282 24894
rect 45838 24946 45890 24958
rect 45838 24882 45890 24894
rect 46174 24946 46226 24958
rect 46174 24882 46226 24894
rect 52558 24946 52610 24958
rect 52558 24882 52610 24894
rect 56814 24946 56866 24958
rect 56814 24882 56866 24894
rect 14478 24834 14530 24846
rect 14478 24770 14530 24782
rect 16494 24834 16546 24846
rect 16494 24770 16546 24782
rect 16606 24834 16658 24846
rect 16606 24770 16658 24782
rect 17614 24834 17666 24846
rect 25342 24834 25394 24846
rect 20514 24782 20526 24834
rect 20578 24782 20590 24834
rect 17614 24770 17666 24782
rect 25342 24770 25394 24782
rect 25902 24834 25954 24846
rect 25902 24770 25954 24782
rect 27694 24834 27746 24846
rect 27694 24770 27746 24782
rect 28926 24834 28978 24846
rect 40910 24834 40962 24846
rect 36082 24782 36094 24834
rect 36146 24782 36158 24834
rect 28926 24770 28978 24782
rect 40910 24770 40962 24782
rect 41134 24834 41186 24846
rect 41134 24770 41186 24782
rect 42142 24834 42194 24846
rect 52782 24834 52834 24846
rect 50194 24782 50206 24834
rect 50258 24782 50270 24834
rect 42142 24770 42194 24782
rect 52782 24770 52834 24782
rect 57822 24834 57874 24846
rect 57822 24770 57874 24782
rect 25230 24722 25282 24734
rect 10210 24670 10222 24722
rect 10274 24670 10286 24722
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 14242 24670 14254 24722
rect 14306 24670 14318 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 18162 24670 18174 24722
rect 18226 24670 18238 24722
rect 19730 24670 19742 24722
rect 19794 24670 19806 24722
rect 23426 24670 23438 24722
rect 23490 24670 23502 24722
rect 25230 24658 25282 24670
rect 25790 24722 25842 24734
rect 25790 24658 25842 24670
rect 27470 24722 27522 24734
rect 27470 24658 27522 24670
rect 28702 24722 28754 24734
rect 32958 24722 33010 24734
rect 29138 24670 29150 24722
rect 29202 24670 29214 24722
rect 29474 24670 29486 24722
rect 29538 24670 29550 24722
rect 28702 24658 28754 24670
rect 32958 24658 33010 24670
rect 33294 24722 33346 24734
rect 41806 24722 41858 24734
rect 33618 24670 33630 24722
rect 33682 24670 33694 24722
rect 34178 24670 34190 24722
rect 34242 24670 34254 24722
rect 35410 24670 35422 24722
rect 35474 24670 35486 24722
rect 33294 24658 33346 24670
rect 41806 24658 41858 24670
rect 42702 24722 42754 24734
rect 52894 24722 52946 24734
rect 43138 24670 43150 24722
rect 43202 24670 43214 24722
rect 49522 24670 49534 24722
rect 49586 24670 49598 24722
rect 42702 24658 42754 24670
rect 52894 24658 52946 24670
rect 56478 24722 56530 24734
rect 56478 24658 56530 24670
rect 56926 24722 56978 24734
rect 56926 24658 56978 24670
rect 57150 24722 57202 24734
rect 57150 24658 57202 24670
rect 15598 24610 15650 24622
rect 18622 24610 18674 24622
rect 23998 24610 24050 24622
rect 38670 24610 38722 24622
rect 10882 24558 10894 24610
rect 10946 24558 10958 24610
rect 13010 24558 13022 24610
rect 13074 24558 13086 24610
rect 14354 24558 14366 24610
rect 14418 24558 14430 24610
rect 17714 24558 17726 24610
rect 17778 24558 17790 24610
rect 22642 24558 22654 24610
rect 22706 24558 22718 24610
rect 23090 24558 23102 24610
rect 23154 24558 23166 24610
rect 29026 24558 29038 24610
rect 29090 24558 29102 24610
rect 31826 24558 31838 24610
rect 31890 24558 31902 24610
rect 38210 24558 38222 24610
rect 38274 24558 38286 24610
rect 15598 24546 15650 24558
rect 18622 24546 18674 24558
rect 23998 24546 24050 24558
rect 38670 24546 38722 24558
rect 41022 24610 41074 24622
rect 41022 24546 41074 24558
rect 43598 24610 43650 24622
rect 43598 24546 43650 24558
rect 44382 24610 44434 24622
rect 44382 24546 44434 24558
rect 44830 24610 44882 24622
rect 44830 24546 44882 24558
rect 45278 24610 45330 24622
rect 53342 24610 53394 24622
rect 52322 24558 52334 24610
rect 52386 24558 52398 24610
rect 57474 24558 57486 24610
rect 57538 24558 57550 24610
rect 45278 24546 45330 24558
rect 53342 24546 53394 24558
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 31502 24162 31554 24174
rect 31502 24098 31554 24110
rect 19406 24050 19458 24062
rect 19406 23986 19458 23998
rect 22318 24050 22370 24062
rect 22318 23986 22370 23998
rect 27694 24050 27746 24062
rect 27694 23986 27746 23998
rect 29150 24050 29202 24062
rect 29150 23986 29202 23998
rect 38446 24050 38498 24062
rect 55122 23998 55134 24050
rect 55186 23998 55198 24050
rect 57250 23998 57262 24050
rect 57314 23998 57326 24050
rect 38446 23986 38498 23998
rect 20302 23938 20354 23950
rect 18946 23886 18958 23938
rect 19010 23886 19022 23938
rect 19842 23886 19854 23938
rect 19906 23886 19918 23938
rect 20302 23874 20354 23886
rect 22206 23938 22258 23950
rect 22206 23874 22258 23886
rect 22878 23938 22930 23950
rect 45502 23938 45554 23950
rect 52670 23938 52722 23950
rect 24882 23886 24894 23938
rect 24946 23886 24958 23938
rect 26898 23886 26910 23938
rect 26962 23886 26974 23938
rect 28018 23886 28030 23938
rect 28082 23886 28094 23938
rect 33730 23886 33742 23938
rect 33794 23886 33806 23938
rect 35746 23886 35758 23938
rect 35810 23886 35822 23938
rect 46162 23886 46174 23938
rect 46226 23886 46238 23938
rect 22878 23874 22930 23886
rect 45502 23874 45554 23886
rect 52670 23874 52722 23886
rect 53230 23938 53282 23950
rect 53230 23874 53282 23886
rect 53790 23938 53842 23950
rect 53790 23874 53842 23886
rect 54126 23938 54178 23950
rect 54126 23874 54178 23886
rect 54462 23938 54514 23950
rect 58034 23886 58046 23938
rect 58098 23886 58110 23938
rect 54462 23874 54514 23886
rect 24334 23826 24386 23838
rect 24334 23762 24386 23774
rect 26350 23826 26402 23838
rect 31614 23826 31666 23838
rect 52894 23826 52946 23838
rect 28242 23774 28254 23826
rect 28306 23774 28318 23826
rect 35970 23774 35982 23826
rect 36034 23774 36046 23826
rect 26350 23762 26402 23774
rect 31614 23762 31666 23774
rect 52894 23762 52946 23774
rect 53454 23826 53506 23838
rect 53454 23762 53506 23774
rect 53678 23826 53730 23838
rect 53678 23762 53730 23774
rect 16606 23714 16658 23726
rect 16606 23650 16658 23662
rect 20750 23714 20802 23726
rect 20750 23650 20802 23662
rect 21982 23714 22034 23726
rect 21982 23650 22034 23662
rect 22430 23714 22482 23726
rect 29262 23714 29314 23726
rect 26786 23662 26798 23714
rect 26850 23662 26862 23714
rect 22430 23650 22482 23662
rect 29262 23650 29314 23662
rect 32062 23714 32114 23726
rect 44942 23714 44994 23726
rect 46510 23714 46562 23726
rect 33506 23662 33518 23714
rect 33570 23662 33582 23714
rect 45826 23662 45838 23714
rect 45890 23662 45902 23714
rect 32062 23650 32114 23662
rect 44942 23650 44994 23662
rect 46510 23650 46562 23662
rect 46622 23714 46674 23726
rect 46622 23650 46674 23662
rect 46734 23714 46786 23726
rect 46734 23650 46786 23662
rect 53006 23714 53058 23726
rect 53006 23650 53058 23662
rect 54238 23714 54290 23726
rect 54238 23650 54290 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 19630 23378 19682 23390
rect 19630 23314 19682 23326
rect 23438 23378 23490 23390
rect 23438 23314 23490 23326
rect 24334 23378 24386 23390
rect 24334 23314 24386 23326
rect 25342 23378 25394 23390
rect 25342 23314 25394 23326
rect 27582 23378 27634 23390
rect 27582 23314 27634 23326
rect 42142 23378 42194 23390
rect 42142 23314 42194 23326
rect 42478 23378 42530 23390
rect 42478 23314 42530 23326
rect 43150 23378 43202 23390
rect 43150 23314 43202 23326
rect 44158 23378 44210 23390
rect 44158 23314 44210 23326
rect 44606 23378 44658 23390
rect 44606 23314 44658 23326
rect 56702 23378 56754 23390
rect 56702 23314 56754 23326
rect 56926 23378 56978 23390
rect 56926 23314 56978 23326
rect 39230 23266 39282 23278
rect 54014 23266 54066 23278
rect 15922 23214 15934 23266
rect 15986 23214 15998 23266
rect 30034 23214 30046 23266
rect 30098 23214 30110 23266
rect 44930 23214 44942 23266
rect 44994 23214 45006 23266
rect 51426 23214 51438 23266
rect 51490 23214 51502 23266
rect 39230 23202 39282 23214
rect 54014 23202 54066 23214
rect 54126 23266 54178 23278
rect 54126 23202 54178 23214
rect 54350 23266 54402 23278
rect 54350 23202 54402 23214
rect 56590 23266 56642 23278
rect 56590 23202 56642 23214
rect 22318 23154 22370 23166
rect 16706 23102 16718 23154
rect 16770 23102 16782 23154
rect 22318 23090 22370 23102
rect 22654 23154 22706 23166
rect 22654 23090 22706 23102
rect 22990 23154 23042 23166
rect 22990 23090 23042 23102
rect 23662 23154 23714 23166
rect 23662 23090 23714 23102
rect 24110 23154 24162 23166
rect 24110 23090 24162 23102
rect 24222 23154 24274 23166
rect 24222 23090 24274 23102
rect 25230 23154 25282 23166
rect 33630 23154 33682 23166
rect 30706 23102 30718 23154
rect 30770 23102 30782 23154
rect 25230 23090 25282 23102
rect 33630 23090 33682 23102
rect 34078 23154 34130 23166
rect 34078 23090 34130 23102
rect 38110 23154 38162 23166
rect 38110 23090 38162 23102
rect 38558 23154 38610 23166
rect 38558 23090 38610 23102
rect 38782 23154 38834 23166
rect 38782 23090 38834 23102
rect 41022 23154 41074 23166
rect 41022 23090 41074 23102
rect 42030 23154 42082 23166
rect 42030 23090 42082 23102
rect 42254 23154 42306 23166
rect 45378 23102 45390 23154
rect 45442 23102 45454 23154
rect 50754 23102 50766 23154
rect 50818 23102 50830 23154
rect 42254 23090 42306 23102
rect 17502 23042 17554 23054
rect 13794 22990 13806 23042
rect 13858 22990 13870 23042
rect 17502 22978 17554 22990
rect 22542 23042 22594 23054
rect 33070 23042 33122 23054
rect 27906 22990 27918 23042
rect 27970 22990 27982 23042
rect 22542 22978 22594 22990
rect 33070 22978 33122 22990
rect 38334 23042 38386 23054
rect 54686 23042 54738 23054
rect 43698 22990 43710 23042
rect 43762 22990 43774 23042
rect 46050 22990 46062 23042
rect 46114 22990 46126 23042
rect 48178 22990 48190 23042
rect 48242 22990 48254 23042
rect 53554 22990 53566 23042
rect 53618 22990 53630 23042
rect 38334 22978 38386 22990
rect 54686 22978 54738 22990
rect 58158 23042 58210 23054
rect 58158 22978 58210 22990
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 33182 22482 33234 22494
rect 45054 22482 45106 22494
rect 36418 22430 36430 22482
rect 36482 22430 36494 22482
rect 40674 22430 40686 22482
rect 40738 22430 40750 22482
rect 44146 22430 44158 22482
rect 44210 22430 44222 22482
rect 33182 22418 33234 22430
rect 45054 22418 45106 22430
rect 45502 22482 45554 22494
rect 45502 22418 45554 22430
rect 45838 22482 45890 22494
rect 51214 22482 51266 22494
rect 47506 22430 47518 22482
rect 47570 22430 47582 22482
rect 50754 22430 50766 22482
rect 50818 22430 50830 22482
rect 45838 22418 45890 22430
rect 51214 22418 51266 22430
rect 24446 22370 24498 22382
rect 24446 22306 24498 22318
rect 26462 22370 26514 22382
rect 26462 22306 26514 22318
rect 26910 22370 26962 22382
rect 45614 22370 45666 22382
rect 33506 22318 33518 22370
rect 33570 22318 33582 22370
rect 37874 22318 37886 22370
rect 37938 22318 37950 22370
rect 38546 22318 38558 22370
rect 38610 22318 38622 22370
rect 41234 22318 41246 22370
rect 41298 22318 41310 22370
rect 26910 22306 26962 22318
rect 45614 22306 45666 22318
rect 45950 22370 46002 22382
rect 45950 22306 46002 22318
rect 46286 22370 46338 22382
rect 46286 22306 46338 22318
rect 46734 22370 46786 22382
rect 54910 22370 54962 22382
rect 47954 22318 47966 22370
rect 48018 22318 48030 22370
rect 46734 22306 46786 22318
rect 54910 22306 54962 22318
rect 56814 22370 56866 22382
rect 56814 22306 56866 22318
rect 57374 22370 57426 22382
rect 57374 22306 57426 22318
rect 57934 22370 57986 22382
rect 57934 22306 57986 22318
rect 23886 22258 23938 22270
rect 23886 22194 23938 22206
rect 25342 22258 25394 22270
rect 25342 22194 25394 22206
rect 27918 22258 27970 22270
rect 37214 22258 37266 22270
rect 34290 22206 34302 22258
rect 34354 22206 34366 22258
rect 27918 22194 27970 22206
rect 37214 22194 37266 22206
rect 37326 22258 37378 22270
rect 37326 22194 37378 22206
rect 37438 22258 37490 22270
rect 47070 22258 47122 22270
rect 54574 22258 54626 22270
rect 42018 22206 42030 22258
rect 42082 22206 42094 22258
rect 47170 22206 47182 22258
rect 47234 22206 47246 22258
rect 48626 22206 48638 22258
rect 48690 22206 48702 22258
rect 37438 22194 37490 22206
rect 47070 22194 47122 22206
rect 54574 22194 54626 22206
rect 55134 22258 55186 22270
rect 55134 22194 55186 22206
rect 56702 22258 56754 22270
rect 56702 22194 56754 22206
rect 57038 22258 57090 22270
rect 57038 22194 57090 22206
rect 46958 22146 47010 22158
rect 28466 22094 28478 22146
rect 28530 22094 28542 22146
rect 46958 22082 47010 22094
rect 54686 22146 54738 22158
rect 54686 22082 54738 22094
rect 56478 22146 56530 22158
rect 56478 22082 56530 22094
rect 57262 22146 57314 22158
rect 57262 22082 57314 22094
rect 57598 22146 57650 22158
rect 57598 22082 57650 22094
rect 57822 22146 57874 22158
rect 57822 22082 57874 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 18622 21810 18674 21822
rect 18622 21746 18674 21758
rect 19294 21810 19346 21822
rect 19294 21746 19346 21758
rect 19966 21810 20018 21822
rect 33630 21810 33682 21822
rect 25330 21758 25342 21810
rect 25394 21758 25406 21810
rect 19966 21746 20018 21758
rect 33630 21746 33682 21758
rect 34414 21810 34466 21822
rect 34414 21746 34466 21758
rect 35534 21810 35586 21822
rect 35534 21746 35586 21758
rect 36766 21810 36818 21822
rect 36766 21746 36818 21758
rect 40350 21810 40402 21822
rect 40350 21746 40402 21758
rect 41470 21810 41522 21822
rect 41470 21746 41522 21758
rect 46398 21810 46450 21822
rect 46398 21746 46450 21758
rect 47070 21810 47122 21822
rect 47070 21746 47122 21758
rect 47294 21810 47346 21822
rect 47294 21746 47346 21758
rect 49646 21810 49698 21822
rect 49646 21746 49698 21758
rect 26350 21698 26402 21710
rect 18274 21646 18286 21698
rect 18338 21646 18350 21698
rect 18946 21646 18958 21698
rect 19010 21646 19022 21698
rect 19618 21646 19630 21698
rect 19682 21646 19694 21698
rect 22418 21646 22430 21698
rect 22482 21646 22494 21698
rect 26350 21634 26402 21646
rect 27806 21698 27858 21710
rect 35758 21698 35810 21710
rect 38110 21698 38162 21710
rect 33954 21646 33966 21698
rect 34018 21646 34030 21698
rect 36082 21646 36094 21698
rect 36146 21646 36158 21698
rect 37090 21646 37102 21698
rect 37154 21646 37166 21698
rect 27806 21634 27858 21646
rect 35758 21634 35810 21646
rect 38110 21634 38162 21646
rect 41582 21698 41634 21710
rect 41582 21634 41634 21646
rect 41806 21698 41858 21710
rect 41806 21634 41858 21646
rect 49758 21698 49810 21710
rect 56926 21698 56978 21710
rect 54338 21646 54350 21698
rect 54402 21646 54414 21698
rect 49758 21634 49810 21646
rect 56926 21634 56978 21646
rect 57150 21698 57202 21710
rect 57150 21634 57202 21646
rect 34302 21586 34354 21598
rect 21746 21534 21758 21586
rect 21810 21534 21822 21586
rect 26786 21534 26798 21586
rect 26850 21534 26862 21586
rect 27234 21534 27246 21586
rect 27298 21534 27310 21586
rect 34302 21522 34354 21534
rect 34526 21586 34578 21598
rect 34526 21522 34578 21534
rect 34862 21586 34914 21598
rect 34862 21522 34914 21534
rect 35086 21586 35138 21598
rect 35086 21522 35138 21534
rect 35646 21586 35698 21598
rect 37774 21586 37826 21598
rect 36306 21534 36318 21586
rect 36370 21534 36382 21586
rect 35646 21522 35698 21534
rect 37774 21522 37826 21534
rect 38334 21586 38386 21598
rect 41134 21586 41186 21598
rect 38994 21534 39006 21586
rect 39058 21534 39070 21586
rect 38334 21522 38386 21534
rect 41134 21522 41186 21534
rect 47406 21586 47458 21598
rect 55582 21586 55634 21598
rect 55122 21534 55134 21586
rect 55186 21534 55198 21586
rect 47406 21522 47458 21534
rect 55582 21522 55634 21534
rect 56478 21586 56530 21598
rect 56478 21522 56530 21534
rect 45390 21474 45442 21486
rect 24546 21422 24558 21474
rect 24610 21422 24622 21474
rect 45390 21410 45442 21422
rect 47854 21474 47906 21486
rect 56702 21474 56754 21486
rect 52210 21422 52222 21474
rect 52274 21422 52286 21474
rect 47854 21410 47906 21422
rect 56702 21410 56754 21422
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 19406 20914 19458 20926
rect 18050 20862 18062 20914
rect 18114 20862 18126 20914
rect 19406 20850 19458 20862
rect 22766 20914 22818 20926
rect 22766 20850 22818 20862
rect 24894 20914 24946 20926
rect 24894 20850 24946 20862
rect 29262 20914 29314 20926
rect 29262 20850 29314 20862
rect 30158 20914 30210 20926
rect 33506 20862 33518 20914
rect 33570 20862 33582 20914
rect 56018 20862 56030 20914
rect 56082 20862 56094 20914
rect 58146 20862 58158 20914
rect 58210 20862 58222 20914
rect 30158 20850 30210 20862
rect 18286 20802 18338 20814
rect 15250 20750 15262 20802
rect 15314 20750 15326 20802
rect 18286 20738 18338 20750
rect 18734 20802 18786 20814
rect 18734 20738 18786 20750
rect 18846 20802 18898 20814
rect 18846 20738 18898 20750
rect 20078 20802 20130 20814
rect 20078 20738 20130 20750
rect 20526 20802 20578 20814
rect 20526 20738 20578 20750
rect 22430 20802 22482 20814
rect 22430 20738 22482 20750
rect 27918 20802 27970 20814
rect 27918 20738 27970 20750
rect 29374 20802 29426 20814
rect 33966 20802 34018 20814
rect 30706 20750 30718 20802
rect 30770 20750 30782 20802
rect 55234 20750 55246 20802
rect 55298 20750 55310 20802
rect 29374 20738 29426 20750
rect 33966 20738 34018 20750
rect 18510 20690 18562 20702
rect 15922 20638 15934 20690
rect 15986 20638 15998 20690
rect 18510 20626 18562 20638
rect 20750 20690 20802 20702
rect 20750 20626 20802 20638
rect 21870 20690 21922 20702
rect 21870 20626 21922 20638
rect 29150 20690 29202 20702
rect 29150 20626 29202 20638
rect 29710 20690 29762 20702
rect 31378 20638 31390 20690
rect 31442 20638 31454 20690
rect 29710 20626 29762 20638
rect 14814 20578 14866 20590
rect 14814 20514 14866 20526
rect 20302 20578 20354 20590
rect 20302 20514 20354 20526
rect 21758 20578 21810 20590
rect 21758 20514 21810 20526
rect 21982 20578 22034 20590
rect 41582 20578 41634 20590
rect 28242 20526 28254 20578
rect 28306 20526 28318 20578
rect 21982 20514 22034 20526
rect 41582 20514 41634 20526
rect 47294 20578 47346 20590
rect 47294 20514 47346 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 18510 20242 18562 20254
rect 18510 20178 18562 20190
rect 31278 20242 31330 20254
rect 31278 20178 31330 20190
rect 37774 20242 37826 20254
rect 37774 20178 37826 20190
rect 58158 20242 58210 20254
rect 58158 20178 58210 20190
rect 18398 20130 18450 20142
rect 31614 20130 31666 20142
rect 20178 20078 20190 20130
rect 20242 20078 20254 20130
rect 26786 20078 26798 20130
rect 26850 20078 26862 20130
rect 27458 20078 27470 20130
rect 27522 20078 27534 20130
rect 28578 20078 28590 20130
rect 28642 20078 28654 20130
rect 18398 20066 18450 20078
rect 31614 20066 31666 20078
rect 32062 20130 32114 20142
rect 32062 20066 32114 20078
rect 32398 20130 32450 20142
rect 32398 20066 32450 20078
rect 40350 20130 40402 20142
rect 40350 20066 40402 20078
rect 41246 20130 41298 20142
rect 41246 20066 41298 20078
rect 46622 20130 46674 20142
rect 46622 20066 46674 20078
rect 47966 20130 48018 20142
rect 47966 20066 48018 20078
rect 18062 20018 18114 20030
rect 18062 19954 18114 19966
rect 18622 20018 18674 20030
rect 31054 20018 31106 20030
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 26562 19966 26574 20018
rect 26626 19966 26638 20018
rect 27234 19966 27246 20018
rect 27298 19966 27310 20018
rect 27906 19966 27918 20018
rect 27970 19966 27982 20018
rect 18622 19954 18674 19966
rect 31054 19954 31106 19966
rect 31390 20018 31442 20030
rect 31390 19954 31442 19966
rect 31950 20018 32002 20030
rect 31950 19954 32002 19966
rect 32174 20018 32226 20030
rect 32174 19954 32226 19966
rect 40910 20018 40962 20030
rect 40910 19954 40962 19966
rect 41470 20018 41522 20030
rect 46846 20018 46898 20030
rect 41794 19966 41806 20018
rect 41858 19966 41870 20018
rect 41470 19954 41522 19966
rect 46846 19954 46898 19966
rect 47070 20018 47122 20030
rect 47070 19954 47122 19966
rect 47518 20018 47570 20030
rect 47518 19954 47570 19966
rect 47742 20018 47794 20030
rect 47742 19954 47794 19966
rect 41022 19906 41074 19918
rect 46286 19906 46338 19918
rect 22306 19854 22318 19906
rect 22370 19854 22382 19906
rect 30706 19854 30718 19906
rect 30770 19854 30782 19906
rect 42578 19854 42590 19906
rect 42642 19854 42654 19906
rect 44706 19854 44718 19906
rect 44770 19854 44782 19906
rect 41022 19842 41074 19854
rect 46286 19842 46338 19854
rect 46734 19906 46786 19918
rect 46734 19842 46786 19854
rect 47630 19906 47682 19918
rect 47630 19842 47682 19854
rect 50318 19906 50370 19918
rect 50318 19842 50370 19854
rect 51214 19906 51266 19918
rect 51214 19842 51266 19854
rect 50082 19742 50094 19794
rect 50146 19791 50158 19794
rect 50306 19791 50318 19794
rect 50146 19745 50318 19791
rect 50146 19742 50158 19745
rect 50306 19742 50318 19745
rect 50370 19742 50382 19794
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 17726 19346 17778 19358
rect 17154 19294 17166 19346
rect 17218 19294 17230 19346
rect 17726 19282 17778 19294
rect 26238 19346 26290 19358
rect 26238 19282 26290 19294
rect 30046 19346 30098 19358
rect 30046 19282 30098 19294
rect 30942 19346 30994 19358
rect 39790 19346 39842 19358
rect 34178 19294 34190 19346
rect 34242 19294 34254 19346
rect 30942 19282 30994 19294
rect 39790 19282 39842 19294
rect 42142 19346 42194 19358
rect 47842 19294 47854 19346
rect 47906 19294 47918 19346
rect 49970 19294 49982 19346
rect 50034 19294 50046 19346
rect 42142 19282 42194 19294
rect 18286 19234 18338 19246
rect 14354 19182 14366 19234
rect 14418 19182 14430 19234
rect 18286 19170 18338 19182
rect 18958 19234 19010 19246
rect 18958 19170 19010 19182
rect 23662 19234 23714 19246
rect 23662 19170 23714 19182
rect 24334 19234 24386 19246
rect 24334 19170 24386 19182
rect 26574 19234 26626 19246
rect 26574 19170 26626 19182
rect 26798 19234 26850 19246
rect 26798 19170 26850 19182
rect 30606 19234 30658 19246
rect 30606 19170 30658 19182
rect 33742 19234 33794 19246
rect 33742 19170 33794 19182
rect 35422 19234 35474 19246
rect 35422 19170 35474 19182
rect 36990 19234 37042 19246
rect 36990 19170 37042 19182
rect 37214 19234 37266 19246
rect 37214 19170 37266 19182
rect 37550 19234 37602 19246
rect 37550 19170 37602 19182
rect 37998 19234 38050 19246
rect 37998 19170 38050 19182
rect 38782 19234 38834 19246
rect 38782 19170 38834 19182
rect 39118 19234 39170 19246
rect 39118 19170 39170 19182
rect 42254 19234 42306 19246
rect 42254 19170 42306 19182
rect 45614 19234 45666 19246
rect 45614 19170 45666 19182
rect 46174 19234 46226 19246
rect 50430 19234 50482 19246
rect 47170 19182 47182 19234
rect 47234 19182 47246 19234
rect 46174 19170 46226 19182
rect 50430 19170 50482 19182
rect 27134 19122 27186 19134
rect 15026 19070 15038 19122
rect 15090 19070 15102 19122
rect 27134 19058 27186 19070
rect 39342 19122 39394 19134
rect 39342 19058 39394 19070
rect 45950 19122 46002 19134
rect 45950 19058 46002 19070
rect 50878 19122 50930 19134
rect 50878 19058 50930 19070
rect 51102 19122 51154 19134
rect 51102 19058 51154 19070
rect 18398 19010 18450 19022
rect 18398 18946 18450 18958
rect 18510 19010 18562 19022
rect 18510 18946 18562 18958
rect 23998 19010 24050 19022
rect 23998 18946 24050 18958
rect 26686 19010 26738 19022
rect 26686 18946 26738 18958
rect 29934 19010 29986 19022
rect 29934 18946 29986 18958
rect 30158 19010 30210 19022
rect 30158 18946 30210 18958
rect 34638 19010 34690 19022
rect 35982 19010 36034 19022
rect 34962 18958 34974 19010
rect 35026 18958 35038 19010
rect 34638 18946 34690 18958
rect 35982 18946 36034 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 37886 19010 37938 19022
rect 37886 18946 37938 18958
rect 38110 19010 38162 19022
rect 38110 18946 38162 18958
rect 38334 19010 38386 19022
rect 38334 18946 38386 18958
rect 38894 19010 38946 19022
rect 38894 18946 38946 18958
rect 41806 19010 41858 19022
rect 41806 18946 41858 18958
rect 42030 19010 42082 19022
rect 42030 18946 42082 18958
rect 45278 19010 45330 19022
rect 45278 18946 45330 18958
rect 45838 19010 45890 19022
rect 45838 18946 45890 18958
rect 50766 19010 50818 19022
rect 50766 18946 50818 18958
rect 51438 19010 51490 19022
rect 51438 18946 51490 18958
rect 51550 19010 51602 19022
rect 51550 18946 51602 18958
rect 51662 19010 51714 19022
rect 51662 18946 51714 18958
rect 51886 19010 51938 19022
rect 51886 18946 51938 18958
rect 52782 19010 52834 19022
rect 52782 18946 52834 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 21758 18674 21810 18686
rect 21758 18610 21810 18622
rect 28478 18674 28530 18686
rect 39566 18674 39618 18686
rect 33842 18622 33854 18674
rect 33906 18622 33918 18674
rect 28478 18610 28530 18622
rect 39566 18610 39618 18622
rect 39678 18674 39730 18686
rect 39678 18610 39730 18622
rect 41246 18674 41298 18686
rect 41246 18610 41298 18622
rect 18510 18562 18562 18574
rect 28702 18562 28754 18574
rect 24434 18510 24446 18562
rect 24498 18510 24510 18562
rect 26002 18510 26014 18562
rect 26066 18510 26078 18562
rect 18510 18498 18562 18510
rect 28702 18498 28754 18510
rect 39790 18562 39842 18574
rect 39790 18498 39842 18510
rect 42142 18562 42194 18574
rect 52558 18562 52610 18574
rect 45826 18510 45838 18562
rect 45890 18510 45902 18562
rect 50866 18510 50878 18562
rect 50930 18510 50942 18562
rect 42142 18498 42194 18510
rect 52558 18498 52610 18510
rect 17950 18450 18002 18462
rect 17950 18386 18002 18398
rect 18062 18450 18114 18462
rect 18062 18386 18114 18398
rect 18286 18450 18338 18462
rect 18286 18386 18338 18398
rect 19070 18450 19122 18462
rect 19070 18386 19122 18398
rect 21982 18450 22034 18462
rect 21982 18386 22034 18398
rect 22430 18450 22482 18462
rect 22430 18386 22482 18398
rect 22990 18450 23042 18462
rect 22990 18386 23042 18398
rect 23214 18450 23266 18462
rect 28590 18450 28642 18462
rect 24210 18398 24222 18450
rect 24274 18398 24286 18450
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 23214 18386 23266 18398
rect 28590 18386 28642 18398
rect 29150 18450 29202 18462
rect 34190 18450 34242 18462
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 29150 18386 29202 18398
rect 34190 18386 34242 18398
rect 34750 18450 34802 18462
rect 40238 18450 40290 18462
rect 35298 18398 35310 18450
rect 35362 18398 35374 18450
rect 35970 18398 35982 18450
rect 36034 18398 36046 18450
rect 34750 18386 34802 18398
rect 40238 18386 40290 18398
rect 41358 18450 41410 18462
rect 41358 18386 41410 18398
rect 41470 18450 41522 18462
rect 42366 18450 42418 18462
rect 41794 18398 41806 18450
rect 41858 18398 41870 18450
rect 41470 18386 41522 18398
rect 42366 18386 42418 18398
rect 42590 18450 42642 18462
rect 42590 18386 42642 18398
rect 43150 18450 43202 18462
rect 43150 18386 43202 18398
rect 43934 18450 43986 18462
rect 43934 18386 43986 18398
rect 44494 18450 44546 18462
rect 52222 18450 52274 18462
rect 53118 18450 53170 18462
rect 45042 18398 45054 18450
rect 45106 18398 45118 18450
rect 50418 18398 50430 18450
rect 50482 18398 50494 18450
rect 51314 18398 51326 18450
rect 51378 18398 51390 18450
rect 52882 18398 52894 18450
rect 52946 18398 52958 18450
rect 44494 18386 44546 18398
rect 52222 18386 52274 18398
rect 53118 18386 53170 18398
rect 21870 18338 21922 18350
rect 21870 18274 21922 18286
rect 23774 18338 23826 18350
rect 31390 18338 31442 18350
rect 38558 18338 38610 18350
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 38098 18286 38110 18338
rect 38162 18286 38174 18338
rect 23774 18274 23826 18286
rect 31390 18274 31442 18286
rect 38558 18274 38610 18286
rect 42254 18338 42306 18350
rect 42254 18274 42306 18286
rect 43598 18338 43650 18350
rect 53566 18338 53618 18350
rect 47954 18286 47966 18338
rect 48018 18286 48030 18338
rect 51090 18286 51102 18338
rect 51154 18286 51166 18338
rect 53218 18286 53230 18338
rect 53282 18286 53294 18338
rect 43598 18274 43650 18286
rect 53566 18274 53618 18286
rect 54462 18338 54514 18350
rect 54462 18274 54514 18286
rect 55134 18338 55186 18350
rect 55134 18274 55186 18286
rect 52334 18226 52386 18238
rect 52334 18162 52386 18174
rect 53790 18226 53842 18238
rect 54574 18226 54626 18238
rect 54114 18174 54126 18226
rect 54178 18174 54190 18226
rect 53790 18162 53842 18174
rect 54574 18162 54626 18174
rect 55246 18226 55298 18238
rect 55246 18162 55298 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 51550 17890 51602 17902
rect 52782 17890 52834 17902
rect 51874 17838 51886 17890
rect 51938 17838 51950 17890
rect 51550 17826 51602 17838
rect 52782 17826 52834 17838
rect 22318 17778 22370 17790
rect 22318 17714 22370 17726
rect 35534 17778 35586 17790
rect 47070 17778 47122 17790
rect 38546 17726 38558 17778
rect 38610 17726 38622 17778
rect 40674 17726 40686 17778
rect 40738 17726 40750 17778
rect 42130 17726 42142 17778
rect 42194 17726 42206 17778
rect 44258 17726 44270 17778
rect 44322 17726 44334 17778
rect 35534 17714 35586 17726
rect 47070 17714 47122 17726
rect 50542 17778 50594 17790
rect 54338 17726 54350 17778
rect 54402 17726 54414 17778
rect 56466 17726 56478 17778
rect 56530 17726 56542 17778
rect 50542 17714 50594 17726
rect 17390 17666 17442 17678
rect 17390 17602 17442 17614
rect 17950 17666 18002 17678
rect 17950 17602 18002 17614
rect 18398 17666 18450 17678
rect 18398 17602 18450 17614
rect 18958 17666 19010 17678
rect 18958 17602 19010 17614
rect 19182 17666 19234 17678
rect 19182 17602 19234 17614
rect 19854 17666 19906 17678
rect 19854 17602 19906 17614
rect 21198 17666 21250 17678
rect 21198 17602 21250 17614
rect 21534 17666 21586 17678
rect 21534 17602 21586 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 23102 17666 23154 17678
rect 23102 17602 23154 17614
rect 30494 17666 30546 17678
rect 30494 17602 30546 17614
rect 30830 17666 30882 17678
rect 30830 17602 30882 17614
rect 31502 17666 31554 17678
rect 31502 17602 31554 17614
rect 32174 17666 32226 17678
rect 44942 17666 44994 17678
rect 35074 17614 35086 17666
rect 35138 17614 35150 17666
rect 37874 17614 37886 17666
rect 37938 17614 37950 17666
rect 41458 17614 41470 17666
rect 41522 17614 41534 17666
rect 32174 17602 32226 17614
rect 44942 17602 44994 17614
rect 46958 17666 47010 17678
rect 46958 17602 47010 17614
rect 47182 17666 47234 17678
rect 47182 17602 47234 17614
rect 50430 17666 50482 17678
rect 50430 17602 50482 17614
rect 50654 17666 50706 17678
rect 50654 17602 50706 17614
rect 50990 17666 51042 17678
rect 50990 17602 51042 17614
rect 51326 17666 51378 17678
rect 51326 17602 51378 17614
rect 52670 17666 52722 17678
rect 52670 17602 52722 17614
rect 53566 17666 53618 17678
rect 57250 17614 57262 17666
rect 57314 17614 57326 17666
rect 53566 17602 53618 17614
rect 17726 17554 17778 17566
rect 31166 17554 31218 17566
rect 58158 17554 58210 17566
rect 22754 17502 22766 17554
rect 22818 17502 22830 17554
rect 53330 17502 53342 17554
rect 53394 17502 53406 17554
rect 57810 17502 57822 17554
rect 57874 17502 57886 17554
rect 17726 17490 17778 17502
rect 31166 17490 31218 17502
rect 58158 17490 58210 17502
rect 17502 17442 17554 17454
rect 17502 17378 17554 17390
rect 18286 17442 18338 17454
rect 18286 17378 18338 17390
rect 18510 17442 18562 17454
rect 18510 17378 18562 17390
rect 19294 17442 19346 17454
rect 19294 17378 19346 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 28366 17442 28418 17454
rect 28366 17378 28418 17390
rect 30718 17442 30770 17454
rect 30718 17378 30770 17390
rect 31614 17442 31666 17454
rect 31614 17378 31666 17390
rect 31726 17442 31778 17454
rect 31726 17378 31778 17390
rect 35982 17442 36034 17454
rect 35982 17378 36034 17390
rect 46622 17442 46674 17454
rect 46622 17378 46674 17390
rect 47406 17442 47458 17454
rect 47406 17378 47458 17390
rect 53118 17442 53170 17454
rect 53118 17378 53170 17390
rect 53454 17442 53506 17454
rect 53454 17378 53506 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 18286 17106 18338 17118
rect 18286 17042 18338 17054
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 33182 17106 33234 17118
rect 33182 17042 33234 17054
rect 51886 17106 51938 17118
rect 51886 17042 51938 17054
rect 52110 17106 52162 17118
rect 52110 17042 52162 17054
rect 57486 17106 57538 17118
rect 57486 17042 57538 17054
rect 58270 17106 58322 17118
rect 58270 17042 58322 17054
rect 19070 16994 19122 17006
rect 27582 16994 27634 17006
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 20626 16942 20638 16994
rect 20690 16942 20702 16994
rect 19070 16930 19122 16942
rect 27582 16930 27634 16942
rect 28142 16994 28194 17006
rect 28142 16930 28194 16942
rect 28702 16994 28754 17006
rect 48974 16994 49026 17006
rect 30370 16942 30382 16994
rect 30434 16942 30446 16994
rect 28702 16930 28754 16942
rect 48974 16930 49026 16942
rect 17614 16882 17666 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 17614 16818 17666 16830
rect 18398 16882 18450 16894
rect 18398 16818 18450 16830
rect 18734 16882 18786 16894
rect 18734 16818 18786 16830
rect 19630 16882 19682 16894
rect 27694 16882 27746 16894
rect 19842 16830 19854 16882
rect 19906 16830 19918 16882
rect 19630 16818 19682 16830
rect 27694 16818 27746 16830
rect 28254 16882 28306 16894
rect 28254 16818 28306 16830
rect 28926 16882 28978 16894
rect 28926 16818 28978 16830
rect 29374 16882 29426 16894
rect 49310 16882 49362 16894
rect 29698 16830 29710 16882
rect 29762 16830 29774 16882
rect 29374 16818 29426 16830
rect 49310 16818 49362 16830
rect 51438 16882 51490 16894
rect 51438 16818 51490 16830
rect 52670 16882 52722 16894
rect 52670 16818 52722 16830
rect 52894 16882 52946 16894
rect 52894 16818 52946 16830
rect 53566 16882 53618 16894
rect 53566 16818 53618 16830
rect 27918 16770 27970 16782
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 22754 16718 22766 16770
rect 22818 16718 22830 16770
rect 27918 16706 27970 16718
rect 28814 16770 28866 16782
rect 41022 16770 41074 16782
rect 32498 16718 32510 16770
rect 32562 16718 32574 16770
rect 28814 16706 28866 16718
rect 41022 16706 41074 16718
rect 41470 16770 41522 16782
rect 41470 16706 41522 16718
rect 51214 16770 51266 16782
rect 51214 16706 51266 16718
rect 51998 16770 52050 16782
rect 51998 16706 52050 16718
rect 53342 16770 53394 16782
rect 53342 16706 53394 16718
rect 53790 16770 53842 16782
rect 53790 16706 53842 16718
rect 54014 16770 54066 16782
rect 54014 16706 54066 16718
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 19742 16210 19794 16222
rect 16706 16158 16718 16210
rect 16770 16158 16782 16210
rect 18834 16158 18846 16210
rect 18898 16158 18910 16210
rect 19742 16146 19794 16158
rect 22430 16210 22482 16222
rect 22430 16146 22482 16158
rect 25230 16210 25282 16222
rect 36094 16210 36146 16222
rect 35634 16158 35646 16210
rect 35698 16158 35710 16210
rect 25230 16146 25282 16158
rect 36094 16146 36146 16158
rect 38222 16210 38274 16222
rect 38222 16146 38274 16158
rect 41470 16210 41522 16222
rect 49298 16158 49310 16210
rect 49362 16158 49374 16210
rect 55234 16158 55246 16210
rect 55298 16158 55310 16210
rect 57362 16158 57374 16210
rect 57426 16158 57438 16210
rect 41470 16146 41522 16158
rect 22766 16098 22818 16110
rect 15922 16046 15934 16098
rect 15986 16046 15998 16098
rect 22766 16034 22818 16046
rect 22990 16098 23042 16110
rect 22990 16034 23042 16046
rect 27694 16098 27746 16110
rect 27694 16034 27746 16046
rect 29262 16098 29314 16110
rect 32398 16098 32450 16110
rect 32050 16046 32062 16098
rect 32114 16046 32126 16098
rect 29262 16034 29314 16046
rect 32398 16034 32450 16046
rect 32622 16098 32674 16110
rect 32622 16034 32674 16046
rect 33630 16098 33682 16110
rect 33630 16034 33682 16046
rect 33966 16098 34018 16110
rect 33966 16034 34018 16046
rect 49534 16098 49586 16110
rect 51650 16046 51662 16098
rect 51714 16046 51726 16098
rect 58034 16046 58046 16098
rect 58098 16046 58110 16098
rect 49534 16034 49586 16046
rect 19294 15986 19346 15998
rect 19294 15922 19346 15934
rect 23326 15986 23378 15998
rect 23326 15922 23378 15934
rect 24446 15986 24498 15998
rect 24446 15922 24498 15934
rect 24670 15986 24722 15998
rect 24670 15922 24722 15934
rect 27470 15986 27522 15998
rect 27470 15922 27522 15934
rect 28142 15986 28194 15998
rect 28142 15922 28194 15934
rect 28366 15986 28418 15998
rect 28366 15922 28418 15934
rect 29374 15986 29426 15998
rect 29374 15922 29426 15934
rect 29710 15986 29762 15998
rect 29710 15922 29762 15934
rect 34302 15986 34354 15998
rect 34302 15922 34354 15934
rect 35310 15986 35362 15998
rect 35310 15922 35362 15934
rect 35534 15986 35586 15998
rect 50542 15986 50594 15998
rect 47842 15934 47854 15986
rect 47906 15934 47918 15986
rect 35534 15922 35586 15934
rect 50542 15922 50594 15934
rect 22990 15874 23042 15886
rect 22990 15810 23042 15822
rect 24558 15874 24610 15886
rect 24558 15810 24610 15822
rect 27918 15874 27970 15886
rect 27918 15810 27970 15822
rect 29486 15874 29538 15886
rect 29486 15810 29538 15822
rect 33070 15874 33122 15886
rect 33070 15810 33122 15822
rect 33966 15874 34018 15886
rect 33966 15810 34018 15822
rect 37886 15874 37938 15886
rect 45726 15874 45778 15886
rect 45378 15822 45390 15874
rect 45442 15822 45454 15874
rect 37886 15810 37938 15822
rect 45726 15810 45778 15822
rect 52110 15874 52162 15886
rect 52110 15810 52162 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 29934 15538 29986 15550
rect 21858 15486 21870 15538
rect 21922 15486 21934 15538
rect 29934 15474 29986 15486
rect 33518 15538 33570 15550
rect 47742 15538 47794 15550
rect 38098 15486 38110 15538
rect 38162 15486 38174 15538
rect 33518 15474 33570 15486
rect 47742 15474 47794 15486
rect 52446 15538 52498 15550
rect 52446 15474 52498 15486
rect 58158 15538 58210 15550
rect 58158 15474 58210 15486
rect 24222 15426 24274 15438
rect 45054 15426 45106 15438
rect 27346 15374 27358 15426
rect 27410 15374 27422 15426
rect 35634 15374 35646 15426
rect 35698 15374 35710 15426
rect 39106 15374 39118 15426
rect 39170 15374 39182 15426
rect 24222 15362 24274 15374
rect 45054 15362 45106 15374
rect 49086 15426 49138 15438
rect 49086 15362 49138 15374
rect 49422 15426 49474 15438
rect 49422 15362 49474 15374
rect 50094 15426 50146 15438
rect 50094 15362 50146 15374
rect 50430 15426 50482 15438
rect 50430 15362 50482 15374
rect 31502 15314 31554 15326
rect 38446 15314 38498 15326
rect 40910 15314 40962 15326
rect 23762 15262 23774 15314
rect 23826 15262 23838 15314
rect 26674 15262 26686 15314
rect 26738 15262 26750 15314
rect 34962 15262 34974 15314
rect 35026 15262 35038 15314
rect 39554 15262 39566 15314
rect 39618 15262 39630 15314
rect 39890 15262 39902 15314
rect 39954 15262 39966 15314
rect 31502 15250 31554 15262
rect 38446 15250 38498 15262
rect 40910 15250 40962 15262
rect 41134 15314 41186 15326
rect 45278 15314 45330 15326
rect 41906 15262 41918 15314
rect 41970 15262 41982 15314
rect 41134 15250 41186 15262
rect 45278 15250 45330 15262
rect 45614 15314 45666 15326
rect 45614 15250 45666 15262
rect 46846 15314 46898 15326
rect 46846 15250 46898 15262
rect 47294 15314 47346 15326
rect 47294 15250 47346 15262
rect 48974 15314 49026 15326
rect 48974 15250 49026 15262
rect 50654 15314 50706 15326
rect 50654 15250 50706 15262
rect 51774 15314 51826 15326
rect 51774 15250 51826 15262
rect 51998 15314 52050 15326
rect 51998 15250 52050 15262
rect 52670 15314 52722 15326
rect 52670 15250 52722 15262
rect 22430 15202 22482 15214
rect 31726 15202 31778 15214
rect 38670 15202 38722 15214
rect 45166 15202 45218 15214
rect 23650 15150 23662 15202
rect 23714 15150 23726 15202
rect 29474 15150 29486 15202
rect 29538 15150 29550 15202
rect 37762 15150 37774 15202
rect 37826 15150 37838 15202
rect 39666 15150 39678 15202
rect 39730 15150 39742 15202
rect 42578 15150 42590 15202
rect 42642 15150 42654 15202
rect 44706 15150 44718 15202
rect 44770 15150 44782 15202
rect 22430 15138 22482 15150
rect 31726 15138 31778 15150
rect 38670 15138 38722 15150
rect 45166 15138 45218 15150
rect 46622 15202 46674 15214
rect 46622 15138 46674 15150
rect 47070 15202 47122 15214
rect 47070 15138 47122 15150
rect 49310 15202 49362 15214
rect 49310 15138 49362 15150
rect 50206 15202 50258 15214
rect 50206 15138 50258 15150
rect 51550 15202 51602 15214
rect 51550 15138 51602 15150
rect 52558 15202 52610 15214
rect 52558 15138 52610 15150
rect 22206 15090 22258 15102
rect 32050 15038 32062 15090
rect 32114 15038 32126 15090
rect 41458 15038 41470 15090
rect 41522 15038 41534 15090
rect 51202 15038 51214 15090
rect 51266 15038 51278 15090
rect 22206 15026 22258 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 50542 14754 50594 14766
rect 50542 14690 50594 14702
rect 52670 14754 52722 14766
rect 52670 14690 52722 14702
rect 52782 14754 52834 14766
rect 52782 14690 52834 14702
rect 18286 14642 18338 14654
rect 27582 14642 27634 14654
rect 50766 14642 50818 14654
rect 54014 14642 54066 14654
rect 24322 14590 24334 14642
rect 24386 14590 24398 14642
rect 26450 14590 26462 14642
rect 26514 14590 26526 14642
rect 34626 14590 34638 14642
rect 34690 14590 34702 14642
rect 38322 14590 38334 14642
rect 38386 14590 38398 14642
rect 41458 14590 41470 14642
rect 41522 14590 41534 14642
rect 53666 14590 53678 14642
rect 53730 14590 53742 14642
rect 54450 14590 54462 14642
rect 54514 14590 54526 14642
rect 18286 14578 18338 14590
rect 27582 14578 27634 14590
rect 50766 14578 50818 14590
rect 54014 14578 54066 14590
rect 18510 14530 18562 14542
rect 35422 14530 35474 14542
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 34962 14478 34974 14530
rect 35026 14478 35038 14530
rect 18510 14466 18562 14478
rect 35422 14466 35474 14478
rect 37550 14530 37602 14542
rect 42590 14530 42642 14542
rect 39778 14478 39790 14530
rect 39842 14478 39854 14530
rect 41682 14478 41694 14530
rect 41746 14478 41758 14530
rect 41906 14478 41918 14530
rect 41970 14478 41982 14530
rect 37550 14466 37602 14478
rect 42590 14466 42642 14478
rect 42814 14530 42866 14542
rect 42814 14466 42866 14478
rect 44718 14530 44770 14542
rect 44718 14466 44770 14478
rect 45054 14530 45106 14542
rect 45054 14466 45106 14478
rect 46846 14530 46898 14542
rect 46846 14466 46898 14478
rect 47182 14530 47234 14542
rect 47182 14466 47234 14478
rect 47854 14530 47906 14542
rect 47854 14466 47906 14478
rect 48078 14530 48130 14542
rect 51102 14530 51154 14542
rect 50194 14478 50206 14530
rect 50258 14478 50270 14530
rect 48078 14466 48130 14478
rect 51102 14466 51154 14478
rect 51214 14530 51266 14542
rect 53566 14530 53618 14542
rect 52098 14478 52110 14530
rect 52162 14478 52174 14530
rect 57250 14478 57262 14530
rect 57314 14478 57326 14530
rect 51214 14466 51266 14478
rect 53566 14466 53618 14478
rect 22654 14418 22706 14430
rect 22654 14354 22706 14366
rect 26798 14418 26850 14430
rect 40910 14418 40962 14430
rect 38994 14366 39006 14418
rect 39058 14366 39070 14418
rect 39554 14366 39566 14418
rect 39618 14366 39630 14418
rect 26798 14354 26850 14366
rect 40910 14354 40962 14366
rect 43038 14418 43090 14430
rect 43038 14354 43090 14366
rect 46622 14418 46674 14430
rect 54126 14418 54178 14430
rect 57822 14418 57874 14430
rect 51762 14366 51774 14418
rect 51826 14366 51838 14418
rect 53330 14366 53342 14418
rect 53394 14366 53406 14418
rect 56578 14366 56590 14418
rect 56642 14366 56654 14418
rect 46622 14354 46674 14366
rect 54126 14354 54178 14366
rect 57822 14354 57874 14366
rect 22094 14306 22146 14318
rect 18834 14254 18846 14306
rect 18898 14254 18910 14306
rect 22094 14242 22146 14254
rect 23214 14306 23266 14318
rect 33742 14306 33794 14318
rect 37886 14306 37938 14318
rect 42702 14306 42754 14318
rect 27122 14254 27134 14306
rect 27186 14254 27198 14306
rect 37202 14254 37214 14306
rect 37266 14254 37278 14306
rect 39218 14254 39230 14306
rect 39282 14254 39294 14306
rect 23214 14242 23266 14254
rect 33742 14242 33794 14254
rect 37886 14242 37938 14254
rect 42702 14242 42754 14254
rect 43710 14306 43762 14318
rect 43710 14242 43762 14254
rect 44942 14306 44994 14318
rect 44942 14242 44994 14254
rect 47070 14306 47122 14318
rect 51550 14306 51602 14318
rect 47506 14254 47518 14306
rect 47570 14254 47582 14306
rect 47070 14242 47122 14254
rect 51550 14242 51602 14254
rect 51886 14306 51938 14318
rect 51886 14242 51938 14254
rect 53118 14306 53170 14318
rect 53118 14242 53170 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 17502 13970 17554 13982
rect 17502 13906 17554 13918
rect 20750 13970 20802 13982
rect 20750 13906 20802 13918
rect 23886 13970 23938 13982
rect 23886 13906 23938 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 40014 13970 40066 13982
rect 40014 13906 40066 13918
rect 42478 13970 42530 13982
rect 42478 13906 42530 13918
rect 43262 13970 43314 13982
rect 43262 13906 43314 13918
rect 47630 13970 47682 13982
rect 47630 13906 47682 13918
rect 47854 13970 47906 13982
rect 47854 13906 47906 13918
rect 50654 13970 50706 13982
rect 50654 13906 50706 13918
rect 50766 13970 50818 13982
rect 50766 13906 50818 13918
rect 34302 13858 34354 13870
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 27906 13806 27918 13858
rect 27970 13806 27982 13858
rect 34302 13794 34354 13806
rect 34526 13858 34578 13870
rect 34526 13794 34578 13806
rect 35310 13858 35362 13870
rect 35310 13794 35362 13806
rect 41470 13858 41522 13870
rect 41470 13794 41522 13806
rect 42814 13858 42866 13870
rect 42814 13794 42866 13806
rect 44046 13858 44098 13870
rect 44046 13794 44098 13806
rect 44158 13858 44210 13870
rect 44158 13794 44210 13806
rect 44942 13858 44994 13870
rect 44942 13794 44994 13806
rect 45166 13858 45218 13870
rect 45166 13794 45218 13806
rect 52782 13858 52834 13870
rect 55234 13806 55246 13858
rect 55298 13806 55310 13858
rect 52782 13794 52834 13806
rect 18286 13746 18338 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 18286 13682 18338 13694
rect 18734 13746 18786 13758
rect 18734 13682 18786 13694
rect 18846 13746 18898 13758
rect 18846 13682 18898 13694
rect 18958 13746 19010 13758
rect 20862 13746 20914 13758
rect 19394 13694 19406 13746
rect 19458 13694 19470 13746
rect 19618 13694 19630 13746
rect 19682 13694 19694 13746
rect 19842 13694 19854 13746
rect 19906 13694 19918 13746
rect 18958 13682 19010 13694
rect 20862 13682 20914 13694
rect 21086 13746 21138 13758
rect 21086 13682 21138 13694
rect 21310 13746 21362 13758
rect 21310 13682 21362 13694
rect 21422 13746 21474 13758
rect 22430 13746 22482 13758
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 21422 13682 21474 13694
rect 22430 13682 22482 13694
rect 22654 13746 22706 13758
rect 22654 13682 22706 13694
rect 22766 13746 22818 13758
rect 22766 13682 22818 13694
rect 22990 13746 23042 13758
rect 22990 13682 23042 13694
rect 23326 13746 23378 13758
rect 33854 13746 33906 13758
rect 23650 13694 23662 13746
rect 23714 13694 23726 13746
rect 27122 13694 27134 13746
rect 27186 13694 27198 13746
rect 33058 13694 33070 13746
rect 33122 13694 33134 13746
rect 23326 13682 23378 13694
rect 33854 13682 33906 13694
rect 34750 13746 34802 13758
rect 39342 13746 39394 13758
rect 41918 13746 41970 13758
rect 35074 13694 35086 13746
rect 35138 13694 35150 13746
rect 39554 13694 39566 13746
rect 39618 13694 39630 13746
rect 41682 13694 41694 13746
rect 41746 13694 41758 13746
rect 34750 13682 34802 13694
rect 39342 13682 39394 13694
rect 41918 13682 41970 13694
rect 42366 13746 42418 13758
rect 42366 13682 42418 13694
rect 42702 13746 42754 13758
rect 42702 13682 42754 13694
rect 44382 13746 44434 13758
rect 50206 13746 50258 13758
rect 47282 13694 47294 13746
rect 47346 13694 47358 13746
rect 44382 13682 44434 13694
rect 50206 13682 50258 13694
rect 50878 13746 50930 13758
rect 50878 13682 50930 13694
rect 52670 13746 52722 13758
rect 55906 13694 55918 13746
rect 55970 13694 55982 13746
rect 52670 13682 52722 13694
rect 22206 13634 22258 13646
rect 30494 13634 30546 13646
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 23762 13582 23774 13634
rect 23826 13582 23838 13634
rect 30034 13582 30046 13634
rect 30098 13582 30110 13634
rect 22206 13570 22258 13582
rect 30494 13570 30546 13582
rect 32062 13634 32114 13646
rect 32062 13570 32114 13582
rect 32398 13634 32450 13646
rect 32398 13570 32450 13582
rect 34078 13634 34130 13646
rect 34078 13570 34130 13582
rect 34974 13634 35026 13646
rect 34974 13570 35026 13582
rect 35758 13634 35810 13646
rect 35758 13570 35810 13582
rect 37550 13634 37602 13646
rect 37550 13570 37602 13582
rect 38110 13634 38162 13646
rect 38110 13570 38162 13582
rect 38446 13634 38498 13646
rect 38446 13570 38498 13582
rect 42142 13634 42194 13646
rect 42142 13570 42194 13582
rect 43710 13634 43762 13646
rect 47742 13634 47794 13646
rect 56702 13634 56754 13646
rect 44930 13582 44942 13634
rect 44994 13582 45006 13634
rect 53106 13582 53118 13634
rect 53170 13582 53182 13634
rect 43710 13570 43762 13582
rect 47742 13570 47794 13582
rect 56702 13570 56754 13582
rect 32510 13522 32562 13534
rect 20402 13470 20414 13522
rect 20466 13470 20478 13522
rect 32510 13458 32562 13470
rect 33070 13522 33122 13534
rect 33070 13458 33122 13470
rect 33406 13522 33458 13534
rect 39006 13522 39058 13534
rect 37650 13470 37662 13522
rect 37714 13519 37726 13522
rect 38098 13519 38110 13522
rect 37714 13473 38110 13519
rect 37714 13470 37726 13473
rect 38098 13470 38110 13473
rect 38162 13470 38174 13522
rect 33406 13458 33458 13470
rect 39006 13458 39058 13470
rect 39118 13522 39170 13534
rect 39118 13458 39170 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 17838 13186 17890 13198
rect 17838 13122 17890 13134
rect 19966 13186 20018 13198
rect 19966 13122 20018 13134
rect 20526 13186 20578 13198
rect 20526 13122 20578 13134
rect 21310 13186 21362 13198
rect 21310 13122 21362 13134
rect 23550 13186 23602 13198
rect 23550 13122 23602 13134
rect 34526 13186 34578 13198
rect 34526 13122 34578 13134
rect 44830 13186 44882 13198
rect 44830 13122 44882 13134
rect 44942 13186 44994 13198
rect 44942 13122 44994 13134
rect 48190 13186 48242 13198
rect 48190 13122 48242 13134
rect 18734 13074 18786 13086
rect 18734 13010 18786 13022
rect 19182 13074 19234 13086
rect 19182 13010 19234 13022
rect 21422 13074 21474 13086
rect 34638 13074 34690 13086
rect 32386 13022 32398 13074
rect 32450 13022 32462 13074
rect 33058 13022 33070 13074
rect 33122 13022 33134 13074
rect 21422 13010 21474 13022
rect 34638 13010 34690 13022
rect 37102 13074 37154 13086
rect 48078 13074 48130 13086
rect 41010 13022 41022 13074
rect 41074 13022 41086 13074
rect 37102 13010 37154 13022
rect 48078 13010 48130 13022
rect 17950 12962 18002 12974
rect 17950 12898 18002 12910
rect 18398 12962 18450 12974
rect 18398 12898 18450 12910
rect 18622 12962 18674 12974
rect 18622 12898 18674 12910
rect 19854 12962 19906 12974
rect 23774 12962 23826 12974
rect 21634 12910 21646 12962
rect 21698 12910 21710 12962
rect 23314 12910 23326 12962
rect 23378 12910 23390 12962
rect 19854 12898 19906 12910
rect 23774 12898 23826 12910
rect 24110 12962 24162 12974
rect 24110 12898 24162 12910
rect 24446 12962 24498 12974
rect 34862 12962 34914 12974
rect 29474 12910 29486 12962
rect 29538 12910 29550 12962
rect 30258 12910 30270 12962
rect 30322 12910 30334 12962
rect 33282 12910 33294 12962
rect 33346 12910 33358 12962
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 24446 12898 24498 12910
rect 34862 12898 34914 12910
rect 35198 12962 35250 12974
rect 35198 12898 35250 12910
rect 35646 12962 35698 12974
rect 35646 12898 35698 12910
rect 35870 12962 35922 12974
rect 35870 12898 35922 12910
rect 36318 12962 36370 12974
rect 43710 12962 43762 12974
rect 39666 12910 39678 12962
rect 39730 12910 39742 12962
rect 36318 12898 36370 12910
rect 43710 12898 43762 12910
rect 45726 12962 45778 12974
rect 47170 12910 47182 12962
rect 47234 12910 47246 12962
rect 45726 12898 45778 12910
rect 18846 12850 18898 12862
rect 18846 12786 18898 12798
rect 20414 12850 20466 12862
rect 20414 12786 20466 12798
rect 22094 12850 22146 12862
rect 22094 12786 22146 12798
rect 22430 12850 22482 12862
rect 22430 12786 22482 12798
rect 22542 12850 22594 12862
rect 22542 12786 22594 12798
rect 22766 12850 22818 12862
rect 22766 12786 22818 12798
rect 22990 12850 23042 12862
rect 22990 12786 23042 12798
rect 24782 12850 24834 12862
rect 24782 12786 24834 12798
rect 34974 12850 35026 12862
rect 47854 12850 47906 12862
rect 42018 12798 42030 12850
rect 42082 12798 42094 12850
rect 45490 12798 45502 12850
rect 45554 12798 45566 12850
rect 47506 12798 47518 12850
rect 47570 12798 47582 12850
rect 34974 12786 35026 12798
rect 47854 12786 47906 12798
rect 17838 12738 17890 12750
rect 17838 12674 17890 12686
rect 19294 12738 19346 12750
rect 19294 12674 19346 12686
rect 19406 12738 19458 12750
rect 19406 12674 19458 12686
rect 19966 12738 20018 12750
rect 19966 12674 20018 12686
rect 23438 12738 23490 12750
rect 23438 12674 23490 12686
rect 24334 12738 24386 12750
rect 24334 12674 24386 12686
rect 25230 12738 25282 12750
rect 35534 12738 35586 12750
rect 33954 12686 33966 12738
rect 34018 12686 34030 12738
rect 25230 12674 25282 12686
rect 35534 12674 35586 12686
rect 38782 12738 38834 12750
rect 38782 12674 38834 12686
rect 42366 12738 42418 12750
rect 42366 12674 42418 12686
rect 42814 12738 42866 12750
rect 42814 12674 42866 12686
rect 43374 12738 43426 12750
rect 45278 12738 45330 12750
rect 44034 12686 44046 12738
rect 44098 12686 44110 12738
rect 43374 12674 43426 12686
rect 45278 12674 45330 12686
rect 45614 12738 45666 12750
rect 45614 12674 45666 12686
rect 47406 12738 47458 12750
rect 47406 12674 47458 12686
rect 51102 12738 51154 12750
rect 51102 12674 51154 12686
rect 51438 12738 51490 12750
rect 51438 12674 51490 12686
rect 53006 12738 53058 12750
rect 53006 12674 53058 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 20862 12402 20914 12414
rect 20862 12338 20914 12350
rect 23326 12402 23378 12414
rect 23326 12338 23378 12350
rect 24222 12402 24274 12414
rect 24222 12338 24274 12350
rect 24558 12402 24610 12414
rect 24558 12338 24610 12350
rect 28366 12402 28418 12414
rect 28366 12338 28418 12350
rect 33070 12402 33122 12414
rect 33070 12338 33122 12350
rect 34526 12402 34578 12414
rect 34526 12338 34578 12350
rect 39006 12402 39058 12414
rect 39006 12338 39058 12350
rect 39902 12402 39954 12414
rect 39902 12338 39954 12350
rect 41134 12402 41186 12414
rect 41134 12338 41186 12350
rect 42590 12402 42642 12414
rect 42590 12338 42642 12350
rect 50654 12402 50706 12414
rect 52110 12402 52162 12414
rect 51650 12350 51662 12402
rect 51714 12350 51726 12402
rect 50654 12338 50706 12350
rect 52110 12338 52162 12350
rect 27358 12290 27410 12302
rect 19506 12238 19518 12290
rect 19570 12238 19582 12290
rect 27358 12226 27410 12238
rect 34862 12290 34914 12302
rect 39118 12290 39170 12302
rect 35970 12238 35982 12290
rect 36034 12238 36046 12290
rect 34862 12226 34914 12238
rect 39118 12226 39170 12238
rect 40910 12290 40962 12302
rect 40910 12226 40962 12238
rect 44718 12290 44770 12302
rect 44718 12226 44770 12238
rect 47742 12290 47794 12302
rect 52222 12290 52274 12302
rect 50978 12238 50990 12290
rect 51042 12238 51054 12290
rect 47742 12226 47794 12238
rect 52222 12226 52274 12238
rect 52670 12290 52722 12302
rect 52670 12226 52722 12238
rect 27134 12178 27186 12190
rect 18274 12126 18286 12178
rect 18338 12126 18350 12178
rect 27134 12114 27186 12126
rect 27470 12178 27522 12190
rect 33294 12178 33346 12190
rect 30146 12126 30158 12178
rect 30210 12126 30222 12178
rect 27470 12114 27522 12126
rect 33294 12114 33346 12126
rect 33742 12178 33794 12190
rect 33742 12114 33794 12126
rect 34302 12178 34354 12190
rect 34302 12114 34354 12126
rect 34638 12178 34690 12190
rect 38782 12178 38834 12190
rect 35298 12126 35310 12178
rect 35362 12126 35374 12178
rect 34638 12114 34690 12126
rect 38782 12114 38834 12126
rect 39230 12178 39282 12190
rect 39230 12114 39282 12126
rect 39566 12178 39618 12190
rect 39566 12114 39618 12126
rect 39902 12178 39954 12190
rect 39902 12114 39954 12126
rect 40238 12178 40290 12190
rect 50318 12178 50370 12190
rect 49858 12126 49870 12178
rect 49922 12126 49934 12178
rect 40238 12114 40290 12126
rect 50318 12114 50370 12126
rect 51326 12178 51378 12190
rect 51326 12114 51378 12126
rect 51886 12178 51938 12190
rect 53330 12126 53342 12178
rect 53394 12126 53406 12178
rect 51886 12114 51938 12126
rect 21198 12066 21250 12078
rect 21198 12002 21250 12014
rect 27918 12066 27970 12078
rect 33182 12066 33234 12078
rect 41694 12066 41746 12078
rect 30818 12014 30830 12066
rect 30882 12014 30894 12066
rect 38098 12014 38110 12066
rect 38162 12014 38174 12066
rect 41234 12014 41246 12066
rect 41298 12014 41310 12066
rect 27918 12002 27970 12014
rect 33182 12002 33234 12014
rect 41694 12002 41746 12014
rect 42142 12066 42194 12078
rect 54450 12014 54462 12066
rect 54514 12014 54526 12066
rect 42142 12002 42194 12014
rect 44606 11954 44658 11966
rect 44146 11902 44158 11954
rect 44210 11951 44222 11954
rect 44370 11951 44382 11954
rect 44210 11905 44382 11951
rect 44210 11902 44222 11905
rect 44370 11902 44382 11905
rect 44434 11902 44446 11954
rect 44606 11890 44658 11902
rect 47854 11954 47906 11966
rect 47854 11890 47906 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 19630 11618 19682 11630
rect 19630 11554 19682 11566
rect 32062 11618 32114 11630
rect 57262 11618 57314 11630
rect 33058 11566 33070 11618
rect 33122 11615 33134 11618
rect 33394 11615 33406 11618
rect 33122 11569 33406 11615
rect 33122 11566 33134 11569
rect 33394 11566 33406 11569
rect 33458 11566 33470 11618
rect 32062 11554 32114 11566
rect 57262 11554 57314 11566
rect 17726 11506 17778 11518
rect 17266 11454 17278 11506
rect 17330 11454 17342 11506
rect 17726 11442 17778 11454
rect 19518 11506 19570 11518
rect 31838 11506 31890 11518
rect 24658 11454 24670 11506
rect 24722 11454 24734 11506
rect 19518 11442 19570 11454
rect 31838 11442 31890 11454
rect 33070 11506 33122 11518
rect 33070 11442 33122 11454
rect 33966 11506 34018 11518
rect 33966 11442 34018 11454
rect 35086 11506 35138 11518
rect 35086 11442 35138 11454
rect 38334 11506 38386 11518
rect 42366 11506 42418 11518
rect 40226 11454 40238 11506
rect 40290 11454 40302 11506
rect 38334 11442 38386 11454
rect 42366 11442 42418 11454
rect 43038 11506 43090 11518
rect 50094 11506 50146 11518
rect 46722 11454 46734 11506
rect 46786 11454 46798 11506
rect 48850 11454 48862 11506
rect 48914 11454 48926 11506
rect 43038 11442 43090 11454
rect 50094 11442 50146 11454
rect 50654 11506 50706 11518
rect 50654 11442 50706 11454
rect 51662 11506 51714 11518
rect 52658 11454 52670 11506
rect 52722 11454 52734 11506
rect 54786 11454 54798 11506
rect 54850 11454 54862 11506
rect 51662 11442 51714 11454
rect 18734 11394 18786 11406
rect 24334 11394 24386 11406
rect 28254 11394 28306 11406
rect 14466 11342 14478 11394
rect 14530 11342 14542 11394
rect 21522 11342 21534 11394
rect 21586 11342 21598 11394
rect 27570 11342 27582 11394
rect 27634 11342 27646 11394
rect 18734 11330 18786 11342
rect 24334 11330 24386 11342
rect 28254 11330 28306 11342
rect 29262 11394 29314 11406
rect 29262 11330 29314 11342
rect 31614 11394 31666 11406
rect 32622 11394 32674 11406
rect 50990 11394 51042 11406
rect 32274 11342 32286 11394
rect 32338 11342 32350 11394
rect 39442 11342 39454 11394
rect 39506 11342 39518 11394
rect 49634 11342 49646 11394
rect 49698 11342 49710 11394
rect 31614 11330 31666 11342
rect 32622 11330 32674 11342
rect 50990 11330 51042 11342
rect 51886 11394 51938 11406
rect 51886 11330 51938 11342
rect 52110 11394 52162 11406
rect 55570 11342 55582 11394
rect 55634 11342 55646 11394
rect 52110 11330 52162 11342
rect 19294 11282 19346 11294
rect 15138 11230 15150 11282
rect 15202 11230 15214 11282
rect 18946 11230 18958 11282
rect 19010 11230 19022 11282
rect 19294 11218 19346 11230
rect 21310 11282 21362 11294
rect 37886 11282 37938 11294
rect 26786 11230 26798 11282
rect 26850 11230 26862 11282
rect 21310 11218 21362 11230
rect 37886 11218 37938 11230
rect 38670 11282 38722 11294
rect 38670 11218 38722 11230
rect 51326 11282 51378 11294
rect 51326 11218 51378 11230
rect 51550 11282 51602 11294
rect 51550 11218 51602 11230
rect 57374 11282 57426 11294
rect 57374 11218 57426 11230
rect 57822 11282 57874 11294
rect 57822 11218 57874 11230
rect 58158 11282 58210 11294
rect 58158 11218 58210 11230
rect 18846 11170 18898 11182
rect 18846 11106 18898 11118
rect 20190 11170 20242 11182
rect 30718 11170 30770 11182
rect 23986 11118 23998 11170
rect 24050 11118 24062 11170
rect 27906 11118 27918 11170
rect 27970 11118 27982 11170
rect 20190 11106 20242 11118
rect 30718 11106 30770 11118
rect 31502 11170 31554 11182
rect 31502 11106 31554 11118
rect 33518 11170 33570 11182
rect 33518 11106 33570 11118
rect 39006 11170 39058 11182
rect 39006 11106 39058 11118
rect 51102 11170 51154 11182
rect 51102 11106 51154 11118
rect 56030 11170 56082 11182
rect 56030 11106 56082 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 15710 10834 15762 10846
rect 15710 10770 15762 10782
rect 18174 10834 18226 10846
rect 18174 10770 18226 10782
rect 25902 10834 25954 10846
rect 25902 10770 25954 10782
rect 26238 10834 26290 10846
rect 26238 10770 26290 10782
rect 26798 10834 26850 10846
rect 26798 10770 26850 10782
rect 42814 10834 42866 10846
rect 51998 10834 52050 10846
rect 50194 10782 50206 10834
rect 50258 10782 50270 10834
rect 42814 10770 42866 10782
rect 51998 10770 52050 10782
rect 15822 10722 15874 10734
rect 15822 10658 15874 10670
rect 18062 10722 18114 10734
rect 18062 10658 18114 10670
rect 18398 10722 18450 10734
rect 18398 10658 18450 10670
rect 18734 10722 18786 10734
rect 26350 10722 26402 10734
rect 23762 10670 23774 10722
rect 23826 10670 23838 10722
rect 18734 10658 18786 10670
rect 26350 10658 26402 10670
rect 27022 10722 27074 10734
rect 27022 10658 27074 10670
rect 31166 10722 31218 10734
rect 31166 10658 31218 10670
rect 31726 10722 31778 10734
rect 51326 10722 51378 10734
rect 43922 10670 43934 10722
rect 43986 10670 43998 10722
rect 47170 10670 47182 10722
rect 47234 10670 47246 10722
rect 31726 10658 31778 10670
rect 51326 10658 51378 10670
rect 51438 10722 51490 10734
rect 51438 10658 51490 10670
rect 52446 10722 52498 10734
rect 52446 10658 52498 10670
rect 17950 10610 18002 10622
rect 25342 10610 25394 10622
rect 24546 10558 24558 10610
rect 24610 10558 24622 10610
rect 17950 10546 18002 10558
rect 25342 10546 25394 10558
rect 26574 10610 26626 10622
rect 26574 10546 26626 10558
rect 27134 10610 27186 10622
rect 30942 10610 30994 10622
rect 30370 10558 30382 10610
rect 30434 10558 30446 10610
rect 27134 10546 27186 10558
rect 30942 10546 30994 10558
rect 31278 10610 31330 10622
rect 46846 10610 46898 10622
rect 41794 10558 41806 10610
rect 41858 10558 41870 10610
rect 43138 10558 43150 10610
rect 43202 10558 43214 10610
rect 31278 10546 31330 10558
rect 46846 10546 46898 10558
rect 49870 10610 49922 10622
rect 49870 10546 49922 10558
rect 51662 10610 51714 10622
rect 51662 10546 51714 10558
rect 58158 10610 58210 10622
rect 58158 10546 58210 10558
rect 42254 10498 42306 10510
rect 49534 10498 49586 10510
rect 21634 10446 21646 10498
rect 21698 10446 21710 10498
rect 27570 10446 27582 10498
rect 27634 10446 27646 10498
rect 29698 10446 29710 10498
rect 29762 10446 29774 10498
rect 46050 10446 46062 10498
rect 46114 10446 46126 10498
rect 42254 10434 42306 10446
rect 49534 10434 49586 10446
rect 50654 10498 50706 10510
rect 50654 10434 50706 10446
rect 18958 10386 19010 10398
rect 18958 10322 19010 10334
rect 19182 10386 19234 10398
rect 19182 10322 19234 10334
rect 19406 10386 19458 10398
rect 19406 10322 19458 10334
rect 19854 10386 19906 10398
rect 19854 10322 19906 10334
rect 26238 10386 26290 10398
rect 26238 10322 26290 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 18062 10050 18114 10062
rect 17714 9998 17726 10050
rect 17778 9998 17790 10050
rect 18062 9986 18114 9998
rect 19518 10050 19570 10062
rect 19518 9986 19570 9998
rect 32734 10050 32786 10062
rect 32734 9986 32786 9998
rect 20078 9938 20130 9950
rect 17266 9886 17278 9938
rect 17330 9886 17342 9938
rect 20078 9874 20130 9886
rect 22206 9938 22258 9950
rect 22206 9874 22258 9886
rect 30494 9938 30546 9950
rect 30494 9874 30546 9886
rect 32286 9938 32338 9950
rect 32286 9874 32338 9886
rect 35422 9938 35474 9950
rect 35422 9874 35474 9886
rect 42590 9938 42642 9950
rect 52658 9886 52670 9938
rect 52722 9886 52734 9938
rect 42590 9874 42642 9886
rect 18286 9826 18338 9838
rect 14466 9774 14478 9826
rect 14530 9774 14542 9826
rect 18286 9762 18338 9774
rect 18734 9826 18786 9838
rect 19630 9826 19682 9838
rect 18946 9774 18958 9826
rect 19010 9774 19022 9826
rect 18734 9762 18786 9774
rect 19630 9762 19682 9774
rect 21758 9826 21810 9838
rect 31838 9826 31890 9838
rect 24882 9774 24894 9826
rect 24946 9774 24958 9826
rect 25330 9774 25342 9826
rect 25394 9774 25406 9826
rect 27458 9774 27470 9826
rect 27522 9774 27534 9826
rect 28018 9774 28030 9826
rect 28082 9774 28094 9826
rect 31154 9774 31166 9826
rect 31218 9774 31230 9826
rect 21758 9762 21810 9774
rect 31838 9762 31890 9774
rect 33182 9826 33234 9838
rect 33182 9762 33234 9774
rect 33406 9826 33458 9838
rect 33406 9762 33458 9774
rect 33742 9826 33794 9838
rect 33742 9762 33794 9774
rect 35646 9826 35698 9838
rect 35646 9762 35698 9774
rect 35870 9826 35922 9838
rect 35870 9762 35922 9774
rect 36094 9826 36146 9838
rect 43486 9826 43538 9838
rect 37650 9774 37662 9826
rect 37714 9774 37726 9826
rect 41458 9774 41470 9826
rect 41522 9774 41534 9826
rect 43026 9774 43038 9826
rect 43090 9774 43102 9826
rect 36094 9762 36146 9774
rect 43486 9762 43538 9774
rect 43822 9826 43874 9838
rect 43822 9762 43874 9774
rect 50766 9826 50818 9838
rect 50766 9762 50818 9774
rect 51102 9826 51154 9838
rect 51102 9762 51154 9774
rect 51438 9826 51490 9838
rect 51438 9762 51490 9774
rect 51774 9826 51826 9838
rect 51774 9762 51826 9774
rect 51998 9826 52050 9838
rect 55570 9774 55582 9826
rect 55634 9774 55646 9826
rect 51998 9762 52050 9774
rect 19294 9714 19346 9726
rect 25902 9714 25954 9726
rect 29934 9714 29986 9726
rect 15138 9662 15150 9714
rect 15202 9662 15214 9714
rect 23426 9662 23438 9714
rect 23490 9662 23502 9714
rect 28578 9662 28590 9714
rect 28642 9662 28654 9714
rect 19294 9650 19346 9662
rect 25902 9650 25954 9662
rect 29934 9650 29986 9662
rect 30718 9714 30770 9726
rect 32734 9714 32786 9726
rect 31490 9662 31502 9714
rect 31554 9662 31566 9714
rect 30718 9650 30770 9662
rect 32734 9650 32786 9662
rect 32846 9714 32898 9726
rect 32846 9650 32898 9662
rect 34078 9714 34130 9726
rect 34078 9650 34130 9662
rect 34414 9714 34466 9726
rect 34414 9650 34466 9662
rect 36542 9714 36594 9726
rect 40350 9714 40402 9726
rect 50878 9714 50930 9726
rect 37762 9662 37774 9714
rect 37826 9662 37838 9714
rect 39554 9662 39566 9714
rect 39618 9662 39630 9714
rect 44146 9662 44158 9714
rect 44210 9662 44222 9714
rect 36542 9650 36594 9662
rect 40350 9650 40402 9662
rect 50878 9650 50930 9662
rect 51662 9714 51714 9726
rect 54786 9662 54798 9714
rect 54850 9662 54862 9714
rect 51662 9650 51714 9662
rect 18846 9602 18898 9614
rect 30046 9602 30098 9614
rect 21410 9550 21422 9602
rect 21474 9550 21486 9602
rect 27010 9550 27022 9602
rect 27074 9550 27086 9602
rect 27570 9550 27582 9602
rect 27634 9550 27646 9602
rect 18846 9538 18898 9550
rect 30046 9538 30098 9550
rect 30382 9602 30434 9614
rect 30382 9538 30434 9550
rect 30606 9602 30658 9614
rect 30606 9538 30658 9550
rect 33406 9602 33458 9614
rect 33406 9538 33458 9550
rect 50430 9602 50482 9614
rect 50430 9538 50482 9550
rect 56030 9602 56082 9614
rect 56030 9538 56082 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 15710 9266 15762 9278
rect 15710 9202 15762 9214
rect 17502 9266 17554 9278
rect 17502 9202 17554 9214
rect 18734 9266 18786 9278
rect 27582 9266 27634 9278
rect 22082 9214 22094 9266
rect 22146 9214 22158 9266
rect 18734 9202 18786 9214
rect 27582 9202 27634 9214
rect 31390 9266 31442 9278
rect 31390 9202 31442 9214
rect 33294 9266 33346 9278
rect 33294 9202 33346 9214
rect 33854 9266 33906 9278
rect 33854 9202 33906 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 41918 9266 41970 9278
rect 41918 9202 41970 9214
rect 44270 9266 44322 9278
rect 44270 9202 44322 9214
rect 50206 9266 50258 9278
rect 50206 9202 50258 9214
rect 51326 9266 51378 9278
rect 51326 9202 51378 9214
rect 15822 9154 15874 9166
rect 15822 9090 15874 9102
rect 18846 9154 18898 9166
rect 33518 9154 33570 9166
rect 31042 9102 31054 9154
rect 31106 9102 31118 9154
rect 18846 9090 18898 9102
rect 33518 9090 33570 9102
rect 33630 9154 33682 9166
rect 33630 9090 33682 9102
rect 35534 9154 35586 9166
rect 35534 9090 35586 9102
rect 37102 9154 37154 9166
rect 37102 9090 37154 9102
rect 37326 9154 37378 9166
rect 37326 9090 37378 9102
rect 37662 9154 37714 9166
rect 37662 9090 37714 9102
rect 39230 9154 39282 9166
rect 39230 9090 39282 9102
rect 39566 9154 39618 9166
rect 42814 9154 42866 9166
rect 43486 9154 43538 9166
rect 49982 9154 50034 9166
rect 39890 9102 39902 9154
rect 39954 9102 39966 9154
rect 42130 9102 42142 9154
rect 42194 9102 42206 9154
rect 43138 9102 43150 9154
rect 43202 9102 43214 9154
rect 43810 9102 43822 9154
rect 43874 9102 43886 9154
rect 39566 9090 39618 9102
rect 42814 9090 42866 9102
rect 43486 9090 43538 9102
rect 49982 9090 50034 9102
rect 18958 9042 19010 9054
rect 22430 9042 22482 9054
rect 19282 8990 19294 9042
rect 19346 8990 19358 9042
rect 18958 8978 19010 8990
rect 22430 8978 22482 8990
rect 35086 9042 35138 9054
rect 35086 8978 35138 8990
rect 35310 9042 35362 9054
rect 50430 9042 50482 9054
rect 42354 8990 42366 9042
rect 42418 8990 42430 9042
rect 44594 8990 44606 9042
rect 44658 8990 44670 9042
rect 35310 8978 35362 8990
rect 50430 8978 50482 8990
rect 35422 8930 35474 8942
rect 35422 8866 35474 8878
rect 37550 8930 37602 8942
rect 50318 8930 50370 8942
rect 45378 8878 45390 8930
rect 45442 8878 45454 8930
rect 47506 8878 47518 8930
rect 47570 8878 47582 8930
rect 37550 8866 37602 8878
rect 50318 8866 50370 8878
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 35310 8482 35362 8494
rect 35310 8418 35362 8430
rect 32510 8370 32562 8382
rect 32510 8306 32562 8318
rect 33630 8370 33682 8382
rect 33630 8306 33682 8318
rect 44942 8370 44994 8382
rect 44942 8306 44994 8318
rect 45390 8370 45442 8382
rect 45390 8306 45442 8318
rect 47406 8370 47458 8382
rect 47406 8306 47458 8318
rect 51214 8370 51266 8382
rect 51214 8306 51266 8318
rect 26910 8258 26962 8270
rect 26910 8194 26962 8206
rect 27358 8258 27410 8270
rect 27358 8194 27410 8206
rect 30942 8258 30994 8270
rect 30942 8194 30994 8206
rect 31502 8258 31554 8270
rect 31502 8194 31554 8206
rect 32174 8258 32226 8270
rect 35534 8258 35586 8270
rect 33954 8206 33966 8258
rect 34018 8206 34030 8258
rect 32174 8194 32226 8206
rect 35534 8194 35586 8206
rect 35870 8258 35922 8270
rect 35870 8194 35922 8206
rect 45166 8258 45218 8270
rect 45166 8194 45218 8206
rect 45614 8258 45666 8270
rect 45614 8194 45666 8206
rect 45838 8258 45890 8270
rect 45838 8194 45890 8206
rect 46286 8258 46338 8270
rect 46286 8194 46338 8206
rect 46398 8258 46450 8270
rect 46398 8194 46450 8206
rect 47182 8258 47234 8270
rect 47182 8194 47234 8206
rect 47518 8258 47570 8270
rect 47518 8194 47570 8206
rect 48414 8258 48466 8270
rect 48414 8194 48466 8206
rect 48638 8258 48690 8270
rect 48638 8194 48690 8206
rect 48862 8258 48914 8270
rect 50990 8258 51042 8270
rect 49522 8206 49534 8258
rect 49586 8206 49598 8258
rect 50418 8206 50430 8258
rect 50482 8206 50494 8258
rect 48862 8194 48914 8206
rect 50990 8194 51042 8206
rect 30606 8146 30658 8158
rect 30606 8082 30658 8094
rect 31166 8146 31218 8158
rect 31166 8082 31218 8094
rect 31614 8146 31666 8158
rect 31614 8082 31666 8094
rect 36318 8146 36370 8158
rect 36318 8082 36370 8094
rect 46622 8146 46674 8158
rect 46622 8082 46674 8094
rect 47854 8146 47906 8158
rect 47854 8082 47906 8094
rect 48190 8146 48242 8158
rect 49858 8094 49870 8146
rect 49922 8094 49934 8146
rect 48190 8082 48242 8094
rect 26686 8034 26738 8046
rect 26686 7970 26738 7982
rect 26798 8034 26850 8046
rect 26798 7970 26850 7982
rect 30718 8034 30770 8046
rect 30718 7970 30770 7982
rect 31726 8034 31778 8046
rect 31726 7970 31778 7982
rect 33742 8034 33794 8046
rect 35982 8034 36034 8046
rect 34962 7982 34974 8034
rect 35026 7982 35038 8034
rect 33742 7970 33794 7982
rect 35982 7970 36034 7982
rect 36094 8034 36146 8046
rect 36094 7970 36146 7982
rect 39006 8034 39058 8046
rect 39678 8034 39730 8046
rect 39330 7982 39342 8034
rect 39394 7982 39406 8034
rect 39006 7970 39058 7982
rect 39678 7970 39730 7982
rect 46174 8034 46226 8046
rect 46174 7970 46226 7982
rect 49310 8034 49362 8046
rect 50530 7982 50542 8034
rect 50594 7982 50606 8034
rect 51538 7982 51550 8034
rect 51602 7982 51614 8034
rect 49310 7970 49362 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 19070 7698 19122 7710
rect 19070 7634 19122 7646
rect 24782 7698 24834 7710
rect 24782 7634 24834 7646
rect 31502 7698 31554 7710
rect 31502 7634 31554 7646
rect 36766 7698 36818 7710
rect 36766 7634 36818 7646
rect 38446 7698 38498 7710
rect 38446 7634 38498 7646
rect 40014 7698 40066 7710
rect 40014 7634 40066 7646
rect 41358 7698 41410 7710
rect 41358 7634 41410 7646
rect 41470 7698 41522 7710
rect 41470 7634 41522 7646
rect 42590 7698 42642 7710
rect 42590 7634 42642 7646
rect 42926 7698 42978 7710
rect 42926 7634 42978 7646
rect 43598 7698 43650 7710
rect 43598 7634 43650 7646
rect 45838 7698 45890 7710
rect 45838 7634 45890 7646
rect 49646 7698 49698 7710
rect 49646 7634 49698 7646
rect 49758 7698 49810 7710
rect 49758 7634 49810 7646
rect 18958 7586 19010 7598
rect 18958 7522 19010 7534
rect 19630 7586 19682 7598
rect 19630 7522 19682 7534
rect 26798 7586 26850 7598
rect 33854 7586 33906 7598
rect 29810 7534 29822 7586
rect 29874 7534 29886 7586
rect 26798 7522 26850 7534
rect 33854 7522 33906 7534
rect 35646 7586 35698 7598
rect 39790 7586 39842 7598
rect 36418 7534 36430 7586
rect 36482 7534 36494 7586
rect 35646 7522 35698 7534
rect 39790 7522 39842 7534
rect 40126 7586 40178 7598
rect 43822 7586 43874 7598
rect 43250 7534 43262 7586
rect 43314 7534 43326 7586
rect 40126 7522 40178 7534
rect 43822 7522 43874 7534
rect 50878 7586 50930 7598
rect 51202 7534 51214 7586
rect 51266 7534 51278 7586
rect 50878 7522 50930 7534
rect 18846 7474 18898 7486
rect 18846 7410 18898 7422
rect 19406 7474 19458 7486
rect 19406 7410 19458 7422
rect 19854 7474 19906 7486
rect 19854 7410 19906 7422
rect 20302 7474 20354 7486
rect 20302 7410 20354 7422
rect 23326 7474 23378 7486
rect 23326 7410 23378 7422
rect 24110 7474 24162 7486
rect 24110 7410 24162 7422
rect 24334 7474 24386 7486
rect 24334 7410 24386 7422
rect 26350 7474 26402 7486
rect 26350 7410 26402 7422
rect 26574 7474 26626 7486
rect 26574 7410 26626 7422
rect 27022 7474 27074 7486
rect 27022 7410 27074 7422
rect 27246 7474 27298 7486
rect 33518 7474 33570 7486
rect 30482 7422 30494 7474
rect 30546 7422 30558 7474
rect 27246 7410 27298 7422
rect 33518 7410 33570 7422
rect 33630 7474 33682 7486
rect 34302 7474 34354 7486
rect 35310 7474 35362 7486
rect 36094 7474 36146 7486
rect 34178 7422 34190 7474
rect 34242 7422 34254 7474
rect 34514 7422 34526 7474
rect 34578 7422 34590 7474
rect 35074 7422 35086 7474
rect 35138 7422 35150 7474
rect 35410 7422 35422 7474
rect 35474 7422 35486 7474
rect 33630 7410 33682 7422
rect 34302 7410 34354 7422
rect 35310 7410 35362 7422
rect 36094 7410 36146 7422
rect 37886 7474 37938 7486
rect 37886 7410 37938 7422
rect 38110 7474 38162 7486
rect 38110 7410 38162 7422
rect 38670 7474 38722 7486
rect 38670 7410 38722 7422
rect 39118 7474 39170 7486
rect 39118 7410 39170 7422
rect 40350 7474 40402 7486
rect 40350 7410 40402 7422
rect 40798 7474 40850 7486
rect 40798 7410 40850 7422
rect 41246 7474 41298 7486
rect 44606 7474 44658 7486
rect 44146 7422 44158 7474
rect 44210 7422 44222 7474
rect 41246 7410 41298 7422
rect 44606 7410 44658 7422
rect 49870 7474 49922 7486
rect 50542 7474 50594 7486
rect 50194 7422 50206 7474
rect 50258 7422 50270 7474
rect 49870 7410 49922 7422
rect 50542 7410 50594 7422
rect 50654 7474 50706 7486
rect 50654 7410 50706 7422
rect 51438 7474 51490 7486
rect 51438 7410 51490 7422
rect 19742 7362 19794 7374
rect 19742 7298 19794 7310
rect 21310 7362 21362 7374
rect 21310 7298 21362 7310
rect 23662 7362 23714 7374
rect 31838 7362 31890 7374
rect 27682 7310 27694 7362
rect 27746 7310 27758 7362
rect 23662 7298 23714 7310
rect 31838 7298 31890 7310
rect 38558 7362 38610 7374
rect 38558 7298 38610 7310
rect 43710 7362 43762 7374
rect 52446 7362 52498 7374
rect 44146 7310 44158 7362
rect 44210 7359 44222 7362
rect 44482 7359 44494 7362
rect 44210 7313 44494 7359
rect 44210 7310 44222 7313
rect 44482 7310 44494 7313
rect 44546 7310 44558 7362
rect 51538 7310 51550 7362
rect 51602 7310 51614 7362
rect 43710 7298 43762 7310
rect 52446 7298 52498 7310
rect 21086 7250 21138 7262
rect 23102 7250 23154 7262
rect 20738 7198 20750 7250
rect 20802 7198 20814 7250
rect 22754 7198 22766 7250
rect 22818 7198 22830 7250
rect 21086 7186 21138 7198
rect 23102 7186 23154 7198
rect 23886 7250 23938 7262
rect 26126 7250 26178 7262
rect 25778 7198 25790 7250
rect 25842 7198 25854 7250
rect 23886 7186 23938 7198
rect 26126 7186 26178 7198
rect 35982 7250 36034 7262
rect 52558 7250 52610 7262
rect 37538 7198 37550 7250
rect 37602 7198 37614 7250
rect 35982 7186 36034 7198
rect 52558 7186 52610 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 19518 6914 19570 6926
rect 19518 6850 19570 6862
rect 19630 6914 19682 6926
rect 19630 6850 19682 6862
rect 21422 6914 21474 6926
rect 21422 6850 21474 6862
rect 23550 6914 23602 6926
rect 23550 6850 23602 6862
rect 26798 6914 26850 6926
rect 26798 6850 26850 6862
rect 26910 6914 26962 6926
rect 26910 6850 26962 6862
rect 38782 6914 38834 6926
rect 38782 6850 38834 6862
rect 38894 6914 38946 6926
rect 38894 6850 38946 6862
rect 40798 6914 40850 6926
rect 40798 6850 40850 6862
rect 40910 6914 40962 6926
rect 40910 6850 40962 6862
rect 41582 6914 41634 6926
rect 41582 6850 41634 6862
rect 50318 6914 50370 6926
rect 50318 6850 50370 6862
rect 20638 6802 20690 6814
rect 18274 6750 18286 6802
rect 18338 6750 18350 6802
rect 18610 6750 18622 6802
rect 18674 6750 18686 6802
rect 20638 6738 20690 6750
rect 21310 6802 21362 6814
rect 32286 6802 32338 6814
rect 22194 6750 22206 6802
rect 22258 6750 22270 6802
rect 24322 6750 24334 6802
rect 24386 6750 24398 6802
rect 25890 6750 25902 6802
rect 25954 6750 25966 6802
rect 21310 6738 21362 6750
rect 32286 6738 32338 6750
rect 36206 6802 36258 6814
rect 41806 6802 41858 6814
rect 41234 6750 41246 6802
rect 41298 6750 41310 6802
rect 36206 6738 36258 6750
rect 41806 6738 41858 6750
rect 48750 6802 48802 6814
rect 48750 6738 48802 6750
rect 49982 6802 50034 6814
rect 49982 6738 50034 6750
rect 50430 6802 50482 6814
rect 52658 6750 52670 6802
rect 52722 6750 52734 6802
rect 50430 6738 50482 6750
rect 18734 6690 18786 6702
rect 15474 6638 15486 6690
rect 15538 6638 15550 6690
rect 18734 6626 18786 6638
rect 20526 6690 20578 6702
rect 20526 6626 20578 6638
rect 23438 6690 23490 6702
rect 25118 6690 25170 6702
rect 24098 6638 24110 6690
rect 24162 6638 24174 6690
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 23438 6626 23490 6638
rect 25118 6626 25170 6638
rect 25454 6690 25506 6702
rect 27582 6690 27634 6702
rect 26226 6638 26238 6690
rect 26290 6638 26302 6690
rect 25454 6626 25506 6638
rect 27582 6626 27634 6638
rect 28030 6690 28082 6702
rect 28030 6626 28082 6638
rect 30158 6690 30210 6702
rect 30158 6626 30210 6638
rect 30270 6690 30322 6702
rect 30270 6626 30322 6638
rect 31278 6690 31330 6702
rect 31278 6626 31330 6638
rect 31950 6690 32002 6702
rect 42926 6690 42978 6702
rect 37874 6638 37886 6690
rect 37938 6638 37950 6690
rect 38210 6638 38222 6690
rect 38274 6638 38286 6690
rect 40226 6638 40238 6690
rect 40290 6638 40302 6690
rect 31950 6626 32002 6638
rect 42926 6626 42978 6638
rect 43486 6690 43538 6702
rect 43486 6626 43538 6638
rect 43934 6690 43986 6702
rect 43934 6626 43986 6638
rect 46398 6690 46450 6702
rect 46398 6626 46450 6638
rect 46846 6690 46898 6702
rect 46846 6626 46898 6638
rect 48414 6690 48466 6702
rect 48414 6626 48466 6638
rect 49758 6690 49810 6702
rect 56030 6690 56082 6702
rect 50978 6638 50990 6690
rect 51042 6638 51054 6690
rect 54786 6638 54798 6690
rect 54850 6638 54862 6690
rect 55458 6638 55470 6690
rect 55522 6638 55534 6690
rect 49758 6626 49810 6638
rect 56030 6626 56082 6638
rect 22206 6578 22258 6590
rect 16146 6526 16158 6578
rect 16210 6526 16222 6578
rect 18946 6526 18958 6578
rect 19010 6526 19022 6578
rect 21970 6526 21982 6578
rect 22034 6526 22046 6578
rect 22206 6514 22258 6526
rect 24782 6578 24834 6590
rect 24782 6514 24834 6526
rect 25230 6578 25282 6590
rect 25230 6514 25282 6526
rect 26014 6578 26066 6590
rect 26014 6514 26066 6526
rect 26574 6578 26626 6590
rect 30942 6578 30994 6590
rect 27234 6526 27246 6578
rect 27298 6526 27310 6578
rect 26574 6514 26626 6526
rect 30942 6514 30994 6526
rect 38558 6578 38610 6590
rect 38558 6514 38610 6526
rect 40014 6578 40066 6590
rect 40014 6514 40066 6526
rect 40574 6578 40626 6590
rect 40574 6514 40626 6526
rect 43262 6578 43314 6590
rect 43262 6514 43314 6526
rect 48526 6578 48578 6590
rect 48526 6514 48578 6526
rect 48862 6578 48914 6590
rect 50766 6578 50818 6590
rect 49410 6526 49422 6578
rect 49474 6526 49486 6578
rect 48862 6514 48914 6526
rect 50766 6514 50818 6526
rect 51214 6578 51266 6590
rect 51214 6514 51266 6526
rect 19182 6466 19234 6478
rect 19182 6402 19234 6414
rect 20302 6466 20354 6478
rect 20302 6402 20354 6414
rect 20750 6466 20802 6478
rect 20750 6402 20802 6414
rect 21758 6466 21810 6478
rect 21758 6402 21810 6414
rect 23886 6466 23938 6478
rect 23886 6402 23938 6414
rect 30718 6466 30770 6478
rect 30718 6402 30770 6414
rect 30830 6466 30882 6478
rect 30830 6402 30882 6414
rect 31390 6466 31442 6478
rect 31390 6402 31442 6414
rect 31502 6466 31554 6478
rect 31502 6402 31554 6414
rect 38110 6466 38162 6478
rect 38110 6402 38162 6414
rect 40126 6466 40178 6478
rect 40126 6402 40178 6414
rect 43150 6466 43202 6478
rect 43150 6402 43202 6414
rect 51102 6466 51154 6478
rect 51102 6402 51154 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 17390 6130 17442 6142
rect 17390 6066 17442 6078
rect 23662 6130 23714 6142
rect 23662 6066 23714 6078
rect 23774 6130 23826 6142
rect 23774 6066 23826 6078
rect 31166 6130 31218 6142
rect 31166 6066 31218 6078
rect 32062 6130 32114 6142
rect 32062 6066 32114 6078
rect 32398 6130 32450 6142
rect 32398 6066 32450 6078
rect 46286 6130 46338 6142
rect 46286 6066 46338 6078
rect 46734 6130 46786 6142
rect 46734 6066 46786 6078
rect 21534 6018 21586 6030
rect 21534 5954 21586 5966
rect 31278 6018 31330 6030
rect 31278 5954 31330 5966
rect 33854 6018 33906 6030
rect 33854 5954 33906 5966
rect 35422 6018 35474 6030
rect 45054 6018 45106 6030
rect 43698 5966 43710 6018
rect 43762 5966 43774 6018
rect 35422 5954 35474 5966
rect 45054 5954 45106 5966
rect 46174 6018 46226 6030
rect 46174 5954 46226 5966
rect 46510 6018 46562 6030
rect 46510 5954 46562 5966
rect 46958 6018 47010 6030
rect 46958 5954 47010 5966
rect 47070 6018 47122 6030
rect 47282 5966 47294 6018
rect 47346 5966 47358 6018
rect 47070 5954 47122 5966
rect 17502 5906 17554 5918
rect 17502 5842 17554 5854
rect 19070 5906 19122 5918
rect 19070 5842 19122 5854
rect 19294 5906 19346 5918
rect 19294 5842 19346 5854
rect 21758 5906 21810 5918
rect 21758 5842 21810 5854
rect 21982 5906 22034 5918
rect 21982 5842 22034 5854
rect 23550 5906 23602 5918
rect 30942 5906 30994 5918
rect 24098 5854 24110 5906
rect 24162 5854 24174 5906
rect 30482 5854 30494 5906
rect 30546 5854 30558 5906
rect 23550 5842 23602 5854
rect 30942 5842 30994 5854
rect 31390 5906 31442 5918
rect 45278 5906 45330 5918
rect 44370 5854 44382 5906
rect 44434 5854 44446 5906
rect 31390 5842 31442 5854
rect 45278 5842 45330 5854
rect 45614 5906 45666 5918
rect 45614 5842 45666 5854
rect 18398 5794 18450 5806
rect 18398 5730 18450 5742
rect 21646 5794 21698 5806
rect 41246 5794 41298 5806
rect 45166 5794 45218 5806
rect 27570 5742 27582 5794
rect 27634 5742 27646 5794
rect 29698 5742 29710 5794
rect 29762 5742 29774 5794
rect 41570 5742 41582 5794
rect 41634 5742 41646 5794
rect 47506 5742 47518 5794
rect 47570 5742 47582 5794
rect 21646 5730 21698 5742
rect 41246 5730 41298 5742
rect 45166 5730 45218 5742
rect 33742 5682 33794 5694
rect 18722 5630 18734 5682
rect 18786 5630 18798 5682
rect 33742 5618 33794 5630
rect 35534 5682 35586 5694
rect 35534 5618 35586 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 20190 5234 20242 5246
rect 20190 5170 20242 5182
rect 21422 5234 21474 5246
rect 21422 5170 21474 5182
rect 23214 5234 23266 5246
rect 23214 5170 23266 5182
rect 25902 5234 25954 5246
rect 25902 5170 25954 5182
rect 31614 5234 31666 5246
rect 31614 5170 31666 5182
rect 32062 5234 32114 5246
rect 40350 5234 40402 5246
rect 33506 5182 33518 5234
rect 33570 5182 33582 5234
rect 35634 5182 35646 5234
rect 35698 5182 35710 5234
rect 36978 5182 36990 5234
rect 37042 5182 37054 5234
rect 32062 5170 32114 5182
rect 40350 5170 40402 5182
rect 40686 5234 40738 5246
rect 40686 5170 40738 5182
rect 44046 5234 44098 5246
rect 44046 5170 44098 5182
rect 44942 5234 44994 5246
rect 44942 5170 44994 5182
rect 45502 5234 45554 5246
rect 51214 5234 51266 5246
rect 47730 5182 47742 5234
rect 47794 5182 47806 5234
rect 49858 5182 49870 5234
rect 49922 5182 49934 5234
rect 45502 5170 45554 5182
rect 51214 5170 51266 5182
rect 30718 5122 30770 5134
rect 30718 5058 30770 5070
rect 30830 5122 30882 5134
rect 30830 5058 30882 5070
rect 31054 5122 31106 5134
rect 31054 5058 31106 5070
rect 31166 5122 31218 5134
rect 45838 5122 45890 5134
rect 32722 5070 32734 5122
rect 32786 5070 32798 5122
rect 39106 5070 39118 5122
rect 39170 5070 39182 5122
rect 39890 5070 39902 5122
rect 39954 5070 39966 5122
rect 31166 5058 31218 5070
rect 45838 5058 45890 5070
rect 46510 5122 46562 5134
rect 50318 5122 50370 5134
rect 47058 5070 47070 5122
rect 47122 5070 47134 5122
rect 46510 5058 46562 5070
rect 50318 5058 50370 5070
rect 20078 4898 20130 4910
rect 20078 4834 20130 4846
rect 23102 4898 23154 4910
rect 23102 4834 23154 4846
rect 26014 4898 26066 4910
rect 26014 4834 26066 4846
rect 40798 4898 40850 4910
rect 40798 4834 40850 4846
rect 45950 4898 46002 4910
rect 45950 4834 46002 4846
rect 46062 4898 46114 4910
rect 46062 4834 46114 4846
rect 51326 4898 51378 4910
rect 51326 4834 51378 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 28590 4562 28642 4574
rect 28590 4498 28642 4510
rect 33182 4562 33234 4574
rect 33182 4498 33234 4510
rect 37662 4562 37714 4574
rect 37662 4498 37714 4510
rect 38222 4562 38274 4574
rect 38222 4498 38274 4510
rect 48750 4562 48802 4574
rect 48750 4498 48802 4510
rect 53902 4562 53954 4574
rect 53902 4498 53954 4510
rect 38110 4450 38162 4462
rect 48862 4450 48914 4462
rect 19058 4398 19070 4450
rect 19122 4398 19134 4450
rect 22306 4398 22318 4450
rect 22370 4398 22382 4450
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 31490 4398 31502 4450
rect 31554 4398 31566 4450
rect 36418 4398 36430 4450
rect 36482 4398 36494 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 44930 4398 44942 4450
rect 44994 4398 45006 4450
rect 52658 4398 52670 4450
rect 52722 4398 52734 4450
rect 38110 4386 38162 4398
rect 48862 4386 48914 4398
rect 57598 4338 57650 4350
rect 18386 4286 18398 4338
rect 18450 4286 18462 4338
rect 21522 4286 21534 4338
rect 21586 4286 21598 4338
rect 25330 4286 25342 4338
rect 25394 4286 25406 4338
rect 32274 4286 32286 4338
rect 32338 4286 32350 4338
rect 37202 4286 37214 4338
rect 37266 4286 37278 4338
rect 40898 4286 40910 4338
rect 40962 4286 40974 4338
rect 44146 4286 44158 4338
rect 44210 4286 44222 4338
rect 53330 4286 53342 4338
rect 53394 4286 53406 4338
rect 57598 4274 57650 4286
rect 58158 4338 58210 4350
rect 58158 4274 58210 4286
rect 57374 4226 57426 4238
rect 21186 4174 21198 4226
rect 21250 4174 21262 4226
rect 24434 4174 24446 4226
rect 24498 4174 24510 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 29362 4174 29374 4226
rect 29426 4174 29438 4226
rect 34290 4174 34302 4226
rect 34354 4174 34366 4226
rect 43810 4174 43822 4226
rect 43874 4174 43886 4226
rect 47058 4174 47070 4226
rect 47122 4174 47134 4226
rect 50530 4174 50542 4226
rect 50594 4174 50606 4226
rect 57374 4162 57426 4174
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 21534 3666 21586 3678
rect 21534 3602 21586 3614
rect 43934 3666 43986 3678
rect 43934 3602 43986 3614
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 8766 66782 8818 66834
rect 9326 66782 9378 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 26126 66446 26178 66498
rect 40798 66446 40850 66498
rect 43822 66446 43874 66498
rect 48414 66446 48466 66498
rect 52222 66446 52274 66498
rect 56030 66446 56082 66498
rect 18846 66334 18898 66386
rect 22878 66334 22930 66386
rect 36990 66334 37042 66386
rect 17614 66222 17666 66274
rect 23550 66222 23602 66274
rect 25118 66222 25170 66274
rect 39230 66222 39282 66274
rect 39790 66222 39842 66274
rect 46174 66222 46226 66274
rect 47406 66222 47458 66274
rect 51214 66222 51266 66274
rect 55022 66222 55074 66274
rect 2942 66110 2994 66162
rect 5518 66110 5570 66162
rect 6974 66110 7026 66162
rect 9326 66110 9378 66162
rect 11006 66110 11058 66162
rect 13134 66110 13186 66162
rect 15038 66110 15090 66162
rect 17054 66110 17106 66162
rect 29150 66110 29202 66162
rect 31166 66110 31218 66162
rect 33182 66110 33234 66162
rect 35198 66110 35250 66162
rect 43038 66110 43090 66162
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 34862 65550 34914 65602
rect 57822 65550 57874 65602
rect 20190 65438 20242 65490
rect 21870 65438 21922 65490
rect 29710 65438 29762 65490
rect 35534 65438 35586 65490
rect 36654 65438 36706 65490
rect 44382 65438 44434 65490
rect 44830 65438 44882 65490
rect 48862 65438 48914 65490
rect 54910 65438 54962 65490
rect 57598 65438 57650 65490
rect 58158 65438 58210 65490
rect 8878 65326 8930 65378
rect 12462 65326 12514 65378
rect 17390 65326 17442 65378
rect 19518 65326 19570 65378
rect 20862 65326 20914 65378
rect 22542 65326 22594 65378
rect 24670 65326 24722 65378
rect 25454 65326 25506 65378
rect 27358 65326 27410 65378
rect 30270 65326 30322 65378
rect 34974 65326 35026 65378
rect 37438 65326 37490 65378
rect 39566 65326 39618 65378
rect 40126 65326 40178 65378
rect 41134 65326 41186 65378
rect 41582 65326 41634 65378
rect 43710 65326 43762 65378
rect 45614 65326 45666 65378
rect 47742 65326 47794 65378
rect 49534 65326 49586 65378
rect 51662 65326 51714 65378
rect 51998 65326 52050 65378
rect 54126 65326 54178 65378
rect 55470 65326 55522 65378
rect 35086 65214 35138 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 23550 64878 23602 64930
rect 42702 64878 42754 64930
rect 47518 64878 47570 64930
rect 50206 64878 50258 64930
rect 51774 64878 51826 64930
rect 8542 64766 8594 64818
rect 12126 64766 12178 64818
rect 20750 64766 20802 64818
rect 26910 64766 26962 64818
rect 33518 64766 33570 64818
rect 35646 64766 35698 64818
rect 41358 64766 41410 64818
rect 44942 64766 44994 64818
rect 45390 64766 45442 64818
rect 55246 64766 55298 64818
rect 5742 64654 5794 64706
rect 9326 64654 9378 64706
rect 13470 64654 13522 64706
rect 17950 64654 18002 64706
rect 23998 64654 24050 64706
rect 27918 64654 27970 64706
rect 29038 64654 29090 64706
rect 29486 64654 29538 64706
rect 30382 64654 30434 64706
rect 36430 64654 36482 64706
rect 37102 64654 37154 64706
rect 38558 64654 38610 64706
rect 41694 64654 41746 64706
rect 49422 64654 49474 64706
rect 54574 64654 54626 64706
rect 58046 64654 58098 64706
rect 6414 64542 6466 64594
rect 9998 64542 10050 64594
rect 12686 64542 12738 64594
rect 13806 64542 13858 64594
rect 18622 64542 18674 64594
rect 23662 64542 23714 64594
rect 24782 64542 24834 64594
rect 30942 64542 30994 64594
rect 32510 64542 32562 64594
rect 32622 64542 32674 64594
rect 32958 64542 33010 64594
rect 39230 64542 39282 64594
rect 50318 64542 50370 64594
rect 51662 64542 51714 64594
rect 57374 64542 57426 64594
rect 12798 64430 12850 64482
rect 13022 64430 13074 64482
rect 13694 64430 13746 64482
rect 21422 64430 21474 64482
rect 23214 64430 23266 64482
rect 27246 64430 27298 64482
rect 27358 64430 27410 64482
rect 27470 64430 27522 64482
rect 28702 64430 28754 64482
rect 29598 64430 29650 64482
rect 29710 64430 29762 64482
rect 30830 64430 30882 64482
rect 31054 64430 31106 64482
rect 31502 64430 31554 64482
rect 32286 64430 32338 64482
rect 33070 64430 33122 64482
rect 33294 64430 33346 64482
rect 52782 64430 52834 64482
rect 54014 64430 54066 64482
rect 54350 64430 54402 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 12798 64094 12850 64146
rect 17614 64094 17666 64146
rect 27806 64094 27858 64146
rect 32286 64094 32338 64146
rect 41582 64094 41634 64146
rect 42030 64094 42082 64146
rect 46734 64094 46786 64146
rect 50430 64094 50482 64146
rect 52334 64094 52386 64146
rect 54574 64094 54626 64146
rect 8542 63982 8594 64034
rect 11454 63982 11506 64034
rect 17726 63982 17778 64034
rect 27470 63982 27522 64034
rect 27582 63982 27634 64034
rect 31950 63982 32002 64034
rect 35198 63982 35250 64034
rect 46846 63982 46898 64034
rect 50878 63982 50930 64034
rect 51214 63982 51266 64034
rect 56030 63982 56082 64034
rect 56814 63982 56866 64034
rect 11790 63870 11842 63922
rect 12462 63870 12514 63922
rect 13582 63870 13634 63922
rect 16830 63870 16882 63922
rect 17278 63870 17330 63922
rect 17838 63870 17890 63922
rect 20190 63870 20242 63922
rect 23438 63870 23490 63922
rect 26686 63870 26738 63922
rect 28030 63870 28082 63922
rect 32062 63870 32114 63922
rect 32510 63870 32562 63922
rect 33518 63870 33570 63922
rect 34638 63870 34690 63922
rect 39454 63870 39506 63922
rect 43374 63870 43426 63922
rect 43822 63870 43874 63922
rect 46398 63870 46450 63922
rect 47070 63870 47122 63922
rect 49534 63870 49586 63922
rect 49646 63870 49698 63922
rect 49982 63870 50034 63922
rect 50094 63870 50146 63922
rect 51326 63870 51378 63922
rect 54126 63870 54178 63922
rect 54798 63870 54850 63922
rect 14254 63758 14306 63810
rect 16382 63758 16434 63810
rect 20862 63758 20914 63810
rect 22990 63758 23042 63810
rect 26350 63758 26402 63810
rect 27134 63758 27186 63810
rect 28814 63758 28866 63810
rect 30942 63758 30994 63810
rect 31726 63758 31778 63810
rect 33182 63758 33234 63810
rect 50430 63758 50482 63810
rect 50766 63758 50818 63810
rect 54686 63758 54738 63810
rect 8430 63646 8482 63698
rect 43038 63646 43090 63698
rect 43374 63646 43426 63698
rect 56590 63646 56642 63698
rect 56926 63646 56978 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 12014 63310 12066 63362
rect 12350 63310 12402 63362
rect 12686 63310 12738 63362
rect 19630 63310 19682 63362
rect 22318 63310 22370 63362
rect 31278 63310 31330 63362
rect 53566 63310 53618 63362
rect 54462 63310 54514 63362
rect 6638 63198 6690 63250
rect 11902 63198 11954 63250
rect 17502 63198 17554 63250
rect 26238 63198 26290 63250
rect 32062 63198 32114 63250
rect 45166 63198 45218 63250
rect 47742 63198 47794 63250
rect 51438 63198 51490 63250
rect 51662 63198 51714 63250
rect 53006 63198 53058 63250
rect 53902 63198 53954 63250
rect 54910 63198 54962 63250
rect 55246 63198 55298 63250
rect 57374 63198 57426 63250
rect 6750 63086 6802 63138
rect 7870 63086 7922 63138
rect 8094 63086 8146 63138
rect 15486 63086 15538 63138
rect 16270 63086 16322 63138
rect 19630 63086 19682 63138
rect 21310 63086 21362 63138
rect 26686 63086 26738 63138
rect 27134 63086 27186 63138
rect 27582 63086 27634 63138
rect 27806 63086 27858 63138
rect 28142 63086 28194 63138
rect 30158 63086 30210 63138
rect 30382 63086 30434 63138
rect 32174 63086 32226 63138
rect 32398 63086 32450 63138
rect 41246 63086 41298 63138
rect 43486 63086 43538 63138
rect 44046 63086 44098 63138
rect 44942 63086 44994 63138
rect 46062 63086 46114 63138
rect 46510 63086 46562 63138
rect 50654 63086 50706 63138
rect 50766 63086 50818 63138
rect 51102 63086 51154 63138
rect 51214 63086 51266 63138
rect 51774 63086 51826 63138
rect 53230 63086 53282 63138
rect 54126 63086 54178 63138
rect 58046 63086 58098 63138
rect 6526 62974 6578 63026
rect 7086 62974 7138 63026
rect 7646 62974 7698 63026
rect 14814 62974 14866 63026
rect 16382 62974 16434 63026
rect 17614 62974 17666 63026
rect 19966 62974 20018 63026
rect 26126 62974 26178 63026
rect 26462 62974 26514 63026
rect 28030 62974 28082 63026
rect 29486 62974 29538 63026
rect 31166 62974 31218 63026
rect 31278 62974 31330 63026
rect 31950 62974 32002 63026
rect 41022 62974 41074 63026
rect 42254 62974 42306 63026
rect 44158 62974 44210 63026
rect 45054 62974 45106 63026
rect 45502 62974 45554 63026
rect 45838 62974 45890 63026
rect 12462 62862 12514 62914
rect 13694 62862 13746 62914
rect 17390 62862 17442 62914
rect 17838 62862 17890 62914
rect 18510 62862 18562 62914
rect 27022 62862 27074 62914
rect 27246 62862 27298 62914
rect 28590 62862 28642 62914
rect 32846 62862 32898 62914
rect 42478 62862 42530 62914
rect 42926 62862 42978 62914
rect 44382 62862 44434 62914
rect 45278 62862 45330 62914
rect 47182 62862 47234 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 7198 62526 7250 62578
rect 7310 62526 7362 62578
rect 7982 62526 8034 62578
rect 13918 62526 13970 62578
rect 14926 62526 14978 62578
rect 16494 62526 16546 62578
rect 16718 62526 16770 62578
rect 19406 62526 19458 62578
rect 19966 62526 20018 62578
rect 29038 62526 29090 62578
rect 44046 62526 44098 62578
rect 44718 62526 44770 62578
rect 45502 62526 45554 62578
rect 45614 62526 45666 62578
rect 47182 62526 47234 62578
rect 52110 62526 52162 62578
rect 6862 62414 6914 62466
rect 8542 62414 8594 62466
rect 10894 62414 10946 62466
rect 13134 62414 13186 62466
rect 14814 62414 14866 62466
rect 18958 62414 19010 62466
rect 28926 62414 28978 62466
rect 37886 62414 37938 62466
rect 39454 62414 39506 62466
rect 41918 62414 41970 62466
rect 43262 62414 43314 62466
rect 47294 62414 47346 62466
rect 52446 62414 52498 62466
rect 56926 62414 56978 62466
rect 57374 62414 57426 62466
rect 7086 62302 7138 62354
rect 7870 62302 7922 62354
rect 8206 62302 8258 62354
rect 8430 62302 8482 62354
rect 8766 62302 8818 62354
rect 9438 62302 9490 62354
rect 10222 62302 10274 62354
rect 12910 62302 12962 62354
rect 13806 62302 13858 62354
rect 15150 62302 15202 62354
rect 16382 62302 16434 62354
rect 19182 62302 19234 62354
rect 19518 62302 19570 62354
rect 19854 62302 19906 62354
rect 20078 62302 20130 62354
rect 20414 62302 20466 62354
rect 29150 62302 29202 62354
rect 29374 62302 29426 62354
rect 37214 62302 37266 62354
rect 38782 62302 38834 62354
rect 41246 62302 41298 62354
rect 42814 62302 42866 62354
rect 43486 62302 43538 62354
rect 43934 62302 43986 62354
rect 44158 62302 44210 62354
rect 44606 62302 44658 62354
rect 44942 62302 44994 62354
rect 45054 62302 45106 62354
rect 45726 62302 45778 62354
rect 45950 62302 46002 62354
rect 46286 62302 46338 62354
rect 46510 62302 46562 62354
rect 46958 62302 47010 62354
rect 48862 62302 48914 62354
rect 53454 62302 53506 62354
rect 56702 62302 56754 62354
rect 57150 62302 57202 62354
rect 57486 62302 57538 62354
rect 10558 62190 10610 62242
rect 15598 62190 15650 62242
rect 20862 62190 20914 62242
rect 27694 62190 27746 62242
rect 30830 62190 30882 62242
rect 31278 62190 31330 62242
rect 37550 62190 37602 62242
rect 38558 62190 38610 62242
rect 41022 62190 41074 62242
rect 42478 62190 42530 62242
rect 46174 62190 46226 62242
rect 49534 62190 49586 62242
rect 51662 62190 51714 62242
rect 52894 62190 52946 62242
rect 55358 62190 55410 62242
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 20302 61742 20354 61794
rect 38222 61742 38274 61794
rect 43374 61742 43426 61794
rect 49198 61742 49250 61794
rect 56366 61742 56418 61794
rect 7534 61630 7586 61682
rect 12238 61630 12290 61682
rect 24558 61630 24610 61682
rect 35870 61630 35922 61682
rect 37438 61630 37490 61682
rect 52782 61630 52834 61682
rect 55022 61630 55074 61682
rect 21758 61518 21810 61570
rect 35646 61518 35698 61570
rect 38558 61518 38610 61570
rect 43374 61518 43426 61570
rect 53118 61518 53170 61570
rect 54350 61518 54402 61570
rect 55470 61518 55522 61570
rect 6414 61406 6466 61458
rect 6750 61406 6802 61458
rect 19966 61406 20018 61458
rect 20414 61406 20466 61458
rect 20638 61406 20690 61458
rect 22430 61406 22482 61458
rect 24894 61406 24946 61458
rect 32734 61406 32786 61458
rect 34414 61406 34466 61458
rect 34974 61406 35026 61458
rect 35982 61406 36034 61458
rect 36990 61406 37042 61458
rect 37214 61406 37266 61458
rect 37550 61406 37602 61458
rect 43710 61406 43762 61458
rect 49086 61406 49138 61458
rect 6190 61294 6242 61346
rect 6302 61294 6354 61346
rect 6862 61294 6914 61346
rect 7086 61294 7138 61346
rect 20190 61294 20242 61346
rect 20750 61294 20802 61346
rect 25006 61294 25058 61346
rect 25566 61294 25618 61346
rect 25902 61294 25954 61346
rect 32398 61294 32450 61346
rect 32622 61294 32674 61346
rect 34526 61294 34578 61346
rect 34750 61294 34802 61346
rect 35086 61294 35138 61346
rect 35198 61294 35250 61346
rect 38334 61294 38386 61346
rect 44942 61294 44994 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 7870 60958 7922 61010
rect 25454 60958 25506 61010
rect 26014 60958 26066 61010
rect 32286 60958 32338 61010
rect 37326 60958 37378 61010
rect 40014 60958 40066 61010
rect 42702 60958 42754 61010
rect 49086 60958 49138 61010
rect 49646 60958 49698 61010
rect 50990 60958 51042 61010
rect 57038 60958 57090 61010
rect 57934 60958 57986 61010
rect 6302 60846 6354 60898
rect 11006 60846 11058 60898
rect 13022 60846 13074 60898
rect 13246 60846 13298 60898
rect 17502 60846 17554 60898
rect 17950 60846 18002 60898
rect 18062 60846 18114 60898
rect 20974 60846 21026 60898
rect 27246 60846 27298 60898
rect 27806 60846 27858 60898
rect 29598 60846 29650 60898
rect 35422 60846 35474 60898
rect 36766 60846 36818 60898
rect 39118 60846 39170 60898
rect 54462 60846 54514 60898
rect 55806 60846 55858 60898
rect 57150 60846 57202 60898
rect 57374 60846 57426 60898
rect 2830 60734 2882 60786
rect 6750 60734 6802 60786
rect 7534 60734 7586 60786
rect 10782 60734 10834 60786
rect 11566 60734 11618 60786
rect 11902 60734 11954 60786
rect 12574 60734 12626 60786
rect 13358 60734 13410 60786
rect 17390 60734 17442 60786
rect 17726 60734 17778 60786
rect 21758 60734 21810 60786
rect 22654 60734 22706 60786
rect 25902 60734 25954 60786
rect 26238 60734 26290 60786
rect 27134 60734 27186 60786
rect 27470 60734 27522 60786
rect 27694 60734 27746 60786
rect 27918 60734 27970 60786
rect 28366 60734 28418 60786
rect 28926 60734 28978 60786
rect 31950 60734 32002 60786
rect 33406 60734 33458 60786
rect 34750 60734 34802 60786
rect 35870 60734 35922 60786
rect 36094 60734 36146 60786
rect 37774 60734 37826 60786
rect 39006 60734 39058 60786
rect 39902 60734 39954 60786
rect 41358 60734 41410 60786
rect 42478 60734 42530 60786
rect 48862 60734 48914 60786
rect 49310 60734 49362 60786
rect 49646 60734 49698 60786
rect 50094 60734 50146 60786
rect 51214 60734 51266 60786
rect 53006 60734 53058 60786
rect 53342 60734 53394 60786
rect 54686 60734 54738 60786
rect 56702 60734 56754 60786
rect 57710 60734 57762 60786
rect 3502 60622 3554 60674
rect 5630 60622 5682 60674
rect 11118 60622 11170 60674
rect 12686 60622 12738 60674
rect 13918 60622 13970 60674
rect 14254 60622 14306 60674
rect 18846 60622 18898 60674
rect 23214 60622 23266 60674
rect 28702 60622 28754 60674
rect 30046 60622 30098 60674
rect 30494 60622 30546 60674
rect 31614 60622 31666 60674
rect 33182 60622 33234 60674
rect 34078 60622 34130 60674
rect 34526 60622 34578 60674
rect 37886 60622 37938 60674
rect 38558 60622 38610 60674
rect 41918 60622 41970 60674
rect 49758 60622 49810 60674
rect 56030 60622 56082 60674
rect 18062 60510 18114 60562
rect 25230 60510 25282 60562
rect 25566 60510 25618 60562
rect 29934 60510 29986 60562
rect 41470 60510 41522 60562
rect 42814 60510 42866 60562
rect 56926 60510 56978 60562
rect 58046 60510 58098 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 6974 60174 7026 60226
rect 17614 60174 17666 60226
rect 18958 60174 19010 60226
rect 22654 60174 22706 60226
rect 28366 60174 28418 60226
rect 32510 60174 32562 60226
rect 34414 60174 34466 60226
rect 34750 60174 34802 60226
rect 44270 60174 44322 60226
rect 5854 60062 5906 60114
rect 9102 60062 9154 60114
rect 11230 60062 11282 60114
rect 11790 60062 11842 60114
rect 15710 60062 15762 60114
rect 17166 60062 17218 60114
rect 25454 60062 25506 60114
rect 27806 60062 27858 60114
rect 32062 60062 32114 60114
rect 34190 60062 34242 60114
rect 38670 60062 38722 60114
rect 42478 60062 42530 60114
rect 49870 60062 49922 60114
rect 54910 60062 54962 60114
rect 55246 60062 55298 60114
rect 6526 59950 6578 60002
rect 7086 59950 7138 60002
rect 7422 59950 7474 60002
rect 8430 59950 8482 60002
rect 11678 59950 11730 60002
rect 12462 59950 12514 60002
rect 12910 59950 12962 60002
rect 14142 59950 14194 60002
rect 15262 59950 15314 60002
rect 16494 59950 16546 60002
rect 16942 59950 16994 60002
rect 18846 59950 18898 60002
rect 19854 59950 19906 60002
rect 20190 59950 20242 60002
rect 23998 59950 24050 60002
rect 25902 59950 25954 60002
rect 26462 59950 26514 60002
rect 28030 59950 28082 60002
rect 29038 59950 29090 60002
rect 29374 59950 29426 60002
rect 31166 59950 31218 60002
rect 31390 59950 31442 60002
rect 32846 59950 32898 60002
rect 33630 59950 33682 60002
rect 40798 59950 40850 60002
rect 41694 59950 41746 60002
rect 47070 59950 47122 60002
rect 50990 59950 51042 60002
rect 51214 59950 51266 60002
rect 51662 59950 51714 60002
rect 51886 59950 51938 60002
rect 52110 59950 52162 60002
rect 58046 59950 58098 60002
rect 12014 59838 12066 59890
rect 13806 59838 13858 59890
rect 16158 59838 16210 59890
rect 16270 59838 16322 59890
rect 22990 59838 23042 59890
rect 23326 59838 23378 59890
rect 24894 59838 24946 59890
rect 26574 59838 26626 59890
rect 29262 59838 29314 59890
rect 32398 59838 32450 59890
rect 33070 59838 33122 59890
rect 33182 59838 33234 59890
rect 44158 59838 44210 59890
rect 47742 59838 47794 59890
rect 50206 59838 50258 59890
rect 57374 59838 57426 59890
rect 21982 59726 22034 59778
rect 22766 59726 22818 59778
rect 26014 59726 26066 59778
rect 27470 59726 27522 59778
rect 30382 59726 30434 59778
rect 30718 59726 30770 59778
rect 32510 59726 32562 59778
rect 40014 59726 40066 59778
rect 40462 59726 40514 59778
rect 40686 59726 40738 59778
rect 40910 59726 40962 59778
rect 50542 59726 50594 59778
rect 51102 59726 51154 59778
rect 51998 59726 52050 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 7646 59390 7698 59442
rect 11342 59390 11394 59442
rect 15038 59390 15090 59442
rect 15150 59390 15202 59442
rect 15710 59390 15762 59442
rect 16718 59390 16770 59442
rect 27022 59390 27074 59442
rect 42254 59390 42306 59442
rect 48078 59390 48130 59442
rect 48862 59390 48914 59442
rect 48974 59390 49026 59442
rect 49534 59390 49586 59442
rect 50430 59390 50482 59442
rect 54686 59390 54738 59442
rect 56030 59390 56082 59442
rect 56814 59390 56866 59442
rect 7534 59278 7586 59330
rect 7758 59278 7810 59330
rect 8206 59278 8258 59330
rect 17614 59278 17666 59330
rect 35646 59278 35698 59330
rect 41470 59278 41522 59330
rect 42366 59278 42418 59330
rect 43038 59278 43090 59330
rect 48190 59278 48242 59330
rect 56926 59278 56978 59330
rect 12238 59166 12290 59218
rect 14478 59166 14530 59218
rect 14926 59166 14978 59218
rect 15934 59166 15986 59218
rect 16494 59166 16546 59218
rect 17726 59166 17778 59218
rect 27358 59166 27410 59218
rect 36542 59166 36594 59218
rect 37102 59166 37154 59218
rect 39902 59166 39954 59218
rect 40798 59166 40850 59218
rect 41246 59166 41298 59218
rect 42030 59166 42082 59218
rect 42142 59166 42194 59218
rect 42590 59166 42642 59218
rect 42926 59166 42978 59218
rect 43262 59166 43314 59218
rect 45278 59166 45330 59218
rect 49310 59166 49362 59218
rect 49422 59166 49474 59218
rect 49982 59166 50034 59218
rect 51438 59166 51490 59218
rect 56590 59166 56642 59218
rect 58158 59166 58210 59218
rect 1822 59054 1874 59106
rect 12798 59054 12850 59106
rect 18062 59054 18114 59106
rect 27806 59054 27858 59106
rect 30942 59054 30994 59106
rect 32286 59054 32338 59106
rect 39454 59054 39506 59106
rect 40350 59054 40402 59106
rect 41022 59054 41074 59106
rect 45726 59054 45778 59106
rect 49646 59054 49698 59106
rect 52110 59054 52162 59106
rect 54238 59054 54290 59106
rect 55582 59054 55634 59106
rect 57710 59054 57762 59106
rect 35758 58942 35810 58994
rect 37214 58942 37266 58994
rect 44942 58942 44994 58994
rect 45278 58942 45330 58994
rect 55582 58942 55634 58994
rect 56142 58942 56194 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 16382 58606 16434 58658
rect 16718 58606 16770 58658
rect 25790 58606 25842 58658
rect 26126 58606 26178 58658
rect 35982 58606 36034 58658
rect 43150 58606 43202 58658
rect 52110 58606 52162 58658
rect 4846 58494 4898 58546
rect 10222 58494 10274 58546
rect 12350 58494 12402 58546
rect 14478 58494 14530 58546
rect 27358 58494 27410 58546
rect 39230 58494 39282 58546
rect 41358 58494 41410 58546
rect 41806 58494 41858 58546
rect 44830 58494 44882 58546
rect 46958 58494 47010 58546
rect 48190 58494 48242 58546
rect 51998 58494 52050 58546
rect 54686 58494 54738 58546
rect 58270 58494 58322 58546
rect 2270 58382 2322 58434
rect 4174 58382 4226 58434
rect 4286 58382 4338 58434
rect 5630 58382 5682 58434
rect 11790 58382 11842 58434
rect 25678 58382 25730 58434
rect 26686 58382 26738 58434
rect 27806 58382 27858 58434
rect 38558 58382 38610 58434
rect 43262 58382 43314 58434
rect 47742 58382 47794 58434
rect 53006 58382 53058 58434
rect 1710 58270 1762 58322
rect 3838 58270 3890 58322
rect 10670 58270 10722 58322
rect 13470 58270 13522 58322
rect 15822 58270 15874 58322
rect 16158 58270 16210 58322
rect 25342 58270 25394 58322
rect 28142 58270 28194 58322
rect 29822 58270 29874 58322
rect 30494 58270 30546 58322
rect 36318 58270 36370 58322
rect 43150 58270 43202 58322
rect 3950 58158 4002 58210
rect 5742 58158 5794 58210
rect 5966 58158 6018 58210
rect 13806 58158 13858 58210
rect 15374 58158 15426 58210
rect 25454 58158 25506 58210
rect 26126 58158 26178 58210
rect 29934 58158 29986 58210
rect 30046 58158 30098 58210
rect 30606 58158 30658 58210
rect 30830 58158 30882 58210
rect 36094 58158 36146 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 6862 57822 6914 57874
rect 9886 57822 9938 57874
rect 10558 57822 10610 57874
rect 20526 57822 20578 57874
rect 25342 57822 25394 57874
rect 28030 57822 28082 57874
rect 44942 57822 44994 57874
rect 51662 57822 51714 57874
rect 52558 57822 52610 57874
rect 2494 57710 2546 57762
rect 4958 57710 5010 57762
rect 13806 57710 13858 57762
rect 19630 57710 19682 57762
rect 19742 57710 19794 57762
rect 22878 57710 22930 57762
rect 23998 57710 24050 57762
rect 27694 57710 27746 57762
rect 30046 57710 30098 57762
rect 36430 57710 36482 57762
rect 39006 57710 39058 57762
rect 43262 57710 43314 57762
rect 1822 57598 1874 57650
rect 5630 57598 5682 57650
rect 6302 57598 6354 57650
rect 7982 57598 8034 57650
rect 8318 57598 8370 57650
rect 8542 57598 8594 57650
rect 9438 57598 9490 57650
rect 10110 57598 10162 57650
rect 10334 57598 10386 57650
rect 10670 57598 10722 57650
rect 13918 57598 13970 57650
rect 19406 57598 19458 57650
rect 20078 57598 20130 57650
rect 20302 57598 20354 57650
rect 20750 57598 20802 57650
rect 22766 57598 22818 57650
rect 23662 57598 23714 57650
rect 24670 57598 24722 57650
rect 25678 57598 25730 57650
rect 26462 57598 26514 57650
rect 27022 57598 27074 57650
rect 28254 57598 28306 57650
rect 30270 57598 30322 57650
rect 30942 57598 30994 57650
rect 32398 57598 32450 57650
rect 37662 57598 37714 57650
rect 42142 57598 42194 57650
rect 44494 57598 44546 57650
rect 51438 57598 51490 57650
rect 51998 57598 52050 57650
rect 4622 57486 4674 57538
rect 5854 57486 5906 57538
rect 8094 57486 8146 57538
rect 9998 57486 10050 57538
rect 13358 57486 13410 57538
rect 23774 57486 23826 57538
rect 31614 57486 31666 57538
rect 32062 57486 32114 57538
rect 33182 57486 33234 57538
rect 36206 57486 36258 57538
rect 42590 57486 42642 57538
rect 43150 57486 43202 57538
rect 51102 57486 51154 57538
rect 51550 57486 51602 57538
rect 6526 57374 6578 57426
rect 13806 57374 13858 57426
rect 22654 57374 22706 57426
rect 32398 57374 32450 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 12238 57038 12290 57090
rect 24670 57038 24722 57090
rect 27246 57038 27298 57090
rect 29822 57038 29874 57090
rect 43598 57038 43650 57090
rect 4510 56926 4562 56978
rect 6078 56926 6130 56978
rect 7422 56926 7474 56978
rect 9550 56926 9602 56978
rect 10670 56926 10722 56978
rect 14142 56926 14194 56978
rect 15038 56926 15090 56978
rect 16158 56926 16210 56978
rect 19406 56926 19458 56978
rect 20190 56926 20242 56978
rect 22094 56926 22146 56978
rect 24222 56926 24274 56978
rect 29934 56926 29986 56978
rect 31614 56926 31666 56978
rect 33742 56926 33794 56978
rect 34974 56926 35026 56978
rect 36318 56926 36370 56978
rect 42366 56926 42418 56978
rect 42702 56926 42754 56978
rect 47070 56926 47122 56978
rect 50430 56926 50482 56978
rect 55358 56926 55410 56978
rect 4622 56814 4674 56866
rect 5070 56814 5122 56866
rect 5518 56814 5570 56866
rect 5966 56814 6018 56866
rect 6750 56814 6802 56866
rect 10558 56814 10610 56866
rect 16494 56814 16546 56866
rect 20302 56814 20354 56866
rect 20750 56814 20802 56866
rect 21310 56814 21362 56866
rect 25454 56814 25506 56866
rect 26126 56814 26178 56866
rect 26686 56814 26738 56866
rect 30158 56814 30210 56866
rect 30830 56814 30882 56866
rect 34526 56814 34578 56866
rect 35982 56814 36034 56866
rect 37102 56814 37154 56866
rect 37326 56814 37378 56866
rect 37998 56814 38050 56866
rect 42254 56814 42306 56866
rect 42926 56814 42978 56866
rect 49982 56814 50034 56866
rect 4398 56702 4450 56754
rect 9886 56702 9938 56754
rect 12014 56702 12066 56754
rect 13806 56702 13858 56754
rect 13918 56702 13970 56754
rect 14254 56702 14306 56754
rect 15150 56702 15202 56754
rect 17278 56702 17330 56754
rect 19854 56702 19906 56754
rect 24782 56702 24834 56754
rect 25118 56702 25170 56754
rect 26798 56702 26850 56754
rect 27134 56702 27186 56754
rect 36094 56702 36146 56754
rect 36430 56702 36482 56754
rect 42478 56702 42530 56754
rect 43262 56702 43314 56754
rect 43486 56702 43538 56754
rect 49198 56702 49250 56754
rect 55582 56702 55634 56754
rect 6190 56590 6242 56642
rect 12574 56590 12626 56642
rect 14030 56590 14082 56642
rect 14702 56590 14754 56642
rect 14926 56590 14978 56642
rect 20078 56590 20130 56642
rect 24670 56590 24722 56642
rect 27694 56590 27746 56642
rect 55358 56590 55410 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 8654 56254 8706 56306
rect 8766 56254 8818 56306
rect 9774 56254 9826 56306
rect 10782 56254 10834 56306
rect 11230 56254 11282 56306
rect 12126 56254 12178 56306
rect 13694 56254 13746 56306
rect 22654 56254 22706 56306
rect 28478 56254 28530 56306
rect 36542 56254 36594 56306
rect 46958 56254 47010 56306
rect 48190 56254 48242 56306
rect 48862 56254 48914 56306
rect 49982 56254 50034 56306
rect 54238 56254 54290 56306
rect 8318 56142 8370 56194
rect 12910 56142 12962 56194
rect 13134 56142 13186 56194
rect 13358 56142 13410 56194
rect 13470 56142 13522 56194
rect 13918 56142 13970 56194
rect 14030 56142 14082 56194
rect 16046 56142 16098 56194
rect 17950 56142 18002 56194
rect 19070 56142 19122 56194
rect 20302 56142 20354 56194
rect 23886 56142 23938 56194
rect 31838 56142 31890 56194
rect 32510 56142 32562 56194
rect 35198 56142 35250 56194
rect 35646 56142 35698 56194
rect 48750 56142 48802 56194
rect 51662 56142 51714 56194
rect 8542 56030 8594 56082
rect 10222 56030 10274 56082
rect 10446 56030 10498 56082
rect 11566 56030 11618 56082
rect 12462 56030 12514 56082
rect 12798 56030 12850 56082
rect 14254 56030 14306 56082
rect 14590 56030 14642 56082
rect 15150 56030 15202 56082
rect 22990 56030 23042 56082
rect 32286 56030 32338 56082
rect 33630 56030 33682 56082
rect 34190 56030 34242 56082
rect 35534 56030 35586 56082
rect 37214 56030 37266 56082
rect 38222 56030 38274 56082
rect 39006 56030 39058 56082
rect 47070 56030 47122 56082
rect 47182 56030 47234 56082
rect 47630 56030 47682 56082
rect 48078 56030 48130 56082
rect 50318 56030 50370 56082
rect 50878 56030 50930 56082
rect 54910 56030 54962 56082
rect 4622 55918 4674 55970
rect 5182 55918 5234 55970
rect 15262 55918 15314 55970
rect 17838 55918 17890 55970
rect 18174 55918 18226 55970
rect 18734 55918 18786 55970
rect 20750 55918 20802 55970
rect 24446 55918 24498 55970
rect 25342 55918 25394 55970
rect 31390 55918 31442 55970
rect 45502 55918 45554 55970
rect 47854 55918 47906 55970
rect 53790 55918 53842 55970
rect 55134 55918 55186 55970
rect 30942 55806 30994 55858
rect 31390 55806 31442 55858
rect 45614 55806 45666 55858
rect 55582 55806 55634 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 4846 55470 4898 55522
rect 32286 55470 32338 55522
rect 35198 55470 35250 55522
rect 43150 55470 43202 55522
rect 11790 55358 11842 55410
rect 23550 55358 23602 55410
rect 23774 55358 23826 55410
rect 33070 55358 33122 55410
rect 34862 55358 34914 55410
rect 40462 55358 40514 55410
rect 41582 55358 41634 55410
rect 42142 55358 42194 55410
rect 45614 55358 45666 55410
rect 47742 55358 47794 55410
rect 52782 55358 52834 55410
rect 55582 55358 55634 55410
rect 57710 55358 57762 55410
rect 2942 55246 2994 55298
rect 3502 55246 3554 55298
rect 3950 55246 4002 55298
rect 4510 55246 4562 55298
rect 11006 55246 11058 55298
rect 11342 55246 11394 55298
rect 14478 55246 14530 55298
rect 23886 55246 23938 55298
rect 28366 55246 28418 55298
rect 29262 55246 29314 55298
rect 30158 55246 30210 55298
rect 30942 55246 30994 55298
rect 31726 55246 31778 55298
rect 32958 55246 33010 55298
rect 33854 55246 33906 55298
rect 34750 55246 34802 55298
rect 37662 55246 37714 55298
rect 41470 55246 41522 55298
rect 42366 55246 42418 55298
rect 42814 55246 42866 55298
rect 44942 55246 44994 55298
rect 53342 55246 53394 55298
rect 54910 55246 54962 55298
rect 58158 55246 58210 55298
rect 3278 55134 3330 55186
rect 4958 55134 5010 55186
rect 29374 55134 29426 55186
rect 30718 55134 30770 55186
rect 31390 55134 31442 55186
rect 32286 55134 32338 55186
rect 32398 55134 32450 55186
rect 38334 55134 38386 55186
rect 40798 55134 40850 55186
rect 49982 55134 50034 55186
rect 3054 55022 3106 55074
rect 3838 55022 3890 55074
rect 4062 55022 4114 55074
rect 4846 55022 4898 55074
rect 11118 55022 11170 55074
rect 12686 55022 12738 55074
rect 13582 55022 13634 55074
rect 14590 55022 14642 55074
rect 18398 55022 18450 55074
rect 27694 55022 27746 55074
rect 27806 55022 27858 55074
rect 27918 55022 27970 55074
rect 30158 55022 30210 55074
rect 31502 55022 31554 55074
rect 43038 55022 43090 55074
rect 44270 55022 44322 55074
rect 49198 55022 49250 55074
rect 49534 55022 49586 55074
rect 50318 55022 50370 55074
rect 52782 55022 52834 55074
rect 52894 55022 52946 55074
rect 53118 55022 53170 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 5070 54686 5122 54738
rect 11006 54686 11058 54738
rect 29486 54686 29538 54738
rect 39566 54686 39618 54738
rect 41022 54686 41074 54738
rect 41582 54686 41634 54738
rect 41694 54686 41746 54738
rect 41806 54686 41858 54738
rect 42478 54686 42530 54738
rect 45502 54686 45554 54738
rect 45950 54686 46002 54738
rect 46622 54686 46674 54738
rect 51886 54686 51938 54738
rect 2494 54574 2546 54626
rect 5406 54574 5458 54626
rect 14590 54574 14642 54626
rect 26686 54574 26738 54626
rect 27022 54574 27074 54626
rect 31502 54574 31554 54626
rect 31950 54574 32002 54626
rect 39454 54574 39506 54626
rect 42366 54574 42418 54626
rect 51214 54574 51266 54626
rect 55806 54574 55858 54626
rect 1822 54462 1874 54514
rect 4958 54462 5010 54514
rect 5182 54462 5234 54514
rect 11342 54462 11394 54514
rect 14254 54462 14306 54514
rect 14478 54462 14530 54514
rect 14814 54462 14866 54514
rect 15150 54462 15202 54514
rect 15486 54462 15538 54514
rect 18286 54462 18338 54514
rect 27246 54462 27298 54514
rect 27582 54462 27634 54514
rect 28142 54462 28194 54514
rect 30830 54462 30882 54514
rect 39790 54462 39842 54514
rect 40014 54462 40066 54514
rect 41470 54462 41522 54514
rect 42030 54462 42082 54514
rect 46062 54462 46114 54514
rect 46398 54462 46450 54514
rect 46622 54462 46674 54514
rect 50878 54462 50930 54514
rect 51662 54462 51714 54514
rect 56478 54462 56530 54514
rect 56814 54462 56866 54514
rect 57150 54462 57202 54514
rect 4622 54350 4674 54402
rect 16718 54350 16770 54402
rect 26798 54350 26850 54402
rect 28478 54350 28530 54402
rect 28926 54350 28978 54402
rect 29150 54350 29202 54402
rect 30606 54350 30658 54402
rect 46846 54350 46898 54402
rect 47182 54350 47234 54402
rect 55134 54350 55186 54402
rect 55918 54350 55970 54402
rect 56702 54350 56754 54402
rect 54574 54238 54626 54290
rect 54910 54238 54962 54290
rect 56030 54238 56082 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 8990 53902 9042 53954
rect 23326 53902 23378 53954
rect 29374 53902 29426 53954
rect 29710 53902 29762 53954
rect 36318 53902 36370 53954
rect 52670 53902 52722 53954
rect 2942 53790 2994 53842
rect 18734 53790 18786 53842
rect 22318 53790 22370 53842
rect 24110 53790 24162 53842
rect 26014 53790 26066 53842
rect 28142 53790 28194 53842
rect 29150 53790 29202 53842
rect 36094 53790 36146 53842
rect 37102 53790 37154 53842
rect 40014 53790 40066 53842
rect 53006 53790 53058 53842
rect 53902 53790 53954 53842
rect 56030 53790 56082 53842
rect 58158 53790 58210 53842
rect 3390 53678 3442 53730
rect 3838 53678 3890 53730
rect 4622 53678 4674 53730
rect 5070 53678 5122 53730
rect 7870 53678 7922 53730
rect 8430 53678 8482 53730
rect 8878 53678 8930 53730
rect 17838 53678 17890 53730
rect 18398 53678 18450 53730
rect 19854 53678 19906 53730
rect 19966 53678 20018 53730
rect 23886 53678 23938 53730
rect 24782 53678 24834 53730
rect 25230 53678 25282 53730
rect 34526 53678 34578 53730
rect 35982 53678 36034 53730
rect 37326 53678 37378 53730
rect 37998 53678 38050 53730
rect 39902 53678 39954 53730
rect 40574 53678 40626 53730
rect 51438 53678 51490 53730
rect 54910 53678 54962 53730
rect 55246 53678 55298 53730
rect 4286 53566 4338 53618
rect 4398 53566 4450 53618
rect 7086 53566 7138 53618
rect 7422 53566 7474 53618
rect 7646 53566 7698 53618
rect 10334 53566 10386 53618
rect 17950 53566 18002 53618
rect 19070 53566 19122 53618
rect 20638 53566 20690 53618
rect 22654 53566 22706 53618
rect 23102 53566 23154 53618
rect 24334 53566 24386 53618
rect 30382 53566 30434 53618
rect 39566 53566 39618 53618
rect 40910 53566 40962 53618
rect 41246 53566 41298 53618
rect 41582 53566 41634 53618
rect 41694 53566 41746 53618
rect 54238 53566 54290 53618
rect 54798 53566 54850 53618
rect 7198 53454 7250 53506
rect 8318 53454 8370 53506
rect 8542 53454 8594 53506
rect 8990 53454 9042 53506
rect 10670 53454 10722 53506
rect 18174 53454 18226 53506
rect 18622 53454 18674 53506
rect 18846 53454 18898 53506
rect 19630 53454 19682 53506
rect 20078 53454 20130 53506
rect 20302 53454 20354 53506
rect 20526 53454 20578 53506
rect 22430 53454 22482 53506
rect 23214 53454 23266 53506
rect 30046 53454 30098 53506
rect 33182 53454 33234 53506
rect 40126 53454 40178 53506
rect 41022 53454 41074 53506
rect 41358 53454 41410 53506
rect 51662 53454 51714 53506
rect 52782 53454 52834 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 14590 53118 14642 53170
rect 23998 53118 24050 53170
rect 24670 53118 24722 53170
rect 25342 53118 25394 53170
rect 31278 53118 31330 53170
rect 36430 53118 36482 53170
rect 45838 53118 45890 53170
rect 46622 53118 46674 53170
rect 46846 53118 46898 53170
rect 47518 53118 47570 53170
rect 47966 53118 48018 53170
rect 55022 53118 55074 53170
rect 5966 53006 6018 53058
rect 8542 53006 8594 53058
rect 12014 53006 12066 53058
rect 12574 53006 12626 53058
rect 14814 53006 14866 53058
rect 18174 53006 18226 53058
rect 21422 53006 21474 53058
rect 23886 53006 23938 53058
rect 36206 53006 36258 53058
rect 36654 53006 36706 53058
rect 51550 53006 51602 53058
rect 5182 52894 5234 52946
rect 8430 52894 8482 52946
rect 8654 52894 8706 52946
rect 8990 52894 9042 52946
rect 10334 52894 10386 52946
rect 11566 52894 11618 52946
rect 12350 52894 12402 52946
rect 12686 52894 12738 52946
rect 14926 52894 14978 52946
rect 17502 52894 17554 52946
rect 20638 52894 20690 52946
rect 24222 52894 24274 52946
rect 31614 52894 31666 52946
rect 32174 52894 32226 52946
rect 33742 52894 33794 52946
rect 34414 52894 34466 52946
rect 35646 52894 35698 52946
rect 35982 52894 36034 52946
rect 36766 52894 36818 52946
rect 42478 52894 42530 52946
rect 46398 52894 46450 52946
rect 47070 52894 47122 52946
rect 50766 52894 50818 52946
rect 54126 52894 54178 52946
rect 54462 52894 54514 52946
rect 58158 52894 58210 52946
rect 8094 52782 8146 52834
rect 9774 52782 9826 52834
rect 10110 52782 10162 52834
rect 10670 52782 10722 52834
rect 11118 52782 11170 52834
rect 13694 52782 13746 52834
rect 20302 52782 20354 52834
rect 23550 52782 23602 52834
rect 31950 52782 32002 52834
rect 33518 52782 33570 52834
rect 41022 52782 41074 52834
rect 43262 52782 43314 52834
rect 45390 52782 45442 52834
rect 46510 52782 46562 52834
rect 53678 52782 53730 52834
rect 57374 52782 57426 52834
rect 57598 52782 57650 52834
rect 13134 52670 13186 52722
rect 32510 52670 32562 52722
rect 45614 52670 45666 52722
rect 46174 52670 46226 52722
rect 47294 52670 47346 52722
rect 47630 52670 47682 52722
rect 54014 52670 54066 52722
rect 54350 52670 54402 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 8766 52334 8818 52386
rect 15710 52334 15762 52386
rect 16158 52334 16210 52386
rect 16494 52334 16546 52386
rect 20414 52334 20466 52386
rect 20750 52334 20802 52386
rect 36094 52334 36146 52386
rect 55918 52334 55970 52386
rect 56142 52334 56194 52386
rect 56254 52334 56306 52386
rect 7310 52222 7362 52274
rect 8206 52222 8258 52274
rect 12350 52222 12402 52274
rect 18510 52222 18562 52274
rect 19406 52222 19458 52274
rect 20190 52222 20242 52274
rect 21534 52222 21586 52274
rect 24558 52222 24610 52274
rect 32398 52222 32450 52274
rect 33630 52222 33682 52274
rect 35982 52222 36034 52274
rect 39454 52222 39506 52274
rect 43262 52222 43314 52274
rect 46734 52222 46786 52274
rect 47630 52222 47682 52274
rect 51214 52222 51266 52274
rect 51774 52222 51826 52274
rect 4622 52110 4674 52162
rect 7982 52110 8034 52162
rect 8654 52110 8706 52162
rect 9662 52110 9714 52162
rect 10222 52110 10274 52162
rect 12910 52110 12962 52162
rect 13582 52110 13634 52162
rect 13918 52110 13970 52162
rect 14478 52110 14530 52162
rect 14814 52110 14866 52162
rect 15038 52110 15090 52162
rect 15262 52110 15314 52162
rect 15934 52110 15986 52162
rect 19182 52110 19234 52162
rect 23102 52110 23154 52162
rect 30942 52110 30994 52162
rect 31950 52110 32002 52162
rect 32286 52110 32338 52162
rect 32734 52110 32786 52162
rect 33294 52110 33346 52162
rect 35646 52110 35698 52162
rect 38894 52110 38946 52162
rect 43822 52110 43874 52162
rect 46622 52110 46674 52162
rect 50542 52110 50594 52162
rect 50990 52110 51042 52162
rect 54126 52110 54178 52162
rect 8766 51998 8818 52050
rect 9998 51998 10050 52050
rect 11454 51998 11506 52050
rect 24334 51998 24386 52050
rect 30718 51998 30770 52050
rect 33742 51998 33794 52050
rect 37662 51998 37714 52050
rect 43150 51998 43202 52050
rect 44158 51998 44210 52050
rect 47070 51998 47122 52050
rect 47294 51998 47346 52050
rect 49758 51998 49810 52050
rect 11790 51886 11842 51938
rect 12238 51886 12290 51938
rect 12462 51886 12514 51938
rect 22542 51886 22594 51938
rect 37998 51886 38050 51938
rect 43374 51886 43426 51938
rect 46846 51886 46898 51938
rect 54462 51886 54514 51938
rect 56254 51886 56306 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 12910 51550 12962 51602
rect 13134 51550 13186 51602
rect 13358 51550 13410 51602
rect 32510 51550 32562 51602
rect 36318 51550 36370 51602
rect 43262 51550 43314 51602
rect 47182 51550 47234 51602
rect 48302 51550 48354 51602
rect 48862 51550 48914 51602
rect 51886 51550 51938 51602
rect 52782 51550 52834 51602
rect 55918 51550 55970 51602
rect 56702 51550 56754 51602
rect 3390 51438 3442 51490
rect 5406 51438 5458 51490
rect 13470 51438 13522 51490
rect 15038 51438 15090 51490
rect 37326 51438 37378 51490
rect 38670 51438 38722 51490
rect 41022 51438 41074 51490
rect 41582 51438 41634 51490
rect 41694 51438 41746 51490
rect 48750 51438 48802 51490
rect 53230 51438 53282 51490
rect 55470 51438 55522 51490
rect 3278 51326 3330 51378
rect 3614 51326 3666 51378
rect 3838 51326 3890 51378
rect 4174 51326 4226 51378
rect 4398 51326 4450 51378
rect 5070 51326 5122 51378
rect 5742 51326 5794 51378
rect 14590 51326 14642 51378
rect 15262 51326 15314 51378
rect 28478 51326 28530 51378
rect 29262 51326 29314 51378
rect 30046 51326 30098 51378
rect 36206 51326 36258 51378
rect 36766 51326 36818 51378
rect 37998 51326 38050 51378
rect 43710 51326 43762 51378
rect 46958 51326 47010 51378
rect 47294 51326 47346 51378
rect 47630 51326 47682 51378
rect 52110 51326 52162 51378
rect 52446 51326 52498 51378
rect 55134 51326 55186 51378
rect 55358 51326 55410 51378
rect 56478 51326 56530 51378
rect 56814 51326 56866 51378
rect 57038 51326 57090 51378
rect 4286 51214 4338 51266
rect 5518 51214 5570 51266
rect 15150 51214 15202 51266
rect 29710 51214 29762 51266
rect 37774 51214 37826 51266
rect 42254 51214 42306 51266
rect 44382 51214 44434 51266
rect 46510 51214 46562 51266
rect 47854 51214 47906 51266
rect 48190 51214 48242 51266
rect 28590 51102 28642 51154
rect 29822 51102 29874 51154
rect 40910 51102 40962 51154
rect 41246 51102 41298 51154
rect 41694 51102 41746 51154
rect 51774 51102 51826 51154
rect 53118 51102 53170 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 5070 50766 5122 50818
rect 5742 50766 5794 50818
rect 14366 50766 14418 50818
rect 41806 50766 41858 50818
rect 4622 50654 4674 50706
rect 9326 50654 9378 50706
rect 11566 50654 11618 50706
rect 28366 50654 28418 50706
rect 29710 50654 29762 50706
rect 33182 50654 33234 50706
rect 35198 50654 35250 50706
rect 36318 50654 36370 50706
rect 38558 50654 38610 50706
rect 40686 50654 40738 50706
rect 44942 50654 44994 50706
rect 56030 50654 56082 50706
rect 58158 50654 58210 50706
rect 1822 50542 1874 50594
rect 4958 50542 5010 50594
rect 5630 50542 5682 50594
rect 9214 50542 9266 50594
rect 9886 50542 9938 50594
rect 25454 50542 25506 50594
rect 29486 50542 29538 50594
rect 30158 50542 30210 50594
rect 30382 50542 30434 50594
rect 30718 50542 30770 50594
rect 30942 50542 30994 50594
rect 32286 50542 32338 50594
rect 32510 50542 32562 50594
rect 33294 50542 33346 50594
rect 35086 50542 35138 50594
rect 41470 50542 41522 50594
rect 41918 50542 41970 50594
rect 42142 50542 42194 50594
rect 42254 50542 42306 50594
rect 42814 50542 42866 50594
rect 44830 50542 44882 50594
rect 45502 50542 45554 50594
rect 45838 50542 45890 50594
rect 46734 50542 46786 50594
rect 47182 50542 47234 50594
rect 47406 50542 47458 50594
rect 55246 50542 55298 50594
rect 2494 50430 2546 50482
rect 5742 50430 5794 50482
rect 8878 50430 8930 50482
rect 10782 50430 10834 50482
rect 11118 50430 11170 50482
rect 14030 50430 14082 50482
rect 19630 50430 19682 50482
rect 25118 50430 25170 50482
rect 26238 50430 26290 50482
rect 30606 50430 30658 50482
rect 47854 50430 47906 50482
rect 13694 50318 13746 50370
rect 14254 50318 14306 50370
rect 19742 50318 19794 50370
rect 45054 50318 45106 50370
rect 46958 50318 47010 50370
rect 47070 50318 47122 50370
rect 54910 50318 54962 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 4510 49982 4562 50034
rect 9438 49982 9490 50034
rect 28478 49982 28530 50034
rect 29374 49982 29426 50034
rect 29486 49982 29538 50034
rect 29934 49982 29986 50034
rect 30158 49982 30210 50034
rect 30494 49982 30546 50034
rect 35422 49982 35474 50034
rect 41022 49982 41074 50034
rect 50878 49982 50930 50034
rect 51102 49982 51154 50034
rect 4062 49870 4114 49922
rect 9662 49870 9714 49922
rect 10222 49870 10274 49922
rect 19294 49870 19346 49922
rect 20414 49870 20466 49922
rect 21534 49870 21586 49922
rect 28366 49870 28418 49922
rect 34078 49870 34130 49922
rect 37774 49870 37826 49922
rect 39342 49870 39394 49922
rect 41918 49870 41970 49922
rect 47294 49870 47346 49922
rect 50766 49870 50818 49922
rect 52222 49870 52274 49922
rect 3390 49758 3442 49810
rect 3950 49758 4002 49810
rect 4286 49758 4338 49810
rect 4734 49758 4786 49810
rect 4846 49758 4898 49810
rect 8654 49758 8706 49810
rect 8878 49758 8930 49810
rect 9774 49758 9826 49810
rect 9998 49758 10050 49810
rect 10334 49758 10386 49810
rect 12686 49758 12738 49810
rect 13246 49758 13298 49810
rect 14366 49758 14418 49810
rect 14814 49758 14866 49810
rect 19182 49758 19234 49810
rect 20302 49758 20354 49810
rect 21198 49758 21250 49810
rect 21422 49758 21474 49810
rect 23774 49758 23826 49810
rect 28702 49758 28754 49810
rect 28814 49758 28866 49810
rect 29262 49758 29314 49810
rect 29822 49758 29874 49810
rect 31502 49758 31554 49810
rect 32062 49758 32114 49810
rect 33406 49758 33458 49810
rect 35086 49758 35138 49810
rect 38670 49758 38722 49810
rect 41246 49758 41298 49810
rect 41358 49758 41410 49810
rect 41470 49758 41522 49810
rect 51998 49758 52050 49810
rect 52670 49758 52722 49810
rect 5406 49646 5458 49698
rect 7982 49646 8034 49698
rect 12350 49646 12402 49698
rect 13918 49646 13970 49698
rect 20526 49646 20578 49698
rect 23662 49646 23714 49698
rect 31166 49646 31218 49698
rect 32398 49646 32450 49698
rect 33742 49646 33794 49698
rect 34862 49646 34914 49698
rect 37214 49646 37266 49698
rect 41806 49646 41858 49698
rect 42142 49646 42194 49698
rect 49870 49646 49922 49698
rect 50430 49646 50482 49698
rect 51662 49646 51714 49698
rect 52446 49646 52498 49698
rect 19294 49534 19346 49586
rect 21534 49534 21586 49586
rect 23438 49534 23490 49586
rect 47406 49534 47458 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 33294 49198 33346 49250
rect 53006 49198 53058 49250
rect 8878 49086 8930 49138
rect 10222 49086 10274 49138
rect 16270 49086 16322 49138
rect 19518 49086 19570 49138
rect 22542 49086 22594 49138
rect 23662 49086 23714 49138
rect 25790 49086 25842 49138
rect 32734 49086 32786 49138
rect 32958 49086 33010 49138
rect 33742 49086 33794 49138
rect 42142 49086 42194 49138
rect 46734 49086 46786 49138
rect 48862 49086 48914 49138
rect 50766 49086 50818 49138
rect 58158 49086 58210 49138
rect 6078 48974 6130 49026
rect 9102 48974 9154 49026
rect 9662 48974 9714 49026
rect 15038 48974 15090 49026
rect 15598 48974 15650 49026
rect 16718 48974 16770 49026
rect 21982 48974 22034 49026
rect 22990 48974 23042 49026
rect 31502 48974 31554 49026
rect 32174 48974 32226 49026
rect 32398 48974 32450 49026
rect 41918 48974 41970 49026
rect 42030 48974 42082 49026
rect 42254 48974 42306 49026
rect 42814 48974 42866 49026
rect 49646 48974 49698 49026
rect 50654 48974 50706 49026
rect 51550 48974 51602 49026
rect 52782 48974 52834 49026
rect 53230 48974 53282 49026
rect 54126 48974 54178 49026
rect 54462 48974 54514 49026
rect 54910 48974 54962 49026
rect 55246 48974 55298 49026
rect 6750 48862 6802 48914
rect 9326 48862 9378 48914
rect 9550 48862 9602 48914
rect 11118 48862 11170 48914
rect 17390 48862 17442 48914
rect 20078 48862 20130 48914
rect 20190 48862 20242 48914
rect 20414 48862 20466 48914
rect 20638 48862 20690 48914
rect 21422 48862 21474 48914
rect 43150 48862 43202 48914
rect 56030 48862 56082 48914
rect 11230 48750 11282 48802
rect 11342 48750 11394 48802
rect 21310 48750 21362 48802
rect 21534 48750 21586 48802
rect 42366 48750 42418 48802
rect 43038 48750 43090 48802
rect 50990 48750 51042 48802
rect 52110 48750 52162 48802
rect 53118 48750 53170 48802
rect 53902 48750 53954 48802
rect 54686 48750 54738 48802
rect 54798 48750 54850 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 8318 48414 8370 48466
rect 8430 48414 8482 48466
rect 8542 48414 8594 48466
rect 19070 48414 19122 48466
rect 22094 48414 22146 48466
rect 24446 48414 24498 48466
rect 27358 48414 27410 48466
rect 32510 48414 32562 48466
rect 41694 48414 41746 48466
rect 42478 48414 42530 48466
rect 55918 48414 55970 48466
rect 4846 48302 4898 48354
rect 6190 48302 6242 48354
rect 8094 48302 8146 48354
rect 8878 48302 8930 48354
rect 10558 48302 10610 48354
rect 13582 48302 13634 48354
rect 15262 48302 15314 48354
rect 15710 48302 15762 48354
rect 20414 48302 20466 48354
rect 23662 48302 23714 48354
rect 28366 48302 28418 48354
rect 37214 48302 37266 48354
rect 42366 48302 42418 48354
rect 43374 48302 43426 48354
rect 53006 48302 53058 48354
rect 55470 48302 55522 48354
rect 55694 48302 55746 48354
rect 4734 48190 4786 48242
rect 5742 48190 5794 48242
rect 5966 48190 6018 48242
rect 6302 48190 6354 48242
rect 11118 48190 11170 48242
rect 11790 48190 11842 48242
rect 13358 48190 13410 48242
rect 14814 48190 14866 48242
rect 15934 48190 15986 48242
rect 19966 48190 20018 48242
rect 22430 48190 22482 48242
rect 27246 48190 27298 48242
rect 27470 48190 27522 48242
rect 27918 48190 27970 48242
rect 28254 48190 28306 48242
rect 35982 48190 36034 48242
rect 37102 48190 37154 48242
rect 43262 48190 43314 48242
rect 43486 48190 43538 48242
rect 43934 48190 43986 48242
rect 49198 48190 49250 48242
rect 50094 48190 50146 48242
rect 53678 48190 53730 48242
rect 56142 48190 56194 48242
rect 5182 48078 5234 48130
rect 8990 48078 9042 48130
rect 12462 48078 12514 48130
rect 13694 48078 13746 48130
rect 15150 48078 15202 48130
rect 19630 48078 19682 48130
rect 20974 48078 21026 48130
rect 23774 48078 23826 48130
rect 36654 48078 36706 48130
rect 41582 48078 41634 48130
rect 48862 48078 48914 48130
rect 49646 48078 49698 48130
rect 50878 48078 50930 48130
rect 54238 48078 54290 48130
rect 54910 48078 54962 48130
rect 24334 47966 24386 48018
rect 24670 47966 24722 48018
rect 28366 47966 28418 48018
rect 42478 47966 42530 48018
rect 50206 47966 50258 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 5630 47630 5682 47682
rect 11118 47630 11170 47682
rect 22654 47630 22706 47682
rect 29374 47630 29426 47682
rect 35422 47630 35474 47682
rect 4622 47518 4674 47570
rect 5070 47518 5122 47570
rect 11230 47518 11282 47570
rect 16270 47518 16322 47570
rect 19070 47518 19122 47570
rect 23102 47518 23154 47570
rect 25790 47518 25842 47570
rect 28478 47518 28530 47570
rect 34638 47518 34690 47570
rect 37438 47518 37490 47570
rect 44270 47518 44322 47570
rect 47742 47518 47794 47570
rect 49758 47518 49810 47570
rect 1822 47406 1874 47458
rect 11118 47406 11170 47458
rect 12238 47406 12290 47458
rect 13358 47406 13410 47458
rect 13694 47406 13746 47458
rect 14030 47406 14082 47458
rect 15822 47406 15874 47458
rect 16046 47406 16098 47458
rect 16382 47406 16434 47458
rect 16606 47406 16658 47458
rect 17614 47406 17666 47458
rect 18174 47406 18226 47458
rect 22878 47406 22930 47458
rect 23662 47406 23714 47458
rect 24558 47406 24610 47458
rect 27470 47406 27522 47458
rect 34750 47406 34802 47458
rect 37662 47406 37714 47458
rect 38110 47406 38162 47458
rect 38446 47406 38498 47458
rect 39006 47406 39058 47458
rect 41694 47406 41746 47458
rect 42478 47406 42530 47458
rect 44830 47406 44882 47458
rect 52670 47406 52722 47458
rect 56254 47406 56306 47458
rect 2494 47294 2546 47346
rect 5742 47294 5794 47346
rect 5966 47294 6018 47346
rect 12574 47294 12626 47346
rect 12910 47294 12962 47346
rect 13582 47294 13634 47346
rect 15486 47294 15538 47346
rect 18286 47294 18338 47346
rect 23998 47294 24050 47346
rect 24894 47294 24946 47346
rect 26126 47294 26178 47346
rect 39118 47294 39170 47346
rect 42590 47294 42642 47346
rect 45614 47294 45666 47346
rect 53454 47294 53506 47346
rect 14590 47182 14642 47234
rect 18622 47182 18674 47234
rect 24334 47182 24386 47234
rect 24782 47182 24834 47234
rect 25454 47182 25506 47234
rect 29486 47182 29538 47234
rect 29598 47182 29650 47234
rect 38558 47182 38610 47234
rect 41358 47182 41410 47234
rect 48526 47182 48578 47234
rect 55694 47182 55746 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 2606 46846 2658 46898
rect 24558 46846 24610 46898
rect 27246 46846 27298 46898
rect 32510 46846 32562 46898
rect 35310 46846 35362 46898
rect 36094 46846 36146 46898
rect 36430 46846 36482 46898
rect 45950 46846 46002 46898
rect 53566 46846 53618 46898
rect 2494 46734 2546 46786
rect 5294 46734 5346 46786
rect 8878 46734 8930 46786
rect 12574 46734 12626 46786
rect 12798 46734 12850 46786
rect 23662 46734 23714 46786
rect 28590 46734 28642 46786
rect 28702 46734 28754 46786
rect 29822 46734 29874 46786
rect 31166 46734 31218 46786
rect 34750 46734 34802 46786
rect 35870 46734 35922 46786
rect 37438 46734 37490 46786
rect 39902 46734 39954 46786
rect 41022 46734 41074 46786
rect 41246 46734 41298 46786
rect 46174 46734 46226 46786
rect 48750 46734 48802 46786
rect 4174 46622 4226 46674
rect 8766 46622 8818 46674
rect 9102 46622 9154 46674
rect 11902 46622 11954 46674
rect 13470 46622 13522 46674
rect 13918 46622 13970 46674
rect 14478 46622 14530 46674
rect 14814 46622 14866 46674
rect 17726 46622 17778 46674
rect 19406 46622 19458 46674
rect 23550 46622 23602 46674
rect 24446 46622 24498 46674
rect 26014 46622 26066 46674
rect 27470 46622 27522 46674
rect 28926 46622 28978 46674
rect 32062 46622 32114 46674
rect 34974 46622 35026 46674
rect 35758 46622 35810 46674
rect 36654 46622 36706 46674
rect 38894 46622 38946 46674
rect 44494 46622 44546 46674
rect 44830 46622 44882 46674
rect 45390 46622 45442 46674
rect 45726 46622 45778 46674
rect 47630 46622 47682 46674
rect 48078 46622 48130 46674
rect 49310 46622 49362 46674
rect 49758 46622 49810 46674
rect 50542 46622 50594 46674
rect 53342 46622 53394 46674
rect 53678 46622 53730 46674
rect 54126 46622 54178 46674
rect 55022 46622 55074 46674
rect 2718 46510 2770 46562
rect 3166 46510 3218 46562
rect 3502 46510 3554 46562
rect 5518 46510 5570 46562
rect 10110 46510 10162 46562
rect 12686 46510 12738 46562
rect 15934 46510 15986 46562
rect 17950 46510 18002 46562
rect 26238 46510 26290 46562
rect 26798 46510 26850 46562
rect 29374 46510 29426 46562
rect 31390 46510 31442 46562
rect 31726 46510 31778 46562
rect 37102 46510 37154 46562
rect 41694 46510 41746 46562
rect 45838 46510 45890 46562
rect 50094 46510 50146 46562
rect 51102 46510 51154 46562
rect 53006 46510 53058 46562
rect 54910 46510 54962 46562
rect 19742 46398 19794 46450
rect 32062 46398 32114 46450
rect 36318 46398 36370 46450
rect 40910 46398 40962 46450
rect 41470 46398 41522 46450
rect 41806 46398 41858 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 9662 46062 9714 46114
rect 18174 46062 18226 46114
rect 27358 46062 27410 46114
rect 29262 46062 29314 46114
rect 9102 45950 9154 46002
rect 9998 45950 10050 46002
rect 12126 45950 12178 46002
rect 14030 45950 14082 46002
rect 17950 45950 18002 46002
rect 20190 45950 20242 46002
rect 29710 45950 29762 46002
rect 31054 45950 31106 46002
rect 37550 45950 37602 46002
rect 39566 45950 39618 46002
rect 41694 45950 41746 46002
rect 42142 45950 42194 46002
rect 50654 45950 50706 46002
rect 50878 45950 50930 46002
rect 55246 45950 55298 46002
rect 9326 45838 9378 45890
rect 12798 45838 12850 45890
rect 15038 45838 15090 45890
rect 15822 45838 15874 45890
rect 17054 45838 17106 45890
rect 17838 45838 17890 45890
rect 27246 45838 27298 45890
rect 27918 45838 27970 45890
rect 29038 45838 29090 45890
rect 30158 45838 30210 45890
rect 33966 45838 34018 45890
rect 37998 45838 38050 45890
rect 38894 45838 38946 45890
rect 45054 45838 45106 45890
rect 45278 45838 45330 45890
rect 45502 45838 45554 45890
rect 48414 45838 48466 45890
rect 49310 45838 49362 45890
rect 58046 45838 58098 45890
rect 15486 45726 15538 45778
rect 33182 45726 33234 45778
rect 49534 45726 49586 45778
rect 49982 45726 50034 45778
rect 51214 45726 51266 45778
rect 57374 45726 57426 45778
rect 8094 45614 8146 45666
rect 8206 45614 8258 45666
rect 8318 45614 8370 45666
rect 8542 45614 8594 45666
rect 13582 45614 13634 45666
rect 14814 45614 14866 45666
rect 15598 45614 15650 45666
rect 20750 45614 20802 45666
rect 21422 45614 21474 45666
rect 23102 45614 23154 45666
rect 28590 45614 28642 45666
rect 34414 45614 34466 45666
rect 45390 45614 45442 45666
rect 45950 45614 46002 45666
rect 48078 45614 48130 45666
rect 50990 45614 51042 45666
rect 54910 45614 54962 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 3054 45278 3106 45330
rect 9662 45278 9714 45330
rect 9774 45278 9826 45330
rect 12462 45278 12514 45330
rect 14478 45278 14530 45330
rect 22318 45278 22370 45330
rect 23662 45278 23714 45330
rect 24110 45278 24162 45330
rect 28702 45278 28754 45330
rect 36654 45278 36706 45330
rect 38446 45278 38498 45330
rect 48302 45278 48354 45330
rect 48750 45278 48802 45330
rect 55918 45278 55970 45330
rect 58158 45278 58210 45330
rect 4958 45166 5010 45218
rect 15374 45166 15426 45218
rect 17502 45166 17554 45218
rect 21758 45166 21810 45218
rect 22206 45166 22258 45218
rect 25230 45166 25282 45218
rect 31838 45166 31890 45218
rect 49086 45166 49138 45218
rect 50766 45166 50818 45218
rect 55694 45166 55746 45218
rect 57150 45166 57202 45218
rect 5070 45054 5122 45106
rect 6078 45054 6130 45106
rect 9550 45054 9602 45106
rect 10110 45054 10162 45106
rect 14590 45054 14642 45106
rect 15822 45054 15874 45106
rect 18062 45054 18114 45106
rect 18622 45054 18674 45106
rect 21646 45054 21698 45106
rect 21982 45054 22034 45106
rect 22430 45054 22482 45106
rect 22878 45054 22930 45106
rect 23326 45054 23378 45106
rect 25902 45054 25954 45106
rect 26238 45054 26290 45106
rect 28478 45054 28530 45106
rect 31726 45054 31778 45106
rect 32510 45054 32562 45106
rect 36206 45054 36258 45106
rect 43822 45054 43874 45106
rect 49982 45054 50034 45106
rect 53342 45054 53394 45106
rect 55470 45054 55522 45106
rect 56030 45054 56082 45106
rect 56590 45054 56642 45106
rect 56814 45054 56866 45106
rect 57038 45054 57090 45106
rect 6750 44942 6802 44994
rect 8878 44942 8930 44994
rect 15710 44942 15762 44994
rect 17614 44942 17666 44994
rect 20974 44942 21026 44994
rect 23102 44942 23154 44994
rect 24670 44942 24722 44994
rect 29150 44942 29202 44994
rect 31950 44942 32002 44994
rect 33294 44942 33346 44994
rect 35422 44942 35474 44994
rect 52894 44942 52946 44994
rect 55134 44942 55186 44994
rect 57598 44942 57650 44994
rect 4958 44830 5010 44882
rect 24446 44830 24498 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 3502 44494 3554 44546
rect 5966 44494 6018 44546
rect 31726 44494 31778 44546
rect 45390 44494 45442 44546
rect 51214 44494 51266 44546
rect 54574 44494 54626 44546
rect 55246 44494 55298 44546
rect 56142 44494 56194 44546
rect 57710 44494 57762 44546
rect 58046 44494 58098 44546
rect 4174 44382 4226 44434
rect 5630 44382 5682 44434
rect 7310 44382 7362 44434
rect 8094 44382 8146 44434
rect 8990 44382 9042 44434
rect 9550 44382 9602 44434
rect 16158 44382 16210 44434
rect 19294 44382 19346 44434
rect 35646 44382 35698 44434
rect 43598 44382 43650 44434
rect 45502 44382 45554 44434
rect 51774 44382 51826 44434
rect 54238 44382 54290 44434
rect 58270 44382 58322 44434
rect 2494 44270 2546 44322
rect 4510 44270 4562 44322
rect 4958 44270 5010 44322
rect 6190 44270 6242 44322
rect 7198 44270 7250 44322
rect 7534 44270 7586 44322
rect 8766 44270 8818 44322
rect 13694 44270 13746 44322
rect 15150 44270 15202 44322
rect 18734 44270 18786 44322
rect 21758 44270 21810 44322
rect 22094 44270 22146 44322
rect 23326 44270 23378 44322
rect 24782 44270 24834 44322
rect 31390 44270 31442 44322
rect 32174 44270 32226 44322
rect 32622 44270 32674 44322
rect 33630 44270 33682 44322
rect 34302 44270 34354 44322
rect 34750 44270 34802 44322
rect 40798 44270 40850 44322
rect 44270 44270 44322 44322
rect 44718 44270 44770 44322
rect 45614 44270 45666 44322
rect 46510 44270 46562 44322
rect 46958 44270 47010 44322
rect 51886 44270 51938 44322
rect 55470 44270 55522 44322
rect 56590 44270 56642 44322
rect 56926 44270 56978 44322
rect 2830 44158 2882 44210
rect 3502 44158 3554 44210
rect 3614 44158 3666 44210
rect 3950 44158 4002 44210
rect 7758 44158 7810 44210
rect 13470 44158 13522 44210
rect 15486 44158 15538 44210
rect 17054 44158 17106 44210
rect 22318 44158 22370 44210
rect 22654 44158 22706 44210
rect 24110 44158 24162 44210
rect 24446 44158 24498 44210
rect 25566 44158 25618 44210
rect 25902 44158 25954 44210
rect 31166 44158 31218 44210
rect 33070 44158 33122 44210
rect 34078 44158 34130 44210
rect 35086 44158 35138 44210
rect 41470 44158 41522 44210
rect 43934 44158 43986 44210
rect 44046 44158 44098 44210
rect 46846 44158 46898 44210
rect 56702 44158 56754 44210
rect 57598 44158 57650 44210
rect 2718 44046 2770 44098
rect 15374 44046 15426 44098
rect 22766 44046 22818 44098
rect 22878 44046 22930 44098
rect 23662 44046 23714 44098
rect 33966 44046 34018 44098
rect 34638 44046 34690 44098
rect 34862 44046 34914 44098
rect 37886 44046 37938 44098
rect 46622 44046 46674 44098
rect 54350 44046 54402 44098
rect 54910 44046 54962 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 4958 43710 5010 43762
rect 14702 43710 14754 43762
rect 23214 43710 23266 43762
rect 32398 43710 32450 43762
rect 37662 43710 37714 43762
rect 2494 43598 2546 43650
rect 5070 43598 5122 43650
rect 5518 43598 5570 43650
rect 13918 43598 13970 43650
rect 16382 43598 16434 43650
rect 17726 43598 17778 43650
rect 18398 43598 18450 43650
rect 22206 43598 22258 43650
rect 22766 43598 22818 43650
rect 29822 43598 29874 43650
rect 36654 43598 36706 43650
rect 38558 43598 38610 43650
rect 46062 43598 46114 43650
rect 57374 43598 57426 43650
rect 57822 43598 57874 43650
rect 1822 43486 1874 43538
rect 13806 43486 13858 43538
rect 14814 43486 14866 43538
rect 15486 43486 15538 43538
rect 17502 43486 17554 43538
rect 19070 43486 19122 43538
rect 22542 43486 22594 43538
rect 29710 43486 29762 43538
rect 29934 43486 29986 43538
rect 30270 43486 30322 43538
rect 31838 43486 31890 43538
rect 32062 43486 32114 43538
rect 37102 43486 37154 43538
rect 37774 43486 37826 43538
rect 39678 43486 39730 43538
rect 41022 43486 41074 43538
rect 41470 43486 41522 43538
rect 45278 43486 45330 43538
rect 52782 43486 52834 43538
rect 53230 43486 53282 43538
rect 4622 43374 4674 43426
rect 16158 43374 16210 43426
rect 17390 43374 17442 43426
rect 19742 43374 19794 43426
rect 21870 43374 21922 43426
rect 22318 43374 22370 43426
rect 38222 43374 38274 43426
rect 40350 43374 40402 43426
rect 42478 43374 42530 43426
rect 44942 43374 44994 43426
rect 48190 43374 48242 43426
rect 54798 43374 54850 43426
rect 57150 43374 57202 43426
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 10110 42926 10162 42978
rect 15934 42926 15986 42978
rect 20190 42926 20242 42978
rect 30942 42926 30994 42978
rect 37102 42926 37154 42978
rect 41358 42926 41410 42978
rect 45614 42926 45666 42978
rect 50094 42926 50146 42978
rect 53566 42926 53618 42978
rect 53678 42926 53730 42978
rect 2942 42814 2994 42866
rect 3726 42814 3778 42866
rect 8430 42814 8482 42866
rect 16382 42814 16434 42866
rect 22094 42814 22146 42866
rect 25342 42814 25394 42866
rect 31278 42814 31330 42866
rect 33518 42814 33570 42866
rect 36430 42814 36482 42866
rect 40238 42814 40290 42866
rect 44158 42814 44210 42866
rect 46734 42814 46786 42866
rect 51662 42814 51714 42866
rect 57038 42814 57090 42866
rect 3614 42702 3666 42754
rect 8878 42702 8930 42754
rect 9662 42702 9714 42754
rect 10110 42702 10162 42754
rect 10558 42702 10610 42754
rect 12574 42702 12626 42754
rect 16494 42702 16546 42754
rect 18174 42702 18226 42754
rect 19630 42702 19682 42754
rect 24782 42702 24834 42754
rect 26014 42702 26066 42754
rect 26238 42702 26290 42754
rect 27134 42702 27186 42754
rect 27470 42702 27522 42754
rect 27694 42702 27746 42754
rect 28366 42702 28418 42754
rect 29150 42702 29202 42754
rect 30046 42702 30098 42754
rect 30942 42702 30994 42754
rect 37774 42702 37826 42754
rect 38110 42702 38162 42754
rect 39342 42702 39394 42754
rect 39790 42702 39842 42754
rect 40798 42702 40850 42754
rect 46622 42702 46674 42754
rect 51550 42702 51602 42754
rect 51774 42702 51826 42754
rect 53902 42702 53954 42754
rect 55918 42702 55970 42754
rect 56478 42702 56530 42754
rect 8766 42590 8818 42642
rect 14142 42590 14194 42642
rect 15598 42590 15650 42642
rect 16830 42590 16882 42642
rect 20302 42590 20354 42642
rect 20750 42590 20802 42642
rect 21310 42590 21362 42642
rect 21646 42590 21698 42642
rect 25006 42590 25058 42642
rect 30606 42590 30658 42642
rect 37214 42590 37266 42642
rect 38558 42590 38610 42642
rect 40574 42590 40626 42642
rect 41694 42590 41746 42642
rect 42030 42590 42082 42642
rect 42254 42590 42306 42642
rect 43934 42590 43986 42642
rect 45614 42590 45666 42642
rect 45726 42590 45778 42642
rect 50206 42590 50258 42642
rect 54014 42590 54066 42642
rect 55470 42590 55522 42642
rect 56926 42590 56978 42642
rect 8990 42478 9042 42530
rect 12350 42478 12402 42530
rect 13806 42478 13858 42530
rect 15822 42478 15874 42530
rect 20526 42478 20578 42530
rect 28478 42478 28530 42530
rect 28702 42478 28754 42530
rect 29262 42478 29314 42530
rect 29486 42478 29538 42530
rect 33182 42478 33234 42530
rect 34078 42478 34130 42530
rect 37102 42478 37154 42530
rect 37662 42478 37714 42530
rect 41470 42478 41522 42530
rect 45166 42478 45218 42530
rect 46398 42478 46450 42530
rect 46846 42478 46898 42530
rect 49646 42478 49698 42530
rect 50094 42478 50146 42530
rect 51998 42478 52050 42530
rect 53118 42478 53170 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 9662 42142 9714 42194
rect 28030 42142 28082 42194
rect 28478 42142 28530 42194
rect 32622 42142 32674 42194
rect 33630 42142 33682 42194
rect 11566 42030 11618 42082
rect 13582 42030 13634 42082
rect 15038 42030 15090 42082
rect 15598 42030 15650 42082
rect 19518 42030 19570 42082
rect 21198 42030 21250 42082
rect 21646 42030 21698 42082
rect 23662 42030 23714 42082
rect 23774 42030 23826 42082
rect 27246 42030 27298 42082
rect 34078 42030 34130 42082
rect 35534 42030 35586 42082
rect 53790 42030 53842 42082
rect 57038 42030 57090 42082
rect 5406 41918 5458 41970
rect 8990 41918 9042 41970
rect 9550 41918 9602 41970
rect 9886 41918 9938 41970
rect 11678 41918 11730 41970
rect 12798 41918 12850 41970
rect 14702 41918 14754 41970
rect 15374 41918 15426 41970
rect 16046 41918 16098 41970
rect 16718 41918 16770 41970
rect 18286 41918 18338 41970
rect 18734 41918 18786 41970
rect 20414 41918 20466 41970
rect 20750 41918 20802 41970
rect 21534 41918 21586 41970
rect 25118 41918 25170 41970
rect 25902 41918 25954 41970
rect 26910 41918 26962 41970
rect 27918 41918 27970 41970
rect 28142 41918 28194 41970
rect 28590 41918 28642 41970
rect 28702 41918 28754 41970
rect 29038 41918 29090 41970
rect 29486 41918 29538 41970
rect 29710 41918 29762 41970
rect 30382 41918 30434 41970
rect 35870 41918 35922 41970
rect 36878 41918 36930 41970
rect 38782 41918 38834 41970
rect 41134 41918 41186 41970
rect 41358 41918 41410 41970
rect 41694 41918 41746 41970
rect 43822 41918 43874 41970
rect 49198 41918 49250 41970
rect 52446 41918 52498 41970
rect 53118 41918 53170 41970
rect 57374 41918 57426 41970
rect 57710 41918 57762 41970
rect 58158 41918 58210 41970
rect 3278 41806 3330 41858
rect 6078 41806 6130 41858
rect 8206 41806 8258 41858
rect 8766 41806 8818 41858
rect 10334 41806 10386 41858
rect 14590 41806 14642 41858
rect 19966 41806 20018 41858
rect 22542 41806 22594 41858
rect 22878 41806 22930 41858
rect 25790 41806 25842 41858
rect 33742 41806 33794 41858
rect 34414 41806 34466 41858
rect 37214 41806 37266 41858
rect 38110 41806 38162 41858
rect 38894 41806 38946 41858
rect 40350 41806 40402 41858
rect 41246 41806 41298 41858
rect 42142 41806 42194 41858
rect 43486 41806 43538 41858
rect 44494 41806 44546 41858
rect 49870 41806 49922 41858
rect 51998 41806 52050 41858
rect 55918 41806 55970 41858
rect 56702 41806 56754 41858
rect 57486 41806 57538 41858
rect 8654 41694 8706 41746
rect 15262 41694 15314 41746
rect 22542 41694 22594 41746
rect 22878 41694 22930 41746
rect 23662 41694 23714 41746
rect 25678 41694 25730 41746
rect 27694 41694 27746 41746
rect 33406 41694 33458 41746
rect 34638 41694 34690 41746
rect 39006 41694 39058 41746
rect 43822 41694 43874 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 27134 41358 27186 41410
rect 32286 41358 32338 41410
rect 44158 41358 44210 41410
rect 45166 41358 45218 41410
rect 50318 41358 50370 41410
rect 52894 41358 52946 41410
rect 2718 41246 2770 41298
rect 4174 41246 4226 41298
rect 21310 41246 21362 41298
rect 22318 41246 22370 41298
rect 23326 41246 23378 41298
rect 23774 41246 23826 41298
rect 24894 41246 24946 41298
rect 27470 41246 27522 41298
rect 32510 41246 32562 41298
rect 33630 41246 33682 41298
rect 34862 41246 34914 41298
rect 36990 41246 37042 41298
rect 38558 41246 38610 41298
rect 40126 41246 40178 41298
rect 43486 41246 43538 41298
rect 45502 41246 45554 41298
rect 50542 41246 50594 41298
rect 52670 41246 52722 41298
rect 4062 41134 4114 41186
rect 5182 41134 5234 41186
rect 5518 41134 5570 41186
rect 8542 41134 8594 41186
rect 9550 41134 9602 41186
rect 15150 41134 15202 41186
rect 15710 41134 15762 41186
rect 17838 41134 17890 41186
rect 19518 41134 19570 41186
rect 20526 41134 20578 41186
rect 21870 41134 21922 41186
rect 23438 41134 23490 41186
rect 25118 41134 25170 41186
rect 25566 41134 25618 41186
rect 25902 41134 25954 41186
rect 28030 41134 28082 41186
rect 29038 41134 29090 41186
rect 32062 41134 32114 41186
rect 33182 41134 33234 41186
rect 33966 41134 34018 41186
rect 34638 41134 34690 41186
rect 34750 41134 34802 41186
rect 35534 41134 35586 41186
rect 35758 41134 35810 41186
rect 36094 41134 36146 41186
rect 37102 41134 37154 41186
rect 37438 41134 37490 41186
rect 43038 41134 43090 41186
rect 51886 41134 51938 41186
rect 51998 41134 52050 41186
rect 53118 41134 53170 41186
rect 55694 41134 55746 41186
rect 57598 41134 57650 41186
rect 2830 41022 2882 41074
rect 3054 41022 3106 41074
rect 3726 41022 3778 41074
rect 5854 41022 5906 41074
rect 9662 41022 9714 41074
rect 12686 41022 12738 41074
rect 16382 41022 16434 41074
rect 17166 41022 17218 41074
rect 18734 41022 18786 41074
rect 19966 41022 20018 41074
rect 20190 41022 20242 41074
rect 26462 41022 26514 41074
rect 26574 41022 26626 41074
rect 26686 41022 26738 41074
rect 29374 41022 29426 41074
rect 42254 41022 42306 41074
rect 44270 41022 44322 41074
rect 51550 41022 51602 41074
rect 55358 41022 55410 41074
rect 57262 41022 57314 41074
rect 5742 40910 5794 40962
rect 8318 40910 8370 40962
rect 12350 40910 12402 40962
rect 14590 40910 14642 40962
rect 20302 40910 20354 40962
rect 27470 40910 27522 40962
rect 27694 40910 27746 40962
rect 29262 40910 29314 40962
rect 34078 40910 34130 40962
rect 34974 40910 35026 40962
rect 35086 40910 35138 40962
rect 44158 40910 44210 40962
rect 45390 40910 45442 40962
rect 50542 40910 50594 40962
rect 51662 40910 51714 40962
rect 53566 40910 53618 40962
rect 56030 40910 56082 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 5070 40574 5122 40626
rect 8094 40574 8146 40626
rect 12238 40574 12290 40626
rect 13582 40574 13634 40626
rect 14590 40574 14642 40626
rect 19742 40574 19794 40626
rect 22542 40574 22594 40626
rect 24334 40574 24386 40626
rect 41134 40574 41186 40626
rect 55694 40574 55746 40626
rect 58158 40574 58210 40626
rect 2494 40462 2546 40514
rect 6190 40462 6242 40514
rect 6526 40462 6578 40514
rect 12462 40462 12514 40514
rect 13358 40462 13410 40514
rect 14366 40462 14418 40514
rect 16718 40462 16770 40514
rect 17950 40462 18002 40514
rect 21198 40462 21250 40514
rect 21310 40462 21362 40514
rect 24110 40462 24162 40514
rect 34862 40462 34914 40514
rect 35646 40462 35698 40514
rect 38782 40462 38834 40514
rect 40238 40462 40290 40514
rect 40350 40462 40402 40514
rect 43486 40462 43538 40514
rect 45950 40462 46002 40514
rect 55918 40462 55970 40514
rect 56702 40462 56754 40514
rect 1822 40350 1874 40402
rect 7870 40350 7922 40402
rect 12574 40350 12626 40402
rect 13806 40350 13858 40402
rect 14254 40350 14306 40402
rect 14814 40350 14866 40402
rect 15150 40350 15202 40402
rect 15710 40350 15762 40402
rect 17502 40350 17554 40402
rect 20302 40350 20354 40402
rect 20862 40350 20914 40402
rect 21870 40350 21922 40402
rect 22990 40350 23042 40402
rect 23774 40350 23826 40402
rect 27134 40350 27186 40402
rect 27806 40350 27858 40402
rect 28926 40350 28978 40402
rect 29262 40350 29314 40402
rect 31390 40350 31442 40402
rect 34526 40350 34578 40402
rect 35758 40350 35810 40402
rect 37998 40350 38050 40402
rect 40798 40350 40850 40402
rect 41246 40350 41298 40402
rect 41358 40350 41410 40402
rect 43822 40350 43874 40402
rect 44718 40350 44770 40402
rect 45166 40350 45218 40402
rect 48750 40350 48802 40402
rect 49310 40350 49362 40402
rect 51662 40350 51714 40402
rect 56030 40350 56082 40402
rect 57038 40350 57090 40402
rect 57486 40350 57538 40402
rect 4622 40238 4674 40290
rect 8542 40238 8594 40290
rect 13694 40238 13746 40290
rect 15374 40238 15426 40290
rect 19182 40238 19234 40290
rect 22654 40238 22706 40290
rect 23438 40238 23490 40290
rect 24446 40238 24498 40290
rect 27582 40238 27634 40290
rect 28030 40238 28082 40290
rect 29374 40238 29426 40290
rect 31166 40238 31218 40290
rect 35870 40238 35922 40290
rect 38110 40238 38162 40290
rect 43710 40238 43762 40290
rect 48078 40238 48130 40290
rect 50990 40238 51042 40290
rect 51774 40238 51826 40290
rect 56926 40238 56978 40290
rect 16606 40126 16658 40178
rect 21310 40126 21362 40178
rect 22318 40126 22370 40178
rect 40238 40126 40290 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 5630 39790 5682 39842
rect 5966 39790 6018 39842
rect 26014 39790 26066 39842
rect 45838 39790 45890 39842
rect 47406 39790 47458 39842
rect 51326 39790 51378 39842
rect 57486 39790 57538 39842
rect 57822 39790 57874 39842
rect 4622 39678 4674 39730
rect 6862 39678 6914 39730
rect 12798 39678 12850 39730
rect 14590 39678 14642 39730
rect 14814 39678 14866 39730
rect 17726 39678 17778 39730
rect 17838 39678 17890 39730
rect 22654 39678 22706 39730
rect 23774 39678 23826 39730
rect 26126 39678 26178 39730
rect 27918 39678 27970 39730
rect 32174 39678 32226 39730
rect 32510 39678 32562 39730
rect 35198 39678 35250 39730
rect 45278 39678 45330 39730
rect 47518 39678 47570 39730
rect 50654 39678 50706 39730
rect 50990 39678 51042 39730
rect 56478 39678 56530 39730
rect 3166 39566 3218 39618
rect 11454 39566 11506 39618
rect 12350 39566 12402 39618
rect 14142 39566 14194 39618
rect 14926 39566 14978 39618
rect 15934 39566 15986 39618
rect 18734 39566 18786 39618
rect 20190 39566 20242 39618
rect 22206 39566 22258 39618
rect 25566 39566 25618 39618
rect 26238 39566 26290 39618
rect 26462 39566 26514 39618
rect 31278 39566 31330 39618
rect 31502 39566 31554 39618
rect 34638 39566 34690 39618
rect 34862 39566 34914 39618
rect 41694 39566 41746 39618
rect 43374 39566 43426 39618
rect 43822 39566 43874 39618
rect 45390 39566 45442 39618
rect 49198 39566 49250 39618
rect 53678 39566 53730 39618
rect 57038 39566 57090 39618
rect 4286 39454 4338 39506
rect 5742 39454 5794 39506
rect 12798 39454 12850 39506
rect 13806 39454 13858 39506
rect 16494 39454 16546 39506
rect 20414 39454 20466 39506
rect 21310 39454 21362 39506
rect 21646 39454 21698 39506
rect 25006 39454 25058 39506
rect 44270 39454 44322 39506
rect 45054 39454 45106 39506
rect 45726 39454 45778 39506
rect 51102 39454 51154 39506
rect 54350 39454 54402 39506
rect 56814 39454 56866 39506
rect 57598 39454 57650 39506
rect 2830 39342 2882 39394
rect 11566 39342 11618 39394
rect 13470 39342 13522 39394
rect 23998 39342 24050 39394
rect 27470 39342 27522 39394
rect 33070 39342 33122 39394
rect 42254 39342 42306 39394
rect 45838 39342 45890 39394
rect 48974 39342 49026 39394
rect 49758 39342 49810 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 6190 39006 6242 39058
rect 8206 39006 8258 39058
rect 8542 39006 8594 39058
rect 13134 39006 13186 39058
rect 18846 39006 18898 39058
rect 19630 39006 19682 39058
rect 27694 39006 27746 39058
rect 27918 39006 27970 39058
rect 44830 39006 44882 39058
rect 48862 39006 48914 39058
rect 53566 39006 53618 39058
rect 54126 39006 54178 39058
rect 7982 38894 8034 38946
rect 12126 38894 12178 38946
rect 12350 38894 12402 38946
rect 17838 38894 17890 38946
rect 20526 38894 20578 38946
rect 30382 38894 30434 38946
rect 37550 38894 37602 38946
rect 37886 38894 37938 38946
rect 39454 38894 39506 38946
rect 50990 38894 51042 38946
rect 57822 38894 57874 38946
rect 6414 38782 6466 38834
rect 6638 38782 6690 38834
rect 7086 38782 7138 38834
rect 7870 38782 7922 38834
rect 11342 38782 11394 38834
rect 12462 38782 12514 38834
rect 12686 38782 12738 38834
rect 15710 38782 15762 38834
rect 16046 38782 16098 38834
rect 20974 38782 21026 38834
rect 21310 38782 21362 38834
rect 23438 38782 23490 38834
rect 23662 38782 23714 38834
rect 24110 38782 24162 38834
rect 25678 38782 25730 38834
rect 27022 38782 27074 38834
rect 27246 38782 27298 38834
rect 28030 38782 28082 38834
rect 30046 38782 30098 38834
rect 30606 38782 30658 38834
rect 32510 38782 32562 38834
rect 34078 38782 34130 38834
rect 34750 38782 34802 38834
rect 39678 38782 39730 38834
rect 40014 38782 40066 38834
rect 50318 38782 50370 38834
rect 58158 38782 58210 38834
rect 6526 38670 6578 38722
rect 7422 38670 7474 38722
rect 11566 38670 11618 38722
rect 15822 38670 15874 38722
rect 22654 38670 22706 38722
rect 23886 38670 23938 38722
rect 25566 38670 25618 38722
rect 26910 38670 26962 38722
rect 29934 38670 29986 38722
rect 32174 38670 32226 38722
rect 34302 38670 34354 38722
rect 34974 38670 35026 38722
rect 39230 38670 39282 38722
rect 45950 38670 46002 38722
rect 46174 38670 46226 38722
rect 49422 38670 49474 38722
rect 53118 38670 53170 38722
rect 53902 38670 53954 38722
rect 54238 38670 54290 38722
rect 56702 38670 56754 38722
rect 57598 38670 57650 38722
rect 11006 38558 11058 38610
rect 15374 38558 15426 38610
rect 24222 38558 24274 38610
rect 26574 38558 26626 38610
rect 30270 38558 30322 38610
rect 30830 38558 30882 38610
rect 31950 38558 32002 38610
rect 46510 38558 46562 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 3950 38222 4002 38274
rect 9774 38222 9826 38274
rect 11790 38222 11842 38274
rect 12238 38222 12290 38274
rect 12574 38222 12626 38274
rect 13694 38222 13746 38274
rect 24558 38222 24610 38274
rect 26014 38222 26066 38274
rect 29262 38222 29314 38274
rect 30494 38222 30546 38274
rect 4510 38110 4562 38162
rect 6862 38110 6914 38162
rect 7758 38110 7810 38162
rect 12798 38110 12850 38162
rect 16606 38110 16658 38162
rect 17950 38110 18002 38162
rect 19742 38110 19794 38162
rect 21198 38110 21250 38162
rect 27022 38110 27074 38162
rect 27582 38110 27634 38162
rect 28142 38110 28194 38162
rect 36318 38110 36370 38162
rect 58158 38166 58210 38218
rect 38334 38110 38386 38162
rect 38782 38110 38834 38162
rect 46398 38110 46450 38162
rect 4062 37998 4114 38050
rect 5854 37998 5906 38050
rect 6190 37998 6242 38050
rect 6414 37998 6466 38050
rect 7198 37998 7250 38050
rect 8766 37998 8818 38050
rect 9438 37998 9490 38050
rect 11454 37998 11506 38050
rect 14030 37998 14082 38050
rect 14814 37998 14866 38050
rect 17054 37998 17106 38050
rect 17614 37998 17666 38050
rect 20190 37998 20242 38050
rect 21310 37998 21362 38050
rect 22990 37998 23042 38050
rect 24222 37998 24274 38050
rect 26126 37998 26178 38050
rect 27134 37998 27186 38050
rect 27470 37998 27522 38050
rect 28590 37998 28642 38050
rect 31278 37998 31330 38050
rect 32958 37998 33010 38050
rect 34414 37998 34466 38050
rect 35310 37998 35362 38050
rect 36542 37998 36594 38050
rect 37102 37998 37154 38050
rect 40238 37998 40290 38050
rect 41582 37998 41634 38050
rect 42142 37998 42194 38050
rect 45390 37998 45442 38050
rect 45838 37998 45890 38050
rect 49310 37998 49362 38050
rect 54910 37998 54962 38050
rect 55358 37998 55410 38050
rect 8654 37886 8706 37938
rect 10670 37886 10722 37938
rect 11230 37886 11282 37938
rect 14702 37886 14754 37938
rect 21534 37886 21586 37938
rect 22094 37886 22146 37938
rect 22766 37886 22818 37938
rect 23998 37886 24050 37938
rect 28142 37886 28194 37938
rect 29262 37886 29314 37938
rect 29374 37886 29426 37938
rect 30606 37886 30658 37938
rect 31838 37886 31890 37938
rect 35086 37886 35138 37938
rect 35646 37886 35698 37938
rect 35982 37886 36034 37938
rect 37326 37886 37378 37938
rect 37662 37886 37714 37938
rect 39006 37886 39058 37938
rect 46062 37886 46114 37938
rect 48526 37886 48578 37938
rect 56030 37886 56082 37938
rect 3950 37774 4002 37826
rect 5966 37774 6018 37826
rect 16158 37774 16210 37826
rect 26014 37774 26066 37826
rect 28366 37774 28418 37826
rect 30494 37774 30546 37826
rect 34862 37774 34914 37826
rect 35534 37774 35586 37826
rect 36206 37774 36258 37826
rect 40798 37774 40850 37826
rect 45278 37774 45330 37826
rect 45950 37774 46002 37826
rect 49758 37774 49810 37826
rect 53566 37774 53618 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 3614 37438 3666 37490
rect 7870 37438 7922 37490
rect 8990 37438 9042 37490
rect 12574 37438 12626 37490
rect 14142 37438 14194 37490
rect 17502 37438 17554 37490
rect 24558 37438 24610 37490
rect 25342 37438 25394 37490
rect 30718 37438 30770 37490
rect 37102 37438 37154 37490
rect 39006 37438 39058 37490
rect 39902 37438 39954 37490
rect 44270 37438 44322 37490
rect 46510 37438 46562 37490
rect 46622 37438 46674 37490
rect 2718 37326 2770 37378
rect 3054 37326 3106 37378
rect 5294 37326 5346 37378
rect 8430 37326 8482 37378
rect 8654 37326 8706 37378
rect 8766 37326 8818 37378
rect 11342 37326 11394 37378
rect 12238 37326 12290 37378
rect 12462 37326 12514 37378
rect 14366 37326 14418 37378
rect 14478 37326 14530 37378
rect 14814 37326 14866 37378
rect 16830 37326 16882 37378
rect 23662 37326 23714 37378
rect 26014 37326 26066 37378
rect 26126 37326 26178 37378
rect 26798 37326 26850 37378
rect 35758 37326 35810 37378
rect 37214 37326 37266 37378
rect 37774 37326 37826 37378
rect 39566 37326 39618 37378
rect 39678 37326 39730 37378
rect 46398 37326 46450 37378
rect 3166 37214 3218 37266
rect 3726 37214 3778 37266
rect 3838 37214 3890 37266
rect 4286 37214 4338 37266
rect 4622 37214 4674 37266
rect 9438 37214 9490 37266
rect 10222 37214 10274 37266
rect 11902 37214 11954 37266
rect 14926 37214 14978 37266
rect 15374 37214 15426 37266
rect 15934 37214 15986 37266
rect 16494 37214 16546 37266
rect 18846 37214 18898 37266
rect 20302 37214 20354 37266
rect 21422 37214 21474 37266
rect 24558 37214 24610 37266
rect 26574 37214 26626 37266
rect 27134 37214 27186 37266
rect 27582 37214 27634 37266
rect 29150 37214 29202 37266
rect 31278 37214 31330 37266
rect 33406 37214 33458 37266
rect 33630 37214 33682 37266
rect 36654 37214 36706 37266
rect 37102 37214 37154 37266
rect 39230 37214 39282 37266
rect 43822 37214 43874 37266
rect 2830 37102 2882 37154
rect 7422 37102 7474 37154
rect 8878 37102 8930 37154
rect 16718 37102 16770 37154
rect 20414 37102 20466 37154
rect 21198 37102 21250 37154
rect 22878 37102 22930 37154
rect 25230 37102 25282 37154
rect 34078 37102 34130 37154
rect 40910 37102 40962 37154
rect 43038 37102 43090 37154
rect 9662 36990 9714 37042
rect 11118 36990 11170 37042
rect 15150 36990 15202 37042
rect 20638 36990 20690 37042
rect 27246 36990 27298 37042
rect 31054 36990 31106 37042
rect 38894 36990 38946 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 23102 36654 23154 36706
rect 24558 36654 24610 36706
rect 27358 36654 27410 36706
rect 35646 36654 35698 36706
rect 36878 36654 36930 36706
rect 40910 36654 40962 36706
rect 41246 36654 41298 36706
rect 2494 36542 2546 36594
rect 4622 36542 4674 36594
rect 5182 36542 5234 36594
rect 9326 36542 9378 36594
rect 11902 36542 11954 36594
rect 15822 36542 15874 36594
rect 16270 36542 16322 36594
rect 17278 36542 17330 36594
rect 22542 36542 22594 36594
rect 24110 36542 24162 36594
rect 27022 36542 27074 36594
rect 28366 36542 28418 36594
rect 30718 36542 30770 36594
rect 33294 36542 33346 36594
rect 35534 36542 35586 36594
rect 37886 36542 37938 36594
rect 52110 36542 52162 36594
rect 52894 36542 52946 36594
rect 56142 36542 56194 36594
rect 56702 36542 56754 36594
rect 1822 36430 1874 36482
rect 8542 36430 8594 36482
rect 11454 36430 11506 36482
rect 12798 36430 12850 36482
rect 13470 36430 13522 36482
rect 15710 36430 15762 36482
rect 16830 36430 16882 36482
rect 17726 36430 17778 36482
rect 18286 36430 18338 36482
rect 18846 36430 18898 36482
rect 19406 36430 19458 36482
rect 22766 36430 22818 36482
rect 23662 36430 23714 36482
rect 23998 36430 24050 36482
rect 24334 36430 24386 36482
rect 24670 36430 24722 36482
rect 26910 36430 26962 36482
rect 33070 36430 33122 36482
rect 35422 36430 35474 36482
rect 36206 36430 36258 36482
rect 37102 36430 37154 36482
rect 37662 36430 37714 36482
rect 49310 36430 49362 36482
rect 53342 36430 53394 36482
rect 8878 36318 8930 36370
rect 11118 36318 11170 36370
rect 11566 36318 11618 36370
rect 17614 36318 17666 36370
rect 19630 36318 19682 36370
rect 32062 36318 32114 36370
rect 37438 36318 37490 36370
rect 44046 36318 44098 36370
rect 49982 36318 50034 36370
rect 54014 36318 54066 36370
rect 8766 36206 8818 36258
rect 9774 36206 9826 36258
rect 10782 36206 10834 36258
rect 11006 36206 11058 36258
rect 12686 36206 12738 36258
rect 13582 36206 13634 36258
rect 13806 36206 13858 36258
rect 20750 36206 20802 36258
rect 21310 36206 21362 36258
rect 21646 36206 21698 36258
rect 27806 36206 27858 36258
rect 31166 36206 31218 36258
rect 32958 36206 33010 36258
rect 41134 36206 41186 36258
rect 41694 36206 41746 36258
rect 43822 36206 43874 36258
rect 43934 36206 43986 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 11678 35870 11730 35922
rect 12910 35870 12962 35922
rect 23326 35870 23378 35922
rect 24222 35870 24274 35922
rect 27246 35870 27298 35922
rect 28366 35870 28418 35922
rect 31390 35870 31442 35922
rect 37326 35870 37378 35922
rect 38334 35870 38386 35922
rect 38782 35870 38834 35922
rect 39006 35870 39058 35922
rect 50430 35870 50482 35922
rect 2270 35758 2322 35810
rect 10334 35758 10386 35810
rect 12798 35758 12850 35810
rect 15038 35758 15090 35810
rect 18846 35758 18898 35810
rect 27358 35758 27410 35810
rect 30942 35758 30994 35810
rect 32398 35758 32450 35810
rect 34974 35758 35026 35810
rect 36318 35758 36370 35810
rect 50990 35870 51042 35922
rect 51214 35870 51266 35922
rect 55134 35870 55186 35922
rect 56814 35870 56866 35922
rect 57710 35870 57762 35922
rect 37438 35758 37490 35810
rect 44830 35758 44882 35810
rect 50766 35758 50818 35810
rect 1822 35646 1874 35698
rect 10110 35646 10162 35698
rect 11342 35646 11394 35698
rect 11678 35646 11730 35698
rect 12014 35646 12066 35698
rect 12350 35646 12402 35698
rect 12574 35646 12626 35698
rect 13918 35646 13970 35698
rect 15822 35646 15874 35698
rect 18510 35646 18562 35698
rect 20302 35646 20354 35698
rect 21086 35646 21138 35698
rect 23998 35646 24050 35698
rect 25342 35646 25394 35698
rect 30494 35646 30546 35698
rect 31390 35646 31442 35698
rect 32510 35646 32562 35698
rect 35982 35646 36034 35698
rect 36430 35646 36482 35698
rect 36654 35646 36706 35698
rect 37662 35646 37714 35698
rect 37998 35646 38050 35698
rect 39118 35646 39170 35698
rect 42478 35646 42530 35698
rect 45502 35646 45554 35698
rect 50654 35646 50706 35698
rect 52110 35646 52162 35698
rect 52894 35646 52946 35698
rect 54910 35646 54962 35698
rect 55358 35646 55410 35698
rect 55582 35646 55634 35698
rect 56590 35646 56642 35698
rect 57038 35646 57090 35698
rect 57150 35646 57202 35698
rect 57598 35646 57650 35698
rect 57934 35646 57986 35698
rect 13582 35534 13634 35586
rect 16046 35534 16098 35586
rect 18622 35534 18674 35586
rect 22878 35534 22930 35586
rect 25678 35534 25730 35586
rect 33630 35534 33682 35586
rect 34190 35534 34242 35586
rect 38222 35534 38274 35586
rect 42702 35534 42754 35586
rect 51998 35534 52050 35586
rect 21646 35422 21698 35474
rect 32398 35422 32450 35474
rect 50318 35422 50370 35474
rect 51774 35422 51826 35474
rect 53118 35422 53170 35474
rect 53454 35422 53506 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 10670 35086 10722 35138
rect 37550 35086 37602 35138
rect 38110 35086 38162 35138
rect 44942 35086 44994 35138
rect 1822 34974 1874 35026
rect 10334 34974 10386 35026
rect 17054 34974 17106 35026
rect 20078 34974 20130 35026
rect 24222 34974 24274 35026
rect 28366 34974 28418 35026
rect 29710 34974 29762 35026
rect 35758 34974 35810 35026
rect 37886 34974 37938 35026
rect 40798 34974 40850 35026
rect 44046 34974 44098 35026
rect 45502 34974 45554 35026
rect 46062 34974 46114 35026
rect 49982 34974 50034 35026
rect 7310 34862 7362 34914
rect 7982 34862 8034 34914
rect 9886 34862 9938 34914
rect 10558 34862 10610 34914
rect 12798 34862 12850 34914
rect 15374 34862 15426 34914
rect 21310 34862 21362 34914
rect 27918 34862 27970 34914
rect 30270 34862 30322 34914
rect 36206 34862 36258 34914
rect 43934 34862 43986 34914
rect 48862 34862 48914 34914
rect 53230 34862 53282 34914
rect 55470 34862 55522 34914
rect 56590 34862 56642 34914
rect 7534 34750 7586 34802
rect 12574 34750 12626 34802
rect 16270 34750 16322 34802
rect 20862 34750 20914 34802
rect 22094 34750 22146 34802
rect 29822 34750 29874 34802
rect 34974 34750 35026 34802
rect 36990 34750 37042 34802
rect 43598 34750 43650 34802
rect 44158 34750 44210 34802
rect 44942 34750 44994 34802
rect 45054 34750 45106 34802
rect 48190 34750 48242 34802
rect 49422 34750 49474 34802
rect 49534 34750 49586 34802
rect 55806 34750 55858 34802
rect 56254 34750 56306 34802
rect 56366 34750 56418 34802
rect 56926 34750 56978 34802
rect 57038 34750 57090 34802
rect 8094 34638 8146 34690
rect 16718 34638 16770 34690
rect 19518 34638 19570 34690
rect 27582 34638 27634 34690
rect 29374 34638 29426 34690
rect 29598 34638 29650 34690
rect 37214 34638 37266 34690
rect 37438 34638 37490 34690
rect 37886 34638 37938 34690
rect 38670 34638 38722 34690
rect 39342 34638 39394 34690
rect 53454 34638 53506 34690
rect 55694 34638 55746 34690
rect 56702 34638 56754 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 7870 34302 7922 34354
rect 8094 34302 8146 34354
rect 9662 34302 9714 34354
rect 15150 34302 15202 34354
rect 19294 34302 19346 34354
rect 20302 34302 20354 34354
rect 29150 34302 29202 34354
rect 29822 34302 29874 34354
rect 34078 34302 34130 34354
rect 41246 34302 41298 34354
rect 41470 34302 41522 34354
rect 42366 34302 42418 34354
rect 44270 34302 44322 34354
rect 44494 34302 44546 34354
rect 54686 34302 54738 34354
rect 8430 34190 8482 34242
rect 10446 34190 10498 34242
rect 10782 34190 10834 34242
rect 17950 34190 18002 34242
rect 30270 34190 30322 34242
rect 30942 34190 30994 34242
rect 31390 34190 31442 34242
rect 34638 34190 34690 34242
rect 47182 34190 47234 34242
rect 54910 34190 54962 34242
rect 56702 34190 56754 34242
rect 7758 34078 7810 34130
rect 8990 34078 9042 34130
rect 10222 34078 10274 34130
rect 16158 34078 16210 34130
rect 17390 34078 17442 34130
rect 20750 34078 20802 34130
rect 23886 34078 23938 34130
rect 28366 34078 28418 34130
rect 28702 34078 28754 34130
rect 28926 34078 28978 34130
rect 30046 34078 30098 34130
rect 30382 34078 30434 34130
rect 30718 34078 30770 34130
rect 31838 34078 31890 34130
rect 34078 34078 34130 34130
rect 36094 34078 36146 34130
rect 36318 34078 36370 34130
rect 37102 34078 37154 34130
rect 39230 34078 39282 34130
rect 39678 34078 39730 34130
rect 40126 34078 40178 34130
rect 41694 34078 41746 34130
rect 42030 34078 42082 34130
rect 43934 34078 43986 34130
rect 44606 34078 44658 34130
rect 45726 34078 45778 34130
rect 45950 34078 46002 34130
rect 55022 34078 55074 34130
rect 57038 34078 57090 34130
rect 57150 34078 57202 34130
rect 9550 33966 9602 34018
rect 11454 33966 11506 34018
rect 16718 33966 16770 34018
rect 19182 33966 19234 34018
rect 21310 33966 21362 34018
rect 23550 33966 23602 34018
rect 25454 33966 25506 34018
rect 27582 33966 27634 34018
rect 28814 33966 28866 34018
rect 31614 33966 31666 34018
rect 33854 33966 33906 34018
rect 37662 33966 37714 34018
rect 38782 33966 38834 34018
rect 41582 33966 41634 34018
rect 46622 33966 46674 34018
rect 46958 33966 47010 34018
rect 47294 33966 47346 34018
rect 47742 33966 47794 34018
rect 56814 33966 56866 34018
rect 9886 33854 9938 33906
rect 36094 33854 36146 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 37550 33518 37602 33570
rect 57038 33518 57090 33570
rect 57598 33518 57650 33570
rect 10894 33406 10946 33458
rect 12686 33406 12738 33458
rect 14142 33406 14194 33458
rect 14590 33406 14642 33458
rect 19406 33406 19458 33458
rect 24222 33406 24274 33458
rect 27918 33406 27970 33458
rect 38110 33406 38162 33458
rect 51214 33406 51266 33458
rect 55582 33406 55634 33458
rect 11230 33294 11282 33346
rect 11678 33294 11730 33346
rect 12238 33294 12290 33346
rect 13022 33294 13074 33346
rect 13806 33294 13858 33346
rect 14814 33294 14866 33346
rect 15822 33294 15874 33346
rect 20190 33294 20242 33346
rect 20638 33294 20690 33346
rect 21422 33294 21474 33346
rect 28142 33294 28194 33346
rect 28366 33294 28418 33346
rect 31838 33294 31890 33346
rect 33630 33294 33682 33346
rect 34302 33294 34354 33346
rect 35086 33294 35138 33346
rect 36990 33294 37042 33346
rect 38446 33294 38498 33346
rect 38894 33294 38946 33346
rect 39790 33294 39842 33346
rect 40238 33294 40290 33346
rect 41246 33294 41298 33346
rect 41694 33294 41746 33346
rect 42030 33294 42082 33346
rect 42366 33294 42418 33346
rect 43934 33294 43986 33346
rect 48302 33294 48354 33346
rect 51886 33294 51938 33346
rect 52782 33294 52834 33346
rect 57150 33294 57202 33346
rect 57486 33294 57538 33346
rect 14254 33182 14306 33234
rect 16718 33182 16770 33234
rect 22094 33182 22146 33234
rect 25790 33182 25842 33234
rect 27806 33182 27858 33234
rect 32398 33182 32450 33234
rect 39118 33182 39170 33234
rect 43710 33182 43762 33234
rect 49086 33182 49138 33234
rect 51550 33182 51602 33234
rect 51998 33182 52050 33234
rect 52110 33182 52162 33234
rect 53454 33182 53506 33234
rect 19966 33070 20018 33122
rect 20078 33070 20130 33122
rect 24670 33070 24722 33122
rect 25118 33070 25170 33122
rect 25454 33070 25506 33122
rect 27582 33070 27634 33122
rect 29486 33070 29538 33122
rect 30942 33070 30994 33122
rect 31278 33070 31330 33122
rect 31502 33070 31554 33122
rect 36206 33070 36258 33122
rect 42030 33070 42082 33122
rect 56030 33070 56082 33122
rect 57038 33070 57090 33122
rect 57598 33070 57650 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 8990 32734 9042 32786
rect 10670 32734 10722 32786
rect 11902 32734 11954 32786
rect 15150 32734 15202 32786
rect 17614 32734 17666 32786
rect 18622 32734 18674 32786
rect 19406 32734 19458 32786
rect 20414 32734 20466 32786
rect 24110 32734 24162 32786
rect 24446 32734 24498 32786
rect 32062 32734 32114 32786
rect 33182 32734 33234 32786
rect 39006 32734 39058 32786
rect 43374 32734 43426 32786
rect 49086 32734 49138 32786
rect 51774 32734 51826 32786
rect 53902 32734 53954 32786
rect 55134 32734 55186 32786
rect 14590 32622 14642 32674
rect 14926 32622 14978 32674
rect 16046 32622 16098 32674
rect 18846 32622 18898 32674
rect 19070 32622 19122 32674
rect 40462 32622 40514 32674
rect 41806 32622 41858 32674
rect 50654 32622 50706 32674
rect 51998 32622 52050 32674
rect 52110 32622 52162 32674
rect 52894 32622 52946 32674
rect 53230 32622 53282 32674
rect 54014 32622 54066 32674
rect 54798 32622 54850 32674
rect 8766 32510 8818 32562
rect 10334 32510 10386 32562
rect 11566 32510 11618 32562
rect 12798 32510 12850 32562
rect 13582 32510 13634 32562
rect 15374 32510 15426 32562
rect 16382 32510 16434 32562
rect 16830 32510 16882 32562
rect 18174 32510 18226 32562
rect 18510 32510 18562 32562
rect 19966 32510 20018 32562
rect 31614 32510 31666 32562
rect 31838 32510 31890 32562
rect 34526 32510 34578 32562
rect 34862 32510 34914 32562
rect 37214 32510 37266 32562
rect 37998 32510 38050 32562
rect 38446 32510 38498 32562
rect 40910 32510 40962 32562
rect 41470 32510 41522 32562
rect 43934 32510 43986 32562
rect 44158 32510 44210 32562
rect 44494 32510 44546 32562
rect 44942 32510 44994 32562
rect 46734 32510 46786 32562
rect 47406 32510 47458 32562
rect 48974 32510 49026 32562
rect 49198 32510 49250 32562
rect 49646 32510 49698 32562
rect 50318 32510 50370 32562
rect 50430 32510 50482 32562
rect 50878 32510 50930 32562
rect 10558 32398 10610 32450
rect 13134 32398 13186 32450
rect 20302 32398 20354 32450
rect 21086 32398 21138 32450
rect 28590 32398 28642 32450
rect 32174 32398 32226 32450
rect 36318 32398 36370 32450
rect 37662 32398 37714 32450
rect 42254 32398 42306 32450
rect 43598 32398 43650 32450
rect 44046 32398 44098 32450
rect 46510 32398 46562 32450
rect 51438 32398 51490 32450
rect 58158 32398 58210 32450
rect 14814 32286 14866 32338
rect 43262 32286 43314 32338
rect 53902 32286 53954 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 35758 31950 35810 32002
rect 43710 31950 43762 32002
rect 44046 31950 44098 32002
rect 49870 31950 49922 32002
rect 7310 31838 7362 31890
rect 8654 31838 8706 31890
rect 12462 31838 12514 31890
rect 14254 31838 14306 31890
rect 18286 31838 18338 31890
rect 18622 31838 18674 31890
rect 19854 31838 19906 31890
rect 26798 31838 26850 31890
rect 30830 31838 30882 31890
rect 32622 31838 32674 31890
rect 34750 31838 34802 31890
rect 37102 31838 37154 31890
rect 39566 31838 39618 31890
rect 41694 31838 41746 31890
rect 42142 31838 42194 31890
rect 45390 31838 45442 31890
rect 56030 31838 56082 31890
rect 58158 31838 58210 31890
rect 7198 31726 7250 31778
rect 8094 31726 8146 31778
rect 8878 31726 8930 31778
rect 10670 31726 10722 31778
rect 11342 31726 11394 31778
rect 12126 31726 12178 31778
rect 12350 31726 12402 31778
rect 13470 31726 13522 31778
rect 13694 31726 13746 31778
rect 13806 31726 13858 31778
rect 15486 31726 15538 31778
rect 19406 31726 19458 31778
rect 23886 31726 23938 31778
rect 31166 31726 31218 31778
rect 32958 31726 33010 31778
rect 33294 31726 33346 31778
rect 34526 31726 34578 31778
rect 35198 31726 35250 31778
rect 35422 31726 35474 31778
rect 37438 31726 37490 31778
rect 37886 31726 37938 31778
rect 38222 31726 38274 31778
rect 38782 31726 38834 31778
rect 44270 31726 44322 31778
rect 48302 31726 48354 31778
rect 49310 31726 49362 31778
rect 50094 31726 50146 31778
rect 55246 31726 55298 31778
rect 16158 31614 16210 31666
rect 24670 31614 24722 31666
rect 47518 31614 47570 31666
rect 49422 31614 49474 31666
rect 49534 31614 49586 31666
rect 15038 31502 15090 31554
rect 27246 31502 27298 31554
rect 48750 31502 48802 31554
rect 50430 31502 50482 31554
rect 50766 31502 50818 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 14030 31166 14082 31218
rect 22542 31166 22594 31218
rect 22766 31166 22818 31218
rect 23326 31166 23378 31218
rect 24110 31166 24162 31218
rect 31054 31166 31106 31218
rect 34526 31166 34578 31218
rect 48974 31166 49026 31218
rect 56926 31166 56978 31218
rect 14478 31054 14530 31106
rect 21982 31054 22034 31106
rect 22094 31054 22146 31106
rect 43038 31054 43090 31106
rect 49982 31054 50034 31106
rect 55358 31054 55410 31106
rect 57822 31054 57874 31106
rect 58158 31054 58210 31106
rect 7198 30942 7250 30994
rect 9998 30942 10050 30994
rect 11790 30942 11842 30994
rect 13918 30942 13970 30994
rect 21534 30942 21586 30994
rect 22318 30942 22370 30994
rect 22878 30942 22930 30994
rect 23102 30942 23154 30994
rect 23438 30942 23490 30994
rect 23998 30942 24050 30994
rect 24334 30942 24386 30994
rect 28142 30942 28194 30994
rect 42366 30942 42418 30994
rect 55134 30942 55186 30994
rect 56590 30942 56642 30994
rect 56814 30942 56866 30994
rect 57262 30942 57314 30994
rect 12238 30830 12290 30882
rect 15710 30830 15762 30882
rect 21198 30830 21250 30882
rect 22094 30830 22146 30882
rect 25454 30830 25506 30882
rect 27694 30830 27746 30882
rect 28814 30830 28866 30882
rect 45166 30830 45218 30882
rect 45614 30830 45666 30882
rect 49870 30830 49922 30882
rect 7758 30718 7810 30770
rect 11566 30718 11618 30770
rect 50206 30718 50258 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 46510 30382 46562 30434
rect 11342 30270 11394 30322
rect 16046 30270 16098 30322
rect 21534 30270 21586 30322
rect 25006 30270 25058 30322
rect 28590 30270 28642 30322
rect 29150 30270 29202 30322
rect 31950 30270 32002 30322
rect 32510 30270 32562 30322
rect 35086 30270 35138 30322
rect 39902 30270 39954 30322
rect 46958 30270 47010 30322
rect 56030 30270 56082 30322
rect 58158 30270 58210 30322
rect 8206 30158 8258 30210
rect 9662 30158 9714 30210
rect 13582 30158 13634 30210
rect 13806 30158 13858 30210
rect 14142 30158 14194 30210
rect 19070 30158 19122 30210
rect 19630 30158 19682 30210
rect 22318 30158 22370 30210
rect 25790 30158 25842 30210
rect 30158 30158 30210 30210
rect 34302 30158 34354 30210
rect 34638 30158 34690 30210
rect 35758 30158 35810 30210
rect 37102 30158 37154 30210
rect 46622 30158 46674 30210
rect 49870 30158 49922 30210
rect 50206 30158 50258 30210
rect 50878 30158 50930 30210
rect 51550 30158 51602 30210
rect 52670 30158 52722 30210
rect 55358 30158 55410 30210
rect 10110 30046 10162 30098
rect 16382 30046 16434 30098
rect 16494 30046 16546 30098
rect 17054 30046 17106 30098
rect 17278 30046 17330 30098
rect 17390 30046 17442 30098
rect 21758 30046 21810 30098
rect 21982 30046 22034 30098
rect 22094 30046 22146 30098
rect 24222 30046 24274 30098
rect 24558 30046 24610 30098
rect 24782 30046 24834 30098
rect 26462 30046 26514 30098
rect 29486 30046 29538 30098
rect 29598 30046 29650 30098
rect 30382 30046 30434 30098
rect 30494 30046 30546 30098
rect 31166 30046 31218 30098
rect 31278 30046 31330 30098
rect 33294 30046 33346 30098
rect 37774 30046 37826 30098
rect 49086 30046 49138 30098
rect 51774 30046 51826 30098
rect 7758 29934 7810 29986
rect 9662 29934 9714 29986
rect 14814 29934 14866 29986
rect 16606 29934 16658 29986
rect 16830 29934 16882 29986
rect 17838 29934 17890 29986
rect 22878 29934 22930 29986
rect 24446 29934 24498 29986
rect 29710 29934 29762 29986
rect 29934 29934 29986 29986
rect 31502 29934 31554 29986
rect 35534 29934 35586 29986
rect 36542 29934 36594 29986
rect 40350 29934 40402 29986
rect 46510 29934 46562 29986
rect 50318 29934 50370 29986
rect 50542 29934 50594 29986
rect 53006 29934 53058 29986
rect 54574 29934 54626 29986
rect 54910 29934 54962 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 10446 29598 10498 29650
rect 20414 29598 20466 29650
rect 21870 29598 21922 29650
rect 22318 29598 22370 29650
rect 23214 29598 23266 29650
rect 24334 29598 24386 29650
rect 25566 29598 25618 29650
rect 26910 29598 26962 29650
rect 27806 29598 27858 29650
rect 28030 29598 28082 29650
rect 28702 29598 28754 29650
rect 34414 29598 34466 29650
rect 34750 29598 34802 29650
rect 35310 29598 35362 29650
rect 37214 29598 37266 29650
rect 42926 29598 42978 29650
rect 43486 29598 43538 29650
rect 51102 29598 51154 29650
rect 53118 29598 53170 29650
rect 56702 29598 56754 29650
rect 56926 29598 56978 29650
rect 57822 29598 57874 29650
rect 9774 29486 9826 29538
rect 11342 29486 11394 29538
rect 12350 29486 12402 29538
rect 21534 29486 21586 29538
rect 21646 29486 21698 29538
rect 22094 29486 22146 29538
rect 22430 29486 22482 29538
rect 22878 29486 22930 29538
rect 23662 29486 23714 29538
rect 25230 29486 25282 29538
rect 27582 29486 27634 29538
rect 27694 29486 27746 29538
rect 28478 29486 28530 29538
rect 30718 29486 30770 29538
rect 30942 29486 30994 29538
rect 31278 29486 31330 29538
rect 51550 29486 51602 29538
rect 53454 29486 53506 29538
rect 57038 29486 57090 29538
rect 4286 29374 4338 29426
rect 7758 29374 7810 29426
rect 9550 29374 9602 29426
rect 10558 29374 10610 29426
rect 13470 29374 13522 29426
rect 14254 29374 14306 29426
rect 15150 29374 15202 29426
rect 15598 29374 15650 29426
rect 17390 29374 17442 29426
rect 21086 29374 21138 29426
rect 23998 29374 24050 29426
rect 24558 29374 24610 29426
rect 28814 29374 28866 29426
rect 31166 29374 31218 29426
rect 35646 29374 35698 29426
rect 36878 29374 36930 29426
rect 36990 29374 37042 29426
rect 37438 29374 37490 29426
rect 50990 29374 51042 29426
rect 51214 29374 51266 29426
rect 5070 29262 5122 29314
rect 7198 29262 7250 29314
rect 8542 29262 8594 29314
rect 11006 29262 11058 29314
rect 18174 29262 18226 29314
rect 21534 29262 21586 29314
rect 27694 29262 27746 29314
rect 29262 29262 29314 29314
rect 29710 29262 29762 29314
rect 31502 29262 31554 29314
rect 31950 29262 32002 29314
rect 35982 29262 36034 29314
rect 40238 29262 40290 29314
rect 44046 29262 44098 29314
rect 53902 29262 53954 29314
rect 58158 29262 58210 29314
rect 13470 29150 13522 29202
rect 40126 29150 40178 29202
rect 42814 29150 42866 29202
rect 43150 29150 43202 29202
rect 43822 29150 43874 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 18174 28814 18226 28866
rect 9102 28702 9154 28754
rect 11118 28702 11170 28754
rect 13470 28702 13522 28754
rect 14926 28702 14978 28754
rect 15822 28702 15874 28754
rect 19630 28702 19682 28754
rect 31950 28702 32002 28754
rect 34078 28702 34130 28754
rect 37886 28702 37938 28754
rect 41470 28702 41522 28754
rect 41918 28702 41970 28754
rect 43486 28702 43538 28754
rect 45278 28702 45330 28754
rect 48526 28702 48578 28754
rect 49534 28702 49586 28754
rect 49758 28702 49810 28754
rect 50654 28702 50706 28754
rect 56590 28702 56642 28754
rect 6974 28590 7026 28642
rect 7310 28590 7362 28642
rect 12910 28590 12962 28642
rect 15374 28590 15426 28642
rect 16606 28590 16658 28642
rect 17390 28590 17442 28642
rect 18062 28590 18114 28642
rect 19182 28590 19234 28642
rect 30270 28590 30322 28642
rect 30606 28590 30658 28642
rect 30942 28590 30994 28642
rect 31166 28590 31218 28642
rect 34862 28590 34914 28642
rect 35310 28590 35362 28642
rect 35870 28590 35922 28642
rect 37326 28590 37378 28642
rect 38670 28590 38722 28642
rect 42702 28590 42754 28642
rect 43038 28590 43090 28642
rect 45614 28590 45666 28642
rect 52782 28590 52834 28642
rect 53230 28590 53282 28642
rect 54238 28590 54290 28642
rect 7870 28478 7922 28530
rect 12350 28478 12402 28530
rect 13694 28478 13746 28530
rect 13918 28478 13970 28530
rect 14814 28478 14866 28530
rect 14926 28478 14978 28530
rect 17502 28478 17554 28530
rect 18174 28478 18226 28530
rect 18846 28478 18898 28530
rect 30718 28478 30770 28530
rect 36094 28478 36146 28530
rect 37774 28478 37826 28530
rect 37998 28478 38050 28530
rect 39342 28478 39394 28530
rect 46398 28478 46450 28530
rect 53566 28478 53618 28530
rect 7422 28366 7474 28418
rect 12798 28366 12850 28418
rect 14030 28366 14082 28418
rect 14254 28366 14306 28418
rect 14590 28366 14642 28418
rect 16942 28366 16994 28418
rect 17054 28366 17106 28418
rect 17166 28366 17218 28418
rect 20750 28366 20802 28418
rect 43374 28366 43426 28418
rect 43598 28366 43650 28418
rect 50094 28366 50146 28418
rect 53006 28366 53058 28418
rect 53454 28366 53506 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 8654 28030 8706 28082
rect 13246 28030 13298 28082
rect 14478 28030 14530 28082
rect 15038 28030 15090 28082
rect 15822 28030 15874 28082
rect 18174 28030 18226 28082
rect 28254 28030 28306 28082
rect 29038 28030 29090 28082
rect 30830 28030 30882 28082
rect 35086 28030 35138 28082
rect 35758 28030 35810 28082
rect 38894 28030 38946 28082
rect 44382 28030 44434 28082
rect 54686 28030 54738 28082
rect 56590 28030 56642 28082
rect 57374 28030 57426 28082
rect 11454 27918 11506 27970
rect 14702 27918 14754 27970
rect 15262 27918 15314 27970
rect 20302 27918 20354 27970
rect 31054 27918 31106 27970
rect 32062 27918 32114 27970
rect 38110 27918 38162 27970
rect 38222 27918 38274 27970
rect 38446 27918 38498 27970
rect 39006 27918 39058 27970
rect 39118 27918 39170 27970
rect 41806 27918 41858 27970
rect 55470 27918 55522 27970
rect 56926 27918 56978 27970
rect 57262 27918 57314 27970
rect 57934 27918 57986 27970
rect 4734 27806 4786 27858
rect 7982 27806 8034 27858
rect 12126 27806 12178 27858
rect 13134 27806 13186 27858
rect 13470 27806 13522 27858
rect 14814 27806 14866 27858
rect 15374 27806 15426 27858
rect 19630 27806 19682 27858
rect 22878 27806 22930 27858
rect 25790 27806 25842 27858
rect 28702 27806 28754 27858
rect 31278 27806 31330 27858
rect 31502 27806 31554 27858
rect 32510 27806 32562 27858
rect 34526 27806 34578 27858
rect 38670 27806 38722 27858
rect 41134 27806 41186 27858
rect 51438 27806 51490 27858
rect 55134 27806 55186 27858
rect 57822 27806 57874 27858
rect 5406 27694 5458 27746
rect 7534 27694 7586 27746
rect 9662 27694 9714 27746
rect 12350 27694 12402 27746
rect 18622 27694 18674 27746
rect 22430 27694 22482 27746
rect 26350 27694 26402 27746
rect 31614 27694 31666 27746
rect 37774 27694 37826 27746
rect 39454 27694 39506 27746
rect 43934 27694 43986 27746
rect 52110 27694 52162 27746
rect 54238 27694 54290 27746
rect 57374 27582 57426 27634
rect 57934 27582 57986 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 7870 27246 7922 27298
rect 8542 27246 8594 27298
rect 24558 27246 24610 27298
rect 12238 27134 12290 27186
rect 13918 27134 13970 27186
rect 15710 27134 15762 27186
rect 18510 27134 18562 27186
rect 29374 27134 29426 27186
rect 31726 27134 31778 27186
rect 33854 27134 33906 27186
rect 38670 27134 38722 27186
rect 40014 27134 40066 27186
rect 41918 27134 41970 27186
rect 58158 27134 58210 27186
rect 6750 27022 6802 27074
rect 7422 27022 7474 27074
rect 9326 27022 9378 27074
rect 11006 27022 11058 27074
rect 11566 27022 11618 27074
rect 14702 27022 14754 27074
rect 15262 27022 15314 27074
rect 25902 27022 25954 27074
rect 26126 27022 26178 27074
rect 26798 27022 26850 27074
rect 28030 27022 28082 27074
rect 30606 27022 30658 27074
rect 30942 27022 30994 27074
rect 37998 27022 38050 27074
rect 40910 27022 40962 27074
rect 45054 27022 45106 27074
rect 52558 27022 52610 27074
rect 53230 27022 53282 27074
rect 53790 27022 53842 27074
rect 55358 27022 55410 27074
rect 6974 26910 7026 26962
rect 10110 26910 10162 26962
rect 13470 26910 13522 26962
rect 14366 26910 14418 26962
rect 15150 26910 15202 26962
rect 24670 26910 24722 26962
rect 25678 26910 25730 26962
rect 26462 26910 26514 26962
rect 38222 26910 38274 26962
rect 44270 26910 44322 26962
rect 44830 26910 44882 26962
rect 45390 26910 45442 26962
rect 52782 26910 52834 26962
rect 53006 26910 53058 26962
rect 53454 26910 53506 26962
rect 56030 26910 56082 26962
rect 14926 26798 14978 26850
rect 18174 26798 18226 26850
rect 18398 26798 18450 26850
rect 24558 26798 24610 26850
rect 25454 26798 25506 26850
rect 25566 26798 25618 26850
rect 26574 26798 26626 26850
rect 27806 26798 27858 26850
rect 28366 26798 28418 26850
rect 29822 26798 29874 26850
rect 43934 26798 43986 26850
rect 44158 26798 44210 26850
rect 44942 26798 44994 26850
rect 53678 26798 53730 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 9550 26462 9602 26514
rect 10670 26462 10722 26514
rect 11566 26462 11618 26514
rect 11790 26462 11842 26514
rect 15598 26462 15650 26514
rect 15934 26462 15986 26514
rect 18174 26462 18226 26514
rect 25118 26462 25170 26514
rect 25342 26462 25394 26514
rect 26462 26462 26514 26514
rect 27358 26462 27410 26514
rect 28478 26462 28530 26514
rect 29038 26462 29090 26514
rect 30270 26462 30322 26514
rect 30830 26462 30882 26514
rect 34414 26462 34466 26514
rect 37662 26462 37714 26514
rect 39230 26462 39282 26514
rect 40126 26462 40178 26514
rect 41918 26462 41970 26514
rect 52334 26462 52386 26514
rect 57038 26462 57090 26514
rect 12350 26350 12402 26402
rect 16494 26350 16546 26402
rect 17390 26350 17442 26402
rect 18062 26350 18114 26402
rect 18622 26350 18674 26402
rect 25454 26350 25506 26402
rect 28814 26350 28866 26402
rect 29598 26350 29650 26402
rect 33966 26350 34018 26402
rect 39790 26350 39842 26402
rect 41470 26350 41522 26402
rect 52558 26350 52610 26402
rect 52670 26350 52722 26402
rect 8766 26238 8818 26290
rect 10446 26238 10498 26290
rect 11118 26238 11170 26290
rect 13246 26238 13298 26290
rect 16830 26238 16882 26290
rect 17726 26238 17778 26290
rect 19182 26238 19234 26290
rect 22766 26238 22818 26290
rect 23774 26238 23826 26290
rect 26126 26238 26178 26290
rect 26350 26238 26402 26290
rect 26574 26238 26626 26290
rect 27134 26238 27186 26290
rect 27470 26238 27522 26290
rect 28254 26238 28306 26290
rect 28590 26238 28642 26290
rect 29150 26238 29202 26290
rect 30158 26238 30210 26290
rect 39454 26238 39506 26290
rect 41134 26238 41186 26290
rect 42590 26238 42642 26290
rect 47630 26238 47682 26290
rect 48190 26238 48242 26290
rect 56590 26238 56642 26290
rect 56926 26238 56978 26290
rect 57262 26238 57314 26290
rect 5630 26126 5682 26178
rect 7870 26126 7922 26178
rect 9998 26126 10050 26178
rect 10558 26126 10610 26178
rect 15038 26126 15090 26178
rect 22318 26126 22370 26178
rect 23214 26126 23266 26178
rect 24110 26126 24162 26178
rect 24334 26126 24386 26178
rect 27246 26126 27298 26178
rect 36766 26126 36818 26178
rect 43262 26126 43314 26178
rect 45390 26126 45442 26178
rect 58158 26126 58210 26178
rect 18174 26014 18226 26066
rect 25902 26014 25954 26066
rect 27806 26014 27858 26066
rect 29486 26014 29538 26066
rect 30270 26014 30322 26066
rect 33854 26014 33906 26066
rect 39118 26014 39170 26066
rect 41022 26014 41074 26066
rect 41358 26014 41410 26066
rect 47294 26014 47346 26066
rect 47630 26014 47682 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 24110 25678 24162 25730
rect 33182 25678 33234 25730
rect 39790 25678 39842 25730
rect 39902 25678 39954 25730
rect 40686 25678 40738 25730
rect 43598 25678 43650 25730
rect 43934 25678 43986 25730
rect 44046 25678 44098 25730
rect 11566 25566 11618 25618
rect 13918 25566 13970 25618
rect 15822 25566 15874 25618
rect 19966 25566 20018 25618
rect 23326 25566 23378 25618
rect 26126 25566 26178 25618
rect 26686 25566 26738 25618
rect 27694 25566 27746 25618
rect 28590 25566 28642 25618
rect 33854 25566 33906 25618
rect 34190 25566 34242 25618
rect 36206 25566 36258 25618
rect 39006 25566 39058 25618
rect 39342 25566 39394 25618
rect 45166 25566 45218 25618
rect 46958 25566 47010 25618
rect 49086 25566 49138 25618
rect 50318 25566 50370 25618
rect 7646 25454 7698 25506
rect 7982 25454 8034 25506
rect 8206 25454 8258 25506
rect 8654 25454 8706 25506
rect 12126 25454 12178 25506
rect 14030 25454 14082 25506
rect 14702 25454 14754 25506
rect 16606 25454 16658 25506
rect 16830 25454 16882 25506
rect 24222 25454 24274 25506
rect 24558 25454 24610 25506
rect 25566 25454 25618 25506
rect 25902 25454 25954 25506
rect 26014 25454 26066 25506
rect 26238 25454 26290 25506
rect 26910 25454 26962 25506
rect 27806 25454 27858 25506
rect 29710 25454 29762 25506
rect 32398 25454 32450 25506
rect 32734 25454 32786 25506
rect 33294 25454 33346 25506
rect 34974 25454 35026 25506
rect 35758 25454 35810 25506
rect 36990 25454 37042 25506
rect 38446 25454 38498 25506
rect 40126 25454 40178 25506
rect 41918 25454 41970 25506
rect 43710 25454 43762 25506
rect 45054 25454 45106 25506
rect 45726 25454 45778 25506
rect 45950 25454 46002 25506
rect 46622 25454 46674 25506
rect 49870 25454 49922 25506
rect 52558 25454 52610 25506
rect 53006 25454 53058 25506
rect 53454 25454 53506 25506
rect 53790 25454 53842 25506
rect 56702 25454 56754 25506
rect 9326 25342 9378 25394
rect 14366 25342 14418 25394
rect 16046 25342 16098 25394
rect 16270 25342 16322 25394
rect 17726 25342 17778 25394
rect 21422 25342 21474 25394
rect 21758 25342 21810 25394
rect 21982 25342 22034 25394
rect 24110 25342 24162 25394
rect 24670 25342 24722 25394
rect 27358 25342 27410 25394
rect 29486 25342 29538 25394
rect 29822 25342 29874 25394
rect 30942 25342 30994 25394
rect 32622 25342 32674 25394
rect 34638 25342 34690 25394
rect 35422 25342 35474 25394
rect 37326 25342 37378 25394
rect 37550 25342 37602 25394
rect 38334 25342 38386 25394
rect 39230 25342 39282 25394
rect 40238 25342 40290 25394
rect 40574 25342 40626 25394
rect 40686 25342 40738 25394
rect 42478 25342 42530 25394
rect 44830 25342 44882 25394
rect 45278 25342 45330 25394
rect 53230 25342 53282 25394
rect 53678 25342 53730 25394
rect 56590 25342 56642 25394
rect 58158 25342 58210 25394
rect 7870 25230 7922 25282
rect 12238 25230 12290 25282
rect 12462 25230 12514 25282
rect 12798 25230 12850 25282
rect 13582 25230 13634 25282
rect 14478 25230 14530 25282
rect 15598 25230 15650 25282
rect 16382 25230 16434 25282
rect 21534 25230 21586 25282
rect 22542 25230 22594 25282
rect 31278 25230 31330 25282
rect 33182 25230 33234 25282
rect 34078 25230 34130 25282
rect 37102 25230 37154 25282
rect 37998 25230 38050 25282
rect 38222 25230 38274 25282
rect 41470 25230 41522 25282
rect 41694 25230 41746 25282
rect 42926 25230 42978 25282
rect 52782 25230 52834 25282
rect 56366 25230 56418 25282
rect 57598 25230 57650 25282
rect 57822 25230 57874 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 8430 24894 8482 24946
rect 8878 24894 8930 24946
rect 13470 24894 13522 24946
rect 14702 24894 14754 24946
rect 15150 24894 15202 24946
rect 16158 24894 16210 24946
rect 16270 24894 16322 24946
rect 17390 24894 17442 24946
rect 19182 24894 19234 24946
rect 25566 24894 25618 24946
rect 26126 24894 26178 24946
rect 27134 24894 27186 24946
rect 28142 24894 28194 24946
rect 29934 24894 29986 24946
rect 31390 24894 31442 24946
rect 39230 24894 39282 24946
rect 45838 24894 45890 24946
rect 46174 24894 46226 24946
rect 52558 24894 52610 24946
rect 56814 24894 56866 24946
rect 14478 24782 14530 24834
rect 16494 24782 16546 24834
rect 16606 24782 16658 24834
rect 17614 24782 17666 24834
rect 20526 24782 20578 24834
rect 25342 24782 25394 24834
rect 25902 24782 25954 24834
rect 27694 24782 27746 24834
rect 28926 24782 28978 24834
rect 36094 24782 36146 24834
rect 40910 24782 40962 24834
rect 41134 24782 41186 24834
rect 42142 24782 42194 24834
rect 50206 24782 50258 24834
rect 52782 24782 52834 24834
rect 57822 24782 57874 24834
rect 10222 24670 10274 24722
rect 14030 24670 14082 24722
rect 14254 24670 14306 24722
rect 17838 24670 17890 24722
rect 18174 24670 18226 24722
rect 19742 24670 19794 24722
rect 23438 24670 23490 24722
rect 25230 24670 25282 24722
rect 25790 24670 25842 24722
rect 27470 24670 27522 24722
rect 28702 24670 28754 24722
rect 29150 24670 29202 24722
rect 29486 24670 29538 24722
rect 32958 24670 33010 24722
rect 33294 24670 33346 24722
rect 33630 24670 33682 24722
rect 34190 24670 34242 24722
rect 35422 24670 35474 24722
rect 41806 24670 41858 24722
rect 42702 24670 42754 24722
rect 43150 24670 43202 24722
rect 49534 24670 49586 24722
rect 52894 24670 52946 24722
rect 56478 24670 56530 24722
rect 56926 24670 56978 24722
rect 57150 24670 57202 24722
rect 10894 24558 10946 24610
rect 13022 24558 13074 24610
rect 14366 24558 14418 24610
rect 15598 24558 15650 24610
rect 17726 24558 17778 24610
rect 18622 24558 18674 24610
rect 22654 24558 22706 24610
rect 23102 24558 23154 24610
rect 23998 24558 24050 24610
rect 29038 24558 29090 24610
rect 31838 24558 31890 24610
rect 38222 24558 38274 24610
rect 38670 24558 38722 24610
rect 41022 24558 41074 24610
rect 43598 24558 43650 24610
rect 44382 24558 44434 24610
rect 44830 24558 44882 24610
rect 45278 24558 45330 24610
rect 52334 24558 52386 24610
rect 53342 24558 53394 24610
rect 57486 24558 57538 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 31502 24110 31554 24162
rect 19406 23998 19458 24050
rect 22318 23998 22370 24050
rect 27694 23998 27746 24050
rect 29150 23998 29202 24050
rect 38446 23998 38498 24050
rect 55134 23998 55186 24050
rect 57262 23998 57314 24050
rect 18958 23886 19010 23938
rect 19854 23886 19906 23938
rect 20302 23886 20354 23938
rect 22206 23886 22258 23938
rect 22878 23886 22930 23938
rect 24894 23886 24946 23938
rect 26910 23886 26962 23938
rect 28030 23886 28082 23938
rect 33742 23886 33794 23938
rect 35758 23886 35810 23938
rect 45502 23886 45554 23938
rect 46174 23886 46226 23938
rect 52670 23886 52722 23938
rect 53230 23886 53282 23938
rect 53790 23886 53842 23938
rect 54126 23886 54178 23938
rect 54462 23886 54514 23938
rect 58046 23886 58098 23938
rect 24334 23774 24386 23826
rect 26350 23774 26402 23826
rect 28254 23774 28306 23826
rect 31614 23774 31666 23826
rect 35982 23774 36034 23826
rect 52894 23774 52946 23826
rect 53454 23774 53506 23826
rect 53678 23774 53730 23826
rect 16606 23662 16658 23714
rect 20750 23662 20802 23714
rect 21982 23662 22034 23714
rect 22430 23662 22482 23714
rect 26798 23662 26850 23714
rect 29262 23662 29314 23714
rect 32062 23662 32114 23714
rect 33518 23662 33570 23714
rect 44942 23662 44994 23714
rect 45838 23662 45890 23714
rect 46510 23662 46562 23714
rect 46622 23662 46674 23714
rect 46734 23662 46786 23714
rect 53006 23662 53058 23714
rect 54238 23662 54290 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 19630 23326 19682 23378
rect 23438 23326 23490 23378
rect 24334 23326 24386 23378
rect 25342 23326 25394 23378
rect 27582 23326 27634 23378
rect 42142 23326 42194 23378
rect 42478 23326 42530 23378
rect 43150 23326 43202 23378
rect 44158 23326 44210 23378
rect 44606 23326 44658 23378
rect 56702 23326 56754 23378
rect 56926 23326 56978 23378
rect 15934 23214 15986 23266
rect 30046 23214 30098 23266
rect 39230 23214 39282 23266
rect 44942 23214 44994 23266
rect 51438 23214 51490 23266
rect 54014 23214 54066 23266
rect 54126 23214 54178 23266
rect 54350 23214 54402 23266
rect 56590 23214 56642 23266
rect 16718 23102 16770 23154
rect 22318 23102 22370 23154
rect 22654 23102 22706 23154
rect 22990 23102 23042 23154
rect 23662 23102 23714 23154
rect 24110 23102 24162 23154
rect 24222 23102 24274 23154
rect 25230 23102 25282 23154
rect 30718 23102 30770 23154
rect 33630 23102 33682 23154
rect 34078 23102 34130 23154
rect 38110 23102 38162 23154
rect 38558 23102 38610 23154
rect 38782 23102 38834 23154
rect 41022 23102 41074 23154
rect 42030 23102 42082 23154
rect 42254 23102 42306 23154
rect 45390 23102 45442 23154
rect 50766 23102 50818 23154
rect 13806 22990 13858 23042
rect 17502 22990 17554 23042
rect 22542 22990 22594 23042
rect 27918 22990 27970 23042
rect 33070 22990 33122 23042
rect 38334 22990 38386 23042
rect 43710 22990 43762 23042
rect 46062 22990 46114 23042
rect 48190 22990 48242 23042
rect 53566 22990 53618 23042
rect 54686 22990 54738 23042
rect 58158 22990 58210 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 33182 22430 33234 22482
rect 36430 22430 36482 22482
rect 40686 22430 40738 22482
rect 44158 22430 44210 22482
rect 45054 22430 45106 22482
rect 45502 22430 45554 22482
rect 45838 22430 45890 22482
rect 47518 22430 47570 22482
rect 50766 22430 50818 22482
rect 51214 22430 51266 22482
rect 24446 22318 24498 22370
rect 26462 22318 26514 22370
rect 26910 22318 26962 22370
rect 33518 22318 33570 22370
rect 37886 22318 37938 22370
rect 38558 22318 38610 22370
rect 41246 22318 41298 22370
rect 45614 22318 45666 22370
rect 45950 22318 46002 22370
rect 46286 22318 46338 22370
rect 46734 22318 46786 22370
rect 47966 22318 48018 22370
rect 54910 22318 54962 22370
rect 56814 22318 56866 22370
rect 57374 22318 57426 22370
rect 57934 22318 57986 22370
rect 23886 22206 23938 22258
rect 25342 22206 25394 22258
rect 27918 22206 27970 22258
rect 34302 22206 34354 22258
rect 37214 22206 37266 22258
rect 37326 22206 37378 22258
rect 37438 22206 37490 22258
rect 42030 22206 42082 22258
rect 47070 22206 47122 22258
rect 47182 22206 47234 22258
rect 48638 22206 48690 22258
rect 54574 22206 54626 22258
rect 55134 22206 55186 22258
rect 56702 22206 56754 22258
rect 57038 22206 57090 22258
rect 28478 22094 28530 22146
rect 46958 22094 47010 22146
rect 54686 22094 54738 22146
rect 56478 22094 56530 22146
rect 57262 22094 57314 22146
rect 57598 22094 57650 22146
rect 57822 22094 57874 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 18622 21758 18674 21810
rect 19294 21758 19346 21810
rect 19966 21758 20018 21810
rect 25342 21758 25394 21810
rect 33630 21758 33682 21810
rect 34414 21758 34466 21810
rect 35534 21758 35586 21810
rect 36766 21758 36818 21810
rect 40350 21758 40402 21810
rect 41470 21758 41522 21810
rect 46398 21758 46450 21810
rect 47070 21758 47122 21810
rect 47294 21758 47346 21810
rect 49646 21758 49698 21810
rect 18286 21646 18338 21698
rect 18958 21646 19010 21698
rect 19630 21646 19682 21698
rect 22430 21646 22482 21698
rect 26350 21646 26402 21698
rect 27806 21646 27858 21698
rect 33966 21646 34018 21698
rect 35758 21646 35810 21698
rect 36094 21646 36146 21698
rect 37102 21646 37154 21698
rect 38110 21646 38162 21698
rect 41582 21646 41634 21698
rect 41806 21646 41858 21698
rect 49758 21646 49810 21698
rect 54350 21646 54402 21698
rect 56926 21646 56978 21698
rect 57150 21646 57202 21698
rect 21758 21534 21810 21586
rect 26798 21534 26850 21586
rect 27246 21534 27298 21586
rect 34302 21534 34354 21586
rect 34526 21534 34578 21586
rect 34862 21534 34914 21586
rect 35086 21534 35138 21586
rect 35646 21534 35698 21586
rect 36318 21534 36370 21586
rect 37774 21534 37826 21586
rect 38334 21534 38386 21586
rect 39006 21534 39058 21586
rect 41134 21534 41186 21586
rect 47406 21534 47458 21586
rect 55134 21534 55186 21586
rect 55582 21534 55634 21586
rect 56478 21534 56530 21586
rect 24558 21422 24610 21474
rect 45390 21422 45442 21474
rect 47854 21422 47906 21474
rect 52222 21422 52274 21474
rect 56702 21422 56754 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 18062 20862 18114 20914
rect 19406 20862 19458 20914
rect 22766 20862 22818 20914
rect 24894 20862 24946 20914
rect 29262 20862 29314 20914
rect 30158 20862 30210 20914
rect 33518 20862 33570 20914
rect 56030 20862 56082 20914
rect 58158 20862 58210 20914
rect 15262 20750 15314 20802
rect 18286 20750 18338 20802
rect 18734 20750 18786 20802
rect 18846 20750 18898 20802
rect 20078 20750 20130 20802
rect 20526 20750 20578 20802
rect 22430 20750 22482 20802
rect 27918 20750 27970 20802
rect 29374 20750 29426 20802
rect 30718 20750 30770 20802
rect 33966 20750 34018 20802
rect 55246 20750 55298 20802
rect 15934 20638 15986 20690
rect 18510 20638 18562 20690
rect 20750 20638 20802 20690
rect 21870 20638 21922 20690
rect 29150 20638 29202 20690
rect 29710 20638 29762 20690
rect 31390 20638 31442 20690
rect 14814 20526 14866 20578
rect 20302 20526 20354 20578
rect 21758 20526 21810 20578
rect 21982 20526 22034 20578
rect 28254 20526 28306 20578
rect 41582 20526 41634 20578
rect 47294 20526 47346 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 18510 20190 18562 20242
rect 31278 20190 31330 20242
rect 37774 20190 37826 20242
rect 58158 20190 58210 20242
rect 18398 20078 18450 20130
rect 20190 20078 20242 20130
rect 26798 20078 26850 20130
rect 27470 20078 27522 20130
rect 28590 20078 28642 20130
rect 31614 20078 31666 20130
rect 32062 20078 32114 20130
rect 32398 20078 32450 20130
rect 40350 20078 40402 20130
rect 41246 20078 41298 20130
rect 46622 20078 46674 20130
rect 47966 20078 48018 20130
rect 18062 19966 18114 20018
rect 18622 19966 18674 20018
rect 18958 19966 19010 20018
rect 19406 19966 19458 20018
rect 26574 19966 26626 20018
rect 27246 19966 27298 20018
rect 27918 19966 27970 20018
rect 31054 19966 31106 20018
rect 31390 19966 31442 20018
rect 31950 19966 32002 20018
rect 32174 19966 32226 20018
rect 40910 19966 40962 20018
rect 41470 19966 41522 20018
rect 41806 19966 41858 20018
rect 46846 19966 46898 20018
rect 47070 19966 47122 20018
rect 47518 19966 47570 20018
rect 47742 19966 47794 20018
rect 22318 19854 22370 19906
rect 30718 19854 30770 19906
rect 41022 19854 41074 19906
rect 42590 19854 42642 19906
rect 44718 19854 44770 19906
rect 46286 19854 46338 19906
rect 46734 19854 46786 19906
rect 47630 19854 47682 19906
rect 50318 19854 50370 19906
rect 51214 19854 51266 19906
rect 50094 19742 50146 19794
rect 50318 19742 50370 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 17166 19294 17218 19346
rect 17726 19294 17778 19346
rect 26238 19294 26290 19346
rect 30046 19294 30098 19346
rect 30942 19294 30994 19346
rect 34190 19294 34242 19346
rect 39790 19294 39842 19346
rect 42142 19294 42194 19346
rect 47854 19294 47906 19346
rect 49982 19294 50034 19346
rect 14366 19182 14418 19234
rect 18286 19182 18338 19234
rect 18958 19182 19010 19234
rect 23662 19182 23714 19234
rect 24334 19182 24386 19234
rect 26574 19182 26626 19234
rect 26798 19182 26850 19234
rect 30606 19182 30658 19234
rect 33742 19182 33794 19234
rect 35422 19182 35474 19234
rect 36990 19182 37042 19234
rect 37214 19182 37266 19234
rect 37550 19182 37602 19234
rect 37998 19182 38050 19234
rect 38782 19182 38834 19234
rect 39118 19182 39170 19234
rect 42254 19182 42306 19234
rect 45614 19182 45666 19234
rect 46174 19182 46226 19234
rect 47182 19182 47234 19234
rect 50430 19182 50482 19234
rect 15038 19070 15090 19122
rect 27134 19070 27186 19122
rect 39342 19070 39394 19122
rect 45950 19070 46002 19122
rect 50878 19070 50930 19122
rect 51102 19070 51154 19122
rect 18398 18958 18450 19010
rect 18510 18958 18562 19010
rect 23998 18958 24050 19010
rect 26686 18958 26738 19010
rect 29934 18958 29986 19010
rect 30158 18958 30210 19010
rect 34638 18958 34690 19010
rect 34974 18958 35026 19010
rect 35982 18958 36034 19010
rect 37102 18958 37154 19010
rect 37886 18958 37938 19010
rect 38110 18958 38162 19010
rect 38334 18958 38386 19010
rect 38894 18958 38946 19010
rect 41806 18958 41858 19010
rect 42030 18958 42082 19010
rect 45278 18958 45330 19010
rect 45838 18958 45890 19010
rect 50766 18958 50818 19010
rect 51438 18958 51490 19010
rect 51550 18958 51602 19010
rect 51662 18958 51714 19010
rect 51886 18958 51938 19010
rect 52782 18958 52834 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 21758 18622 21810 18674
rect 28478 18622 28530 18674
rect 33854 18622 33906 18674
rect 39566 18622 39618 18674
rect 39678 18622 39730 18674
rect 41246 18622 41298 18674
rect 18510 18510 18562 18562
rect 24446 18510 24498 18562
rect 26014 18510 26066 18562
rect 28702 18510 28754 18562
rect 39790 18510 39842 18562
rect 42142 18510 42194 18562
rect 45838 18510 45890 18562
rect 50878 18510 50930 18562
rect 52558 18510 52610 18562
rect 17950 18398 18002 18450
rect 18062 18398 18114 18450
rect 18286 18398 18338 18450
rect 19070 18398 19122 18450
rect 21982 18398 22034 18450
rect 22430 18398 22482 18450
rect 22990 18398 23042 18450
rect 23214 18398 23266 18450
rect 24222 18398 24274 18450
rect 25342 18398 25394 18450
rect 28590 18398 28642 18450
rect 29150 18398 29202 18450
rect 33630 18398 33682 18450
rect 34190 18398 34242 18450
rect 34750 18398 34802 18450
rect 35310 18398 35362 18450
rect 35982 18398 36034 18450
rect 40238 18398 40290 18450
rect 41358 18398 41410 18450
rect 41470 18398 41522 18450
rect 41806 18398 41858 18450
rect 42366 18398 42418 18450
rect 42590 18398 42642 18450
rect 43150 18398 43202 18450
rect 43934 18398 43986 18450
rect 44494 18398 44546 18450
rect 45054 18398 45106 18450
rect 50430 18398 50482 18450
rect 51326 18398 51378 18450
rect 52222 18398 52274 18450
rect 52894 18398 52946 18450
rect 53118 18398 53170 18450
rect 21870 18286 21922 18338
rect 23774 18286 23826 18338
rect 28142 18286 28194 18338
rect 31390 18286 31442 18338
rect 38110 18286 38162 18338
rect 38558 18286 38610 18338
rect 42254 18286 42306 18338
rect 43598 18286 43650 18338
rect 47966 18286 48018 18338
rect 51102 18286 51154 18338
rect 53230 18286 53282 18338
rect 53566 18286 53618 18338
rect 54462 18286 54514 18338
rect 55134 18286 55186 18338
rect 52334 18174 52386 18226
rect 53790 18174 53842 18226
rect 54126 18174 54178 18226
rect 54574 18174 54626 18226
rect 55246 18174 55298 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 51550 17838 51602 17890
rect 51886 17838 51938 17890
rect 52782 17838 52834 17890
rect 22318 17726 22370 17778
rect 35534 17726 35586 17778
rect 38558 17726 38610 17778
rect 40686 17726 40738 17778
rect 42142 17726 42194 17778
rect 44270 17726 44322 17778
rect 47070 17726 47122 17778
rect 50542 17726 50594 17778
rect 54350 17726 54402 17778
rect 56478 17726 56530 17778
rect 17390 17614 17442 17666
rect 17950 17614 18002 17666
rect 18398 17614 18450 17666
rect 18958 17614 19010 17666
rect 19182 17614 19234 17666
rect 19854 17614 19906 17666
rect 21198 17614 21250 17666
rect 21534 17614 21586 17666
rect 21870 17614 21922 17666
rect 23102 17614 23154 17666
rect 30494 17614 30546 17666
rect 30830 17614 30882 17666
rect 31502 17614 31554 17666
rect 32174 17614 32226 17666
rect 35086 17614 35138 17666
rect 37886 17614 37938 17666
rect 41470 17614 41522 17666
rect 44942 17614 44994 17666
rect 46958 17614 47010 17666
rect 47182 17614 47234 17666
rect 50430 17614 50482 17666
rect 50654 17614 50706 17666
rect 50990 17614 51042 17666
rect 51326 17614 51378 17666
rect 52670 17614 52722 17666
rect 53566 17614 53618 17666
rect 57262 17614 57314 17666
rect 17726 17502 17778 17554
rect 22766 17502 22818 17554
rect 31166 17502 31218 17554
rect 53342 17502 53394 17554
rect 57822 17502 57874 17554
rect 58158 17502 58210 17554
rect 17502 17390 17554 17442
rect 18286 17390 18338 17442
rect 18510 17390 18562 17442
rect 19294 17390 19346 17442
rect 19406 17390 19458 17442
rect 21422 17390 21474 17442
rect 28366 17390 28418 17442
rect 30718 17390 30770 17442
rect 31614 17390 31666 17442
rect 31726 17390 31778 17442
rect 35982 17390 36034 17442
rect 46622 17390 46674 17442
rect 47406 17390 47458 17442
rect 53118 17390 53170 17442
rect 53454 17390 53506 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 18286 17054 18338 17106
rect 18734 17054 18786 17106
rect 33182 17054 33234 17106
rect 51886 17054 51938 17106
rect 52110 17054 52162 17106
rect 57486 17054 57538 17106
rect 58270 17054 58322 17106
rect 14702 16942 14754 16994
rect 19070 16942 19122 16994
rect 20638 16942 20690 16994
rect 27582 16942 27634 16994
rect 28142 16942 28194 16994
rect 28702 16942 28754 16994
rect 30382 16942 30434 16994
rect 48974 16942 49026 16994
rect 14030 16830 14082 16882
rect 17614 16830 17666 16882
rect 18398 16830 18450 16882
rect 18734 16830 18786 16882
rect 19630 16830 19682 16882
rect 19854 16830 19906 16882
rect 27694 16830 27746 16882
rect 28254 16830 28306 16882
rect 28926 16830 28978 16882
rect 29374 16830 29426 16882
rect 29710 16830 29762 16882
rect 49310 16830 49362 16882
rect 51438 16830 51490 16882
rect 52670 16830 52722 16882
rect 52894 16830 52946 16882
rect 53566 16830 53618 16882
rect 16830 16718 16882 16770
rect 22766 16718 22818 16770
rect 27918 16718 27970 16770
rect 28814 16718 28866 16770
rect 32510 16718 32562 16770
rect 41022 16718 41074 16770
rect 41470 16718 41522 16770
rect 51214 16718 51266 16770
rect 51998 16718 52050 16770
rect 53342 16718 53394 16770
rect 53790 16718 53842 16770
rect 54014 16718 54066 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 16718 16158 16770 16210
rect 18846 16158 18898 16210
rect 19742 16158 19794 16210
rect 22430 16158 22482 16210
rect 25230 16158 25282 16210
rect 35646 16158 35698 16210
rect 36094 16158 36146 16210
rect 38222 16158 38274 16210
rect 41470 16158 41522 16210
rect 49310 16158 49362 16210
rect 55246 16158 55298 16210
rect 57374 16158 57426 16210
rect 15934 16046 15986 16098
rect 22766 16046 22818 16098
rect 22990 16046 23042 16098
rect 27694 16046 27746 16098
rect 29262 16046 29314 16098
rect 32062 16046 32114 16098
rect 32398 16046 32450 16098
rect 32622 16046 32674 16098
rect 33630 16046 33682 16098
rect 33966 16046 34018 16098
rect 49534 16046 49586 16098
rect 51662 16046 51714 16098
rect 58046 16046 58098 16098
rect 19294 15934 19346 15986
rect 23326 15934 23378 15986
rect 24446 15934 24498 15986
rect 24670 15934 24722 15986
rect 27470 15934 27522 15986
rect 28142 15934 28194 15986
rect 28366 15934 28418 15986
rect 29374 15934 29426 15986
rect 29710 15934 29762 15986
rect 34302 15934 34354 15986
rect 35310 15934 35362 15986
rect 35534 15934 35586 15986
rect 47854 15934 47906 15986
rect 50542 15934 50594 15986
rect 22990 15822 23042 15874
rect 24558 15822 24610 15874
rect 27918 15822 27970 15874
rect 29486 15822 29538 15874
rect 33070 15822 33122 15874
rect 33966 15822 34018 15874
rect 37886 15822 37938 15874
rect 45390 15822 45442 15874
rect 45726 15822 45778 15874
rect 52110 15822 52162 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 21870 15486 21922 15538
rect 29934 15486 29986 15538
rect 33518 15486 33570 15538
rect 38110 15486 38162 15538
rect 47742 15486 47794 15538
rect 52446 15486 52498 15538
rect 58158 15486 58210 15538
rect 24222 15374 24274 15426
rect 27358 15374 27410 15426
rect 35646 15374 35698 15426
rect 39118 15374 39170 15426
rect 45054 15374 45106 15426
rect 49086 15374 49138 15426
rect 49422 15374 49474 15426
rect 50094 15374 50146 15426
rect 50430 15374 50482 15426
rect 23774 15262 23826 15314
rect 26686 15262 26738 15314
rect 31502 15262 31554 15314
rect 34974 15262 35026 15314
rect 38446 15262 38498 15314
rect 39566 15262 39618 15314
rect 39902 15262 39954 15314
rect 40910 15262 40962 15314
rect 41134 15262 41186 15314
rect 41918 15262 41970 15314
rect 45278 15262 45330 15314
rect 45614 15262 45666 15314
rect 46846 15262 46898 15314
rect 47294 15262 47346 15314
rect 48974 15262 49026 15314
rect 50654 15262 50706 15314
rect 51774 15262 51826 15314
rect 51998 15262 52050 15314
rect 52670 15262 52722 15314
rect 22430 15150 22482 15202
rect 23662 15150 23714 15202
rect 29486 15150 29538 15202
rect 31726 15150 31778 15202
rect 37774 15150 37826 15202
rect 38670 15150 38722 15202
rect 39678 15150 39730 15202
rect 42590 15150 42642 15202
rect 44718 15150 44770 15202
rect 45166 15150 45218 15202
rect 46622 15150 46674 15202
rect 47070 15150 47122 15202
rect 49310 15150 49362 15202
rect 50206 15150 50258 15202
rect 51550 15150 51602 15202
rect 52558 15150 52610 15202
rect 22206 15038 22258 15090
rect 32062 15038 32114 15090
rect 41470 15038 41522 15090
rect 51214 15038 51266 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 50542 14702 50594 14754
rect 52670 14702 52722 14754
rect 52782 14702 52834 14754
rect 18286 14590 18338 14642
rect 24334 14590 24386 14642
rect 26462 14590 26514 14642
rect 27582 14590 27634 14642
rect 34638 14590 34690 14642
rect 38334 14590 38386 14642
rect 41470 14590 41522 14642
rect 50766 14590 50818 14642
rect 53678 14590 53730 14642
rect 54014 14590 54066 14642
rect 54462 14590 54514 14642
rect 18510 14478 18562 14530
rect 23550 14478 23602 14530
rect 34974 14478 35026 14530
rect 35422 14478 35474 14530
rect 37550 14478 37602 14530
rect 39790 14478 39842 14530
rect 41694 14478 41746 14530
rect 41918 14478 41970 14530
rect 42590 14478 42642 14530
rect 42814 14478 42866 14530
rect 44718 14478 44770 14530
rect 45054 14478 45106 14530
rect 46846 14478 46898 14530
rect 47182 14478 47234 14530
rect 47854 14478 47906 14530
rect 48078 14478 48130 14530
rect 50206 14478 50258 14530
rect 51102 14478 51154 14530
rect 51214 14478 51266 14530
rect 52110 14478 52162 14530
rect 53566 14478 53618 14530
rect 57262 14478 57314 14530
rect 22654 14366 22706 14418
rect 26798 14366 26850 14418
rect 39006 14366 39058 14418
rect 39566 14366 39618 14418
rect 40910 14366 40962 14418
rect 43038 14366 43090 14418
rect 46622 14366 46674 14418
rect 51774 14366 51826 14418
rect 53342 14366 53394 14418
rect 54126 14366 54178 14418
rect 56590 14366 56642 14418
rect 57822 14366 57874 14418
rect 18846 14254 18898 14306
rect 22094 14254 22146 14306
rect 23214 14254 23266 14306
rect 27134 14254 27186 14306
rect 33742 14254 33794 14306
rect 37214 14254 37266 14306
rect 37886 14254 37938 14306
rect 39230 14254 39282 14306
rect 42702 14254 42754 14306
rect 43710 14254 43762 14306
rect 44942 14254 44994 14306
rect 47070 14254 47122 14306
rect 47518 14254 47570 14306
rect 51550 14254 51602 14306
rect 51886 14254 51938 14306
rect 53118 14254 53170 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 17502 13918 17554 13970
rect 20750 13918 20802 13970
rect 23886 13918 23938 13970
rect 24334 13918 24386 13970
rect 40014 13918 40066 13970
rect 42478 13918 42530 13970
rect 43262 13918 43314 13970
rect 47630 13918 47682 13970
rect 47854 13918 47906 13970
rect 50654 13918 50706 13970
rect 50766 13918 50818 13970
rect 14702 13806 14754 13858
rect 27918 13806 27970 13858
rect 34302 13806 34354 13858
rect 34526 13806 34578 13858
rect 35310 13806 35362 13858
rect 41470 13806 41522 13858
rect 42814 13806 42866 13858
rect 44046 13806 44098 13858
rect 44158 13806 44210 13858
rect 44942 13806 44994 13858
rect 45166 13806 45218 13858
rect 52782 13806 52834 13858
rect 55246 13806 55298 13858
rect 14030 13694 14082 13746
rect 18286 13694 18338 13746
rect 18734 13694 18786 13746
rect 18846 13694 18898 13746
rect 18958 13694 19010 13746
rect 19406 13694 19458 13746
rect 19630 13694 19682 13746
rect 19854 13694 19906 13746
rect 20862 13694 20914 13746
rect 21086 13694 21138 13746
rect 21310 13694 21362 13746
rect 21422 13694 21474 13746
rect 21758 13694 21810 13746
rect 22430 13694 22482 13746
rect 22654 13694 22706 13746
rect 22766 13694 22818 13746
rect 22990 13694 23042 13746
rect 23326 13694 23378 13746
rect 23662 13694 23714 13746
rect 27134 13694 27186 13746
rect 33070 13694 33122 13746
rect 33854 13694 33906 13746
rect 34750 13694 34802 13746
rect 35086 13694 35138 13746
rect 39342 13694 39394 13746
rect 39566 13694 39618 13746
rect 41694 13694 41746 13746
rect 41918 13694 41970 13746
rect 42366 13694 42418 13746
rect 42702 13694 42754 13746
rect 44382 13694 44434 13746
rect 47294 13694 47346 13746
rect 50206 13694 50258 13746
rect 50878 13694 50930 13746
rect 52670 13694 52722 13746
rect 55918 13694 55970 13746
rect 16830 13582 16882 13634
rect 22206 13582 22258 13634
rect 23774 13582 23826 13634
rect 30046 13582 30098 13634
rect 30494 13582 30546 13634
rect 32062 13582 32114 13634
rect 32398 13582 32450 13634
rect 34078 13582 34130 13634
rect 34974 13582 35026 13634
rect 35758 13582 35810 13634
rect 37550 13582 37602 13634
rect 38110 13582 38162 13634
rect 38446 13582 38498 13634
rect 42142 13582 42194 13634
rect 43710 13582 43762 13634
rect 44942 13582 44994 13634
rect 47742 13582 47794 13634
rect 53118 13582 53170 13634
rect 56702 13582 56754 13634
rect 20414 13470 20466 13522
rect 32510 13470 32562 13522
rect 33070 13470 33122 13522
rect 33406 13470 33458 13522
rect 37662 13470 37714 13522
rect 38110 13470 38162 13522
rect 39006 13470 39058 13522
rect 39118 13470 39170 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17838 13134 17890 13186
rect 19966 13134 20018 13186
rect 20526 13134 20578 13186
rect 21310 13134 21362 13186
rect 23550 13134 23602 13186
rect 34526 13134 34578 13186
rect 44830 13134 44882 13186
rect 44942 13134 44994 13186
rect 48190 13134 48242 13186
rect 18734 13022 18786 13074
rect 19182 13022 19234 13074
rect 21422 13022 21474 13074
rect 32398 13022 32450 13074
rect 33070 13022 33122 13074
rect 34638 13022 34690 13074
rect 37102 13022 37154 13074
rect 41022 13022 41074 13074
rect 48078 13022 48130 13074
rect 17950 12910 18002 12962
rect 18398 12910 18450 12962
rect 18622 12910 18674 12962
rect 19854 12910 19906 12962
rect 21646 12910 21698 12962
rect 23326 12910 23378 12962
rect 23774 12910 23826 12962
rect 24110 12910 24162 12962
rect 24446 12910 24498 12962
rect 29486 12910 29538 12962
rect 30270 12910 30322 12962
rect 33294 12910 33346 12962
rect 33630 12910 33682 12962
rect 34862 12910 34914 12962
rect 35198 12910 35250 12962
rect 35646 12910 35698 12962
rect 35870 12910 35922 12962
rect 36318 12910 36370 12962
rect 39678 12910 39730 12962
rect 43710 12910 43762 12962
rect 45726 12910 45778 12962
rect 47182 12910 47234 12962
rect 18846 12798 18898 12850
rect 20414 12798 20466 12850
rect 22094 12798 22146 12850
rect 22430 12798 22482 12850
rect 22542 12798 22594 12850
rect 22766 12798 22818 12850
rect 22990 12798 23042 12850
rect 24782 12798 24834 12850
rect 34974 12798 35026 12850
rect 42030 12798 42082 12850
rect 45502 12798 45554 12850
rect 47518 12798 47570 12850
rect 47854 12798 47906 12850
rect 17838 12686 17890 12738
rect 19294 12686 19346 12738
rect 19406 12686 19458 12738
rect 19966 12686 20018 12738
rect 23438 12686 23490 12738
rect 24334 12686 24386 12738
rect 25230 12686 25282 12738
rect 33966 12686 34018 12738
rect 35534 12686 35586 12738
rect 38782 12686 38834 12738
rect 42366 12686 42418 12738
rect 42814 12686 42866 12738
rect 43374 12686 43426 12738
rect 44046 12686 44098 12738
rect 45278 12686 45330 12738
rect 45614 12686 45666 12738
rect 47406 12686 47458 12738
rect 51102 12686 51154 12738
rect 51438 12686 51490 12738
rect 53006 12686 53058 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 20862 12350 20914 12402
rect 23326 12350 23378 12402
rect 24222 12350 24274 12402
rect 24558 12350 24610 12402
rect 28366 12350 28418 12402
rect 33070 12350 33122 12402
rect 34526 12350 34578 12402
rect 39006 12350 39058 12402
rect 39902 12350 39954 12402
rect 41134 12350 41186 12402
rect 42590 12350 42642 12402
rect 50654 12350 50706 12402
rect 51662 12350 51714 12402
rect 52110 12350 52162 12402
rect 19518 12238 19570 12290
rect 27358 12238 27410 12290
rect 34862 12238 34914 12290
rect 35982 12238 36034 12290
rect 39118 12238 39170 12290
rect 40910 12238 40962 12290
rect 44718 12238 44770 12290
rect 47742 12238 47794 12290
rect 50990 12238 51042 12290
rect 52222 12238 52274 12290
rect 52670 12238 52722 12290
rect 18286 12126 18338 12178
rect 27134 12126 27186 12178
rect 27470 12126 27522 12178
rect 30158 12126 30210 12178
rect 33294 12126 33346 12178
rect 33742 12126 33794 12178
rect 34302 12126 34354 12178
rect 34638 12126 34690 12178
rect 35310 12126 35362 12178
rect 38782 12126 38834 12178
rect 39230 12126 39282 12178
rect 39566 12126 39618 12178
rect 39902 12126 39954 12178
rect 40238 12126 40290 12178
rect 49870 12126 49922 12178
rect 50318 12126 50370 12178
rect 51326 12126 51378 12178
rect 51886 12126 51938 12178
rect 53342 12126 53394 12178
rect 21198 12014 21250 12066
rect 27918 12014 27970 12066
rect 30830 12014 30882 12066
rect 33182 12014 33234 12066
rect 38110 12014 38162 12066
rect 41246 12014 41298 12066
rect 41694 12014 41746 12066
rect 42142 12014 42194 12066
rect 54462 12014 54514 12066
rect 44158 11902 44210 11954
rect 44382 11902 44434 11954
rect 44606 11902 44658 11954
rect 47854 11902 47906 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19630 11566 19682 11618
rect 32062 11566 32114 11618
rect 33070 11566 33122 11618
rect 33406 11566 33458 11618
rect 57262 11566 57314 11618
rect 17278 11454 17330 11506
rect 17726 11454 17778 11506
rect 19518 11454 19570 11506
rect 24670 11454 24722 11506
rect 31838 11454 31890 11506
rect 33070 11454 33122 11506
rect 33966 11454 34018 11506
rect 35086 11454 35138 11506
rect 38334 11454 38386 11506
rect 40238 11454 40290 11506
rect 42366 11454 42418 11506
rect 43038 11454 43090 11506
rect 46734 11454 46786 11506
rect 48862 11454 48914 11506
rect 50094 11454 50146 11506
rect 50654 11454 50706 11506
rect 51662 11454 51714 11506
rect 52670 11454 52722 11506
rect 54798 11454 54850 11506
rect 14478 11342 14530 11394
rect 18734 11342 18786 11394
rect 21534 11342 21586 11394
rect 24334 11342 24386 11394
rect 27582 11342 27634 11394
rect 28254 11342 28306 11394
rect 29262 11342 29314 11394
rect 31614 11342 31666 11394
rect 32286 11342 32338 11394
rect 32622 11342 32674 11394
rect 39454 11342 39506 11394
rect 49646 11342 49698 11394
rect 50990 11342 51042 11394
rect 51886 11342 51938 11394
rect 52110 11342 52162 11394
rect 55582 11342 55634 11394
rect 15150 11230 15202 11282
rect 18958 11230 19010 11282
rect 19294 11230 19346 11282
rect 21310 11230 21362 11282
rect 26798 11230 26850 11282
rect 37886 11230 37938 11282
rect 38670 11230 38722 11282
rect 51326 11230 51378 11282
rect 51550 11230 51602 11282
rect 57374 11230 57426 11282
rect 57822 11230 57874 11282
rect 58158 11230 58210 11282
rect 18846 11118 18898 11170
rect 20190 11118 20242 11170
rect 23998 11118 24050 11170
rect 27918 11118 27970 11170
rect 30718 11118 30770 11170
rect 31502 11118 31554 11170
rect 33518 11118 33570 11170
rect 39006 11118 39058 11170
rect 51102 11118 51154 11170
rect 56030 11118 56082 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 15710 10782 15762 10834
rect 18174 10782 18226 10834
rect 25902 10782 25954 10834
rect 26238 10782 26290 10834
rect 26798 10782 26850 10834
rect 42814 10782 42866 10834
rect 50206 10782 50258 10834
rect 51998 10782 52050 10834
rect 15822 10670 15874 10722
rect 18062 10670 18114 10722
rect 18398 10670 18450 10722
rect 18734 10670 18786 10722
rect 23774 10670 23826 10722
rect 26350 10670 26402 10722
rect 27022 10670 27074 10722
rect 31166 10670 31218 10722
rect 31726 10670 31778 10722
rect 43934 10670 43986 10722
rect 47182 10670 47234 10722
rect 51326 10670 51378 10722
rect 51438 10670 51490 10722
rect 52446 10670 52498 10722
rect 17950 10558 18002 10610
rect 24558 10558 24610 10610
rect 25342 10558 25394 10610
rect 26574 10558 26626 10610
rect 27134 10558 27186 10610
rect 30382 10558 30434 10610
rect 30942 10558 30994 10610
rect 31278 10558 31330 10610
rect 41806 10558 41858 10610
rect 43150 10558 43202 10610
rect 46846 10558 46898 10610
rect 49870 10558 49922 10610
rect 51662 10558 51714 10610
rect 58158 10558 58210 10610
rect 21646 10446 21698 10498
rect 27582 10446 27634 10498
rect 29710 10446 29762 10498
rect 42254 10446 42306 10498
rect 46062 10446 46114 10498
rect 49534 10446 49586 10498
rect 50654 10446 50706 10498
rect 18958 10334 19010 10386
rect 19182 10334 19234 10386
rect 19406 10334 19458 10386
rect 19854 10334 19906 10386
rect 26238 10334 26290 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 17726 9998 17778 10050
rect 18062 9998 18114 10050
rect 19518 9998 19570 10050
rect 32734 9998 32786 10050
rect 17278 9886 17330 9938
rect 20078 9886 20130 9938
rect 22206 9886 22258 9938
rect 30494 9886 30546 9938
rect 32286 9886 32338 9938
rect 35422 9886 35474 9938
rect 42590 9886 42642 9938
rect 52670 9886 52722 9938
rect 14478 9774 14530 9826
rect 18286 9774 18338 9826
rect 18734 9774 18786 9826
rect 18958 9774 19010 9826
rect 19630 9774 19682 9826
rect 21758 9774 21810 9826
rect 24894 9774 24946 9826
rect 25342 9774 25394 9826
rect 27470 9774 27522 9826
rect 28030 9774 28082 9826
rect 31166 9774 31218 9826
rect 31838 9774 31890 9826
rect 33182 9774 33234 9826
rect 33406 9774 33458 9826
rect 33742 9774 33794 9826
rect 35646 9774 35698 9826
rect 35870 9774 35922 9826
rect 36094 9774 36146 9826
rect 37662 9774 37714 9826
rect 41470 9774 41522 9826
rect 43038 9774 43090 9826
rect 43486 9774 43538 9826
rect 43822 9774 43874 9826
rect 50766 9774 50818 9826
rect 51102 9774 51154 9826
rect 51438 9774 51490 9826
rect 51774 9774 51826 9826
rect 51998 9774 52050 9826
rect 55582 9774 55634 9826
rect 15150 9662 15202 9714
rect 19294 9662 19346 9714
rect 23438 9662 23490 9714
rect 25902 9662 25954 9714
rect 28590 9662 28642 9714
rect 29934 9662 29986 9714
rect 30718 9662 30770 9714
rect 31502 9662 31554 9714
rect 32734 9662 32786 9714
rect 32846 9662 32898 9714
rect 34078 9662 34130 9714
rect 34414 9662 34466 9714
rect 36542 9662 36594 9714
rect 37774 9662 37826 9714
rect 39566 9662 39618 9714
rect 40350 9662 40402 9714
rect 44158 9662 44210 9714
rect 50878 9662 50930 9714
rect 51662 9662 51714 9714
rect 54798 9662 54850 9714
rect 18846 9550 18898 9602
rect 21422 9550 21474 9602
rect 27022 9550 27074 9602
rect 27582 9550 27634 9602
rect 30046 9550 30098 9602
rect 30382 9550 30434 9602
rect 30606 9550 30658 9602
rect 33406 9550 33458 9602
rect 50430 9550 50482 9602
rect 56030 9550 56082 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 15710 9214 15762 9266
rect 17502 9214 17554 9266
rect 18734 9214 18786 9266
rect 22094 9214 22146 9266
rect 27582 9214 27634 9266
rect 31390 9214 31442 9266
rect 33294 9214 33346 9266
rect 33854 9214 33906 9266
rect 40238 9214 40290 9266
rect 41918 9214 41970 9266
rect 44270 9214 44322 9266
rect 50206 9214 50258 9266
rect 51326 9214 51378 9266
rect 15822 9102 15874 9154
rect 18846 9102 18898 9154
rect 31054 9102 31106 9154
rect 33518 9102 33570 9154
rect 33630 9102 33682 9154
rect 35534 9102 35586 9154
rect 37102 9102 37154 9154
rect 37326 9102 37378 9154
rect 37662 9102 37714 9154
rect 39230 9102 39282 9154
rect 39566 9102 39618 9154
rect 39902 9102 39954 9154
rect 42142 9102 42194 9154
rect 42814 9102 42866 9154
rect 43150 9102 43202 9154
rect 43486 9102 43538 9154
rect 43822 9102 43874 9154
rect 49982 9102 50034 9154
rect 18958 8990 19010 9042
rect 19294 8990 19346 9042
rect 22430 8990 22482 9042
rect 35086 8990 35138 9042
rect 35310 8990 35362 9042
rect 42366 8990 42418 9042
rect 44606 8990 44658 9042
rect 50430 8990 50482 9042
rect 35422 8878 35474 8930
rect 37550 8878 37602 8930
rect 45390 8878 45442 8930
rect 47518 8878 47570 8930
rect 50318 8878 50370 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 35310 8430 35362 8482
rect 32510 8318 32562 8370
rect 33630 8318 33682 8370
rect 44942 8318 44994 8370
rect 45390 8318 45442 8370
rect 47406 8318 47458 8370
rect 51214 8318 51266 8370
rect 26910 8206 26962 8258
rect 27358 8206 27410 8258
rect 30942 8206 30994 8258
rect 31502 8206 31554 8258
rect 32174 8206 32226 8258
rect 33966 8206 34018 8258
rect 35534 8206 35586 8258
rect 35870 8206 35922 8258
rect 45166 8206 45218 8258
rect 45614 8206 45666 8258
rect 45838 8206 45890 8258
rect 46286 8206 46338 8258
rect 46398 8206 46450 8258
rect 47182 8206 47234 8258
rect 47518 8206 47570 8258
rect 48414 8206 48466 8258
rect 48638 8206 48690 8258
rect 48862 8206 48914 8258
rect 49534 8206 49586 8258
rect 50430 8206 50482 8258
rect 50990 8206 51042 8258
rect 30606 8094 30658 8146
rect 31166 8094 31218 8146
rect 31614 8094 31666 8146
rect 36318 8094 36370 8146
rect 46622 8094 46674 8146
rect 47854 8094 47906 8146
rect 48190 8094 48242 8146
rect 49870 8094 49922 8146
rect 26686 7982 26738 8034
rect 26798 7982 26850 8034
rect 30718 7982 30770 8034
rect 31726 7982 31778 8034
rect 33742 7982 33794 8034
rect 34974 7982 35026 8034
rect 35982 7982 36034 8034
rect 36094 7982 36146 8034
rect 39006 7982 39058 8034
rect 39342 7982 39394 8034
rect 39678 7982 39730 8034
rect 46174 7982 46226 8034
rect 49310 7982 49362 8034
rect 50542 7982 50594 8034
rect 51550 7982 51602 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 19070 7646 19122 7698
rect 24782 7646 24834 7698
rect 31502 7646 31554 7698
rect 36766 7646 36818 7698
rect 38446 7646 38498 7698
rect 40014 7646 40066 7698
rect 41358 7646 41410 7698
rect 41470 7646 41522 7698
rect 42590 7646 42642 7698
rect 42926 7646 42978 7698
rect 43598 7646 43650 7698
rect 45838 7646 45890 7698
rect 49646 7646 49698 7698
rect 49758 7646 49810 7698
rect 18958 7534 19010 7586
rect 19630 7534 19682 7586
rect 26798 7534 26850 7586
rect 29822 7534 29874 7586
rect 33854 7534 33906 7586
rect 35646 7534 35698 7586
rect 36430 7534 36482 7586
rect 39790 7534 39842 7586
rect 40126 7534 40178 7586
rect 43262 7534 43314 7586
rect 43822 7534 43874 7586
rect 50878 7534 50930 7586
rect 51214 7534 51266 7586
rect 18846 7422 18898 7474
rect 19406 7422 19458 7474
rect 19854 7422 19906 7474
rect 20302 7422 20354 7474
rect 23326 7422 23378 7474
rect 24110 7422 24162 7474
rect 24334 7422 24386 7474
rect 26350 7422 26402 7474
rect 26574 7422 26626 7474
rect 27022 7422 27074 7474
rect 27246 7422 27298 7474
rect 30494 7422 30546 7474
rect 33518 7422 33570 7474
rect 33630 7422 33682 7474
rect 34190 7422 34242 7474
rect 34302 7422 34354 7474
rect 34526 7422 34578 7474
rect 35086 7422 35138 7474
rect 35310 7422 35362 7474
rect 35422 7422 35474 7474
rect 36094 7422 36146 7474
rect 37886 7422 37938 7474
rect 38110 7422 38162 7474
rect 38670 7422 38722 7474
rect 39118 7422 39170 7474
rect 40350 7422 40402 7474
rect 40798 7422 40850 7474
rect 41246 7422 41298 7474
rect 44158 7422 44210 7474
rect 44606 7422 44658 7474
rect 49870 7422 49922 7474
rect 50206 7422 50258 7474
rect 50542 7422 50594 7474
rect 50654 7422 50706 7474
rect 51438 7422 51490 7474
rect 19742 7310 19794 7362
rect 21310 7310 21362 7362
rect 23662 7310 23714 7362
rect 27694 7310 27746 7362
rect 31838 7310 31890 7362
rect 38558 7310 38610 7362
rect 43710 7310 43762 7362
rect 44158 7310 44210 7362
rect 44494 7310 44546 7362
rect 51550 7310 51602 7362
rect 52446 7310 52498 7362
rect 20750 7198 20802 7250
rect 21086 7198 21138 7250
rect 22766 7198 22818 7250
rect 23102 7198 23154 7250
rect 23886 7198 23938 7250
rect 25790 7198 25842 7250
rect 26126 7198 26178 7250
rect 35982 7198 36034 7250
rect 37550 7198 37602 7250
rect 52558 7198 52610 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19518 6862 19570 6914
rect 19630 6862 19682 6914
rect 21422 6862 21474 6914
rect 23550 6862 23602 6914
rect 26798 6862 26850 6914
rect 26910 6862 26962 6914
rect 38782 6862 38834 6914
rect 38894 6862 38946 6914
rect 40798 6862 40850 6914
rect 40910 6862 40962 6914
rect 41582 6862 41634 6914
rect 50318 6862 50370 6914
rect 18286 6750 18338 6802
rect 18622 6750 18674 6802
rect 20638 6750 20690 6802
rect 21310 6750 21362 6802
rect 22206 6750 22258 6802
rect 24334 6750 24386 6802
rect 25902 6750 25954 6802
rect 32286 6750 32338 6802
rect 36206 6750 36258 6802
rect 41246 6750 41298 6802
rect 41806 6750 41858 6802
rect 48750 6750 48802 6802
rect 49982 6750 50034 6802
rect 50430 6750 50482 6802
rect 52670 6750 52722 6802
rect 15486 6638 15538 6690
rect 18734 6638 18786 6690
rect 20526 6638 20578 6690
rect 23438 6638 23490 6690
rect 24110 6638 24162 6690
rect 24446 6638 24498 6690
rect 25118 6638 25170 6690
rect 25454 6638 25506 6690
rect 26238 6638 26290 6690
rect 27582 6638 27634 6690
rect 28030 6638 28082 6690
rect 30158 6638 30210 6690
rect 30270 6638 30322 6690
rect 31278 6638 31330 6690
rect 31950 6638 32002 6690
rect 37886 6638 37938 6690
rect 38222 6638 38274 6690
rect 40238 6638 40290 6690
rect 42926 6638 42978 6690
rect 43486 6638 43538 6690
rect 43934 6638 43986 6690
rect 46398 6638 46450 6690
rect 46846 6638 46898 6690
rect 48414 6638 48466 6690
rect 49758 6638 49810 6690
rect 50990 6638 51042 6690
rect 54798 6638 54850 6690
rect 55470 6638 55522 6690
rect 56030 6638 56082 6690
rect 16158 6526 16210 6578
rect 18958 6526 19010 6578
rect 21982 6526 22034 6578
rect 22206 6526 22258 6578
rect 24782 6526 24834 6578
rect 25230 6526 25282 6578
rect 26014 6526 26066 6578
rect 26574 6526 26626 6578
rect 27246 6526 27298 6578
rect 30942 6526 30994 6578
rect 38558 6526 38610 6578
rect 40014 6526 40066 6578
rect 40574 6526 40626 6578
rect 43262 6526 43314 6578
rect 48526 6526 48578 6578
rect 48862 6526 48914 6578
rect 49422 6526 49474 6578
rect 50766 6526 50818 6578
rect 51214 6526 51266 6578
rect 19182 6414 19234 6466
rect 20302 6414 20354 6466
rect 20750 6414 20802 6466
rect 21758 6414 21810 6466
rect 23886 6414 23938 6466
rect 30718 6414 30770 6466
rect 30830 6414 30882 6466
rect 31390 6414 31442 6466
rect 31502 6414 31554 6466
rect 38110 6414 38162 6466
rect 40126 6414 40178 6466
rect 43150 6414 43202 6466
rect 51102 6414 51154 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 17390 6078 17442 6130
rect 23662 6078 23714 6130
rect 23774 6078 23826 6130
rect 31166 6078 31218 6130
rect 32062 6078 32114 6130
rect 32398 6078 32450 6130
rect 46286 6078 46338 6130
rect 46734 6078 46786 6130
rect 21534 5966 21586 6018
rect 31278 5966 31330 6018
rect 33854 5966 33906 6018
rect 35422 5966 35474 6018
rect 43710 5966 43762 6018
rect 45054 5966 45106 6018
rect 46174 5966 46226 6018
rect 46510 5966 46562 6018
rect 46958 5966 47010 6018
rect 47070 5966 47122 6018
rect 47294 5966 47346 6018
rect 17502 5854 17554 5906
rect 19070 5854 19122 5906
rect 19294 5854 19346 5906
rect 21758 5854 21810 5906
rect 21982 5854 22034 5906
rect 23550 5854 23602 5906
rect 24110 5854 24162 5906
rect 30494 5854 30546 5906
rect 30942 5854 30994 5906
rect 31390 5854 31442 5906
rect 44382 5854 44434 5906
rect 45278 5854 45330 5906
rect 45614 5854 45666 5906
rect 18398 5742 18450 5794
rect 21646 5742 21698 5794
rect 27582 5742 27634 5794
rect 29710 5742 29762 5794
rect 41246 5742 41298 5794
rect 41582 5742 41634 5794
rect 45166 5742 45218 5794
rect 47518 5742 47570 5794
rect 18734 5630 18786 5682
rect 33742 5630 33794 5682
rect 35534 5630 35586 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 20190 5182 20242 5234
rect 21422 5182 21474 5234
rect 23214 5182 23266 5234
rect 25902 5182 25954 5234
rect 31614 5182 31666 5234
rect 32062 5182 32114 5234
rect 33518 5182 33570 5234
rect 35646 5182 35698 5234
rect 36990 5182 37042 5234
rect 40350 5182 40402 5234
rect 40686 5182 40738 5234
rect 44046 5182 44098 5234
rect 44942 5182 44994 5234
rect 45502 5182 45554 5234
rect 47742 5182 47794 5234
rect 49870 5182 49922 5234
rect 51214 5182 51266 5234
rect 30718 5070 30770 5122
rect 30830 5070 30882 5122
rect 31054 5070 31106 5122
rect 31166 5070 31218 5122
rect 32734 5070 32786 5122
rect 39118 5070 39170 5122
rect 39902 5070 39954 5122
rect 45838 5070 45890 5122
rect 46510 5070 46562 5122
rect 47070 5070 47122 5122
rect 50318 5070 50370 5122
rect 20078 4846 20130 4898
rect 23102 4846 23154 4898
rect 26014 4846 26066 4898
rect 40798 4846 40850 4898
rect 45950 4846 46002 4898
rect 46062 4846 46114 4898
rect 51326 4846 51378 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 28590 4510 28642 4562
rect 33182 4510 33234 4562
rect 37662 4510 37714 4562
rect 38222 4510 38274 4562
rect 48750 4510 48802 4562
rect 53902 4510 53954 4562
rect 19070 4398 19122 4450
rect 22318 4398 22370 4450
rect 26014 4398 26066 4450
rect 31502 4398 31554 4450
rect 36430 4398 36482 4450
rect 38110 4398 38162 4450
rect 41694 4398 41746 4450
rect 44942 4398 44994 4450
rect 48862 4398 48914 4450
rect 52670 4398 52722 4450
rect 18398 4286 18450 4338
rect 21534 4286 21586 4338
rect 25342 4286 25394 4338
rect 32286 4286 32338 4338
rect 37214 4286 37266 4338
rect 40910 4286 40962 4338
rect 44158 4286 44210 4338
rect 53342 4286 53394 4338
rect 57598 4286 57650 4338
rect 58158 4286 58210 4338
rect 21198 4174 21250 4226
rect 24446 4174 24498 4226
rect 28142 4174 28194 4226
rect 29374 4174 29426 4226
rect 34302 4174 34354 4226
rect 43822 4174 43874 4226
rect 47070 4174 47122 4226
rect 50542 4174 50594 4226
rect 57374 4174 57426 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 21534 3614 21586 3666
rect 43934 3614 43986 3666
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 2688 69200 2800 70000
rect 4704 69200 4816 70000
rect 6720 69200 6832 70000
rect 8736 69200 8848 70000
rect 10752 69200 10864 70000
rect 12768 69200 12880 70000
rect 14784 69200 14896 70000
rect 16800 69200 16912 70000
rect 18816 69200 18928 70000
rect 20832 69200 20944 70000
rect 22848 69200 22960 70000
rect 24864 69200 24976 70000
rect 26880 69200 26992 70000
rect 28896 69200 29008 70000
rect 30912 69200 31024 70000
rect 32928 69200 33040 70000
rect 34944 69200 35056 70000
rect 36960 69200 37072 70000
rect 38976 69200 39088 70000
rect 40992 69200 41104 70000
rect 43008 69200 43120 70000
rect 45024 69200 45136 70000
rect 47040 69200 47152 70000
rect 49056 69200 49168 70000
rect 51072 69200 51184 70000
rect 53088 69200 53200 70000
rect 55104 69200 55216 70000
rect 57120 69200 57232 70000
rect 2716 67228 2772 69200
rect 2716 67172 2996 67228
rect 2940 66162 2996 67172
rect 4732 66836 4788 69200
rect 6748 67228 6804 69200
rect 6748 67172 7028 67228
rect 4732 66770 4788 66780
rect 5516 66836 5572 66846
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 2940 66110 2942 66162
rect 2994 66110 2996 66162
rect 2940 66098 2996 66110
rect 5516 66162 5572 66780
rect 5516 66110 5518 66162
rect 5570 66110 5572 66162
rect 5516 66098 5572 66110
rect 6972 66162 7028 67172
rect 8764 66834 8820 69200
rect 10780 67228 10836 69200
rect 12796 67228 12852 69200
rect 14812 67228 14868 69200
rect 16828 67228 16884 69200
rect 10780 67172 11060 67228
rect 12796 67172 13188 67228
rect 14812 67172 15092 67228
rect 16828 67172 17108 67228
rect 8764 66782 8766 66834
rect 8818 66782 8820 66834
rect 8764 66770 8820 66782
rect 9324 66834 9380 66846
rect 9324 66782 9326 66834
rect 9378 66782 9380 66834
rect 6972 66110 6974 66162
rect 7026 66110 7028 66162
rect 6972 66098 7028 66110
rect 9324 66162 9380 66782
rect 9324 66110 9326 66162
rect 9378 66110 9380 66162
rect 9324 66098 9380 66110
rect 11004 66162 11060 67172
rect 11004 66110 11006 66162
rect 11058 66110 11060 66162
rect 11004 66098 11060 66110
rect 13132 66162 13188 67172
rect 13132 66110 13134 66162
rect 13186 66110 13188 66162
rect 13132 66098 13188 66110
rect 15036 66162 15092 67172
rect 15036 66110 15038 66162
rect 15090 66110 15092 66162
rect 15036 66098 15092 66110
rect 17052 66162 17108 67172
rect 18844 66386 18900 69200
rect 20860 67228 20916 69200
rect 20860 67172 21140 67228
rect 18844 66334 18846 66386
rect 18898 66334 18900 66386
rect 18844 66322 18900 66334
rect 17612 66276 17668 66286
rect 17052 66110 17054 66162
rect 17106 66110 17108 66162
rect 17052 66098 17108 66110
rect 17388 66274 17668 66276
rect 17388 66222 17614 66274
rect 17666 66222 17668 66274
rect 17388 66220 17668 66222
rect 8876 65378 8932 65390
rect 8876 65326 8878 65378
rect 8930 65326 8932 65378
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 8540 64818 8596 64830
rect 8540 64766 8542 64818
rect 8594 64766 8596 64818
rect 5740 64708 5796 64718
rect 5796 64652 5908 64708
rect 5740 64614 5796 64652
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 2828 60786 2884 60798
rect 2828 60734 2830 60786
rect 2882 60734 2884 60786
rect 1820 59108 1876 59118
rect 1708 59106 1876 59108
rect 1708 59054 1822 59106
rect 1874 59054 1876 59106
rect 1708 59052 1876 59054
rect 1708 58324 1764 59052
rect 1820 59042 1876 59052
rect 1708 58230 1764 58268
rect 1820 58660 1876 58670
rect 1820 57650 1876 58604
rect 2828 58660 2884 60734
rect 3500 60674 3556 60686
rect 3500 60622 3502 60674
rect 3554 60622 3556 60674
rect 3500 59444 3556 60622
rect 5628 60676 5684 60686
rect 5628 60582 5684 60620
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 3500 59378 3556 59388
rect 5852 60114 5908 64652
rect 6412 64596 6468 64606
rect 6412 64594 6692 64596
rect 6412 64542 6414 64594
rect 6466 64542 6692 64594
rect 6412 64540 6692 64542
rect 6412 64530 6468 64540
rect 6636 63250 6692 64540
rect 8540 64034 8596 64766
rect 8876 64708 8932 65326
rect 12460 65380 12516 65390
rect 12460 65378 12628 65380
rect 12460 65326 12462 65378
rect 12514 65326 12628 65378
rect 12460 65324 12628 65326
rect 12460 65314 12516 65324
rect 12124 64818 12180 64830
rect 12124 64766 12126 64818
rect 12178 64766 12180 64818
rect 8876 64642 8932 64652
rect 9324 64708 9380 64718
rect 9324 64614 9380 64652
rect 8540 63982 8542 64034
rect 8594 63982 8596 64034
rect 8540 63970 8596 63982
rect 9996 64594 10052 64606
rect 9996 64542 9998 64594
rect 10050 64542 10052 64594
rect 6636 63198 6638 63250
rect 6690 63198 6692 63250
rect 6636 63186 6692 63198
rect 8428 63698 8484 63710
rect 8428 63646 8430 63698
rect 8482 63646 8484 63698
rect 6748 63138 6804 63150
rect 6748 63086 6750 63138
rect 6802 63086 6804 63138
rect 6524 63028 6580 63038
rect 6524 62934 6580 62972
rect 6748 62356 6804 63086
rect 7868 63138 7924 63150
rect 7868 63086 7870 63138
rect 7922 63086 7924 63138
rect 7084 63028 7140 63038
rect 7308 63028 7364 63038
rect 7084 63026 7252 63028
rect 7084 62974 7086 63026
rect 7138 62974 7252 63026
rect 7084 62972 7252 62974
rect 7084 62962 7140 62972
rect 7196 62578 7252 62972
rect 7196 62526 7198 62578
rect 7250 62526 7252 62578
rect 7196 62514 7252 62526
rect 7308 62578 7364 62972
rect 7644 63028 7700 63038
rect 7644 62934 7700 62972
rect 7308 62526 7310 62578
rect 7362 62526 7364 62578
rect 7308 62514 7364 62526
rect 6748 61684 6804 62300
rect 6860 62466 6916 62478
rect 6860 62414 6862 62466
rect 6914 62414 6916 62466
rect 6860 61796 6916 62414
rect 7084 62356 7140 62366
rect 7084 62262 7140 62300
rect 7868 62354 7924 63086
rect 8092 63140 8148 63150
rect 8428 63140 8484 63646
rect 9996 63364 10052 64542
rect 11788 64596 11844 64606
rect 11452 64036 11508 64046
rect 11452 63942 11508 63980
rect 11788 63922 11844 64540
rect 12124 64036 12180 64766
rect 12572 64708 12628 65324
rect 17388 65378 17444 66220
rect 17612 66210 17668 66220
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 20188 65492 20244 65502
rect 17388 65326 17390 65378
rect 17442 65326 17444 65378
rect 17388 65314 17444 65326
rect 17612 65380 17668 65390
rect 11788 63870 11790 63922
rect 11842 63870 11844 63922
rect 11788 63858 11844 63870
rect 11900 63980 12124 64036
rect 9996 63298 10052 63308
rect 11900 63250 11956 63980
rect 12124 63970 12180 63980
rect 12236 64484 12292 64494
rect 12012 63364 12068 63374
rect 12236 63364 12292 64428
rect 12460 63922 12516 63934
rect 12460 63870 12462 63922
rect 12514 63870 12516 63922
rect 12012 63362 12292 63364
rect 12012 63310 12014 63362
rect 12066 63310 12292 63362
rect 12012 63308 12292 63310
rect 12348 63364 12404 63374
rect 12012 63298 12068 63308
rect 12348 63270 12404 63308
rect 11900 63198 11902 63250
rect 11954 63198 11956 63250
rect 11900 63186 11956 63198
rect 8092 63138 8484 63140
rect 8092 63086 8094 63138
rect 8146 63086 8484 63138
rect 8092 63084 8484 63086
rect 12460 63140 12516 63870
rect 12572 63924 12628 64652
rect 13468 64706 13524 64718
rect 13468 64654 13470 64706
rect 13522 64654 13524 64706
rect 12684 64596 12740 64606
rect 12684 64502 12740 64540
rect 12796 64484 12852 64494
rect 13020 64484 13076 64494
rect 12796 64390 12852 64428
rect 12908 64482 13076 64484
rect 12908 64430 13022 64482
rect 13074 64430 13076 64482
rect 12908 64428 13076 64430
rect 12796 64148 12852 64158
rect 12572 63858 12628 63868
rect 12684 64146 12852 64148
rect 12684 64094 12798 64146
rect 12850 64094 12852 64146
rect 12684 64092 12852 64094
rect 12684 63362 12740 64092
rect 12796 64082 12852 64092
rect 12684 63310 12686 63362
rect 12738 63310 12740 63362
rect 12684 63298 12740 63310
rect 12460 63084 12628 63140
rect 7980 62580 8036 62590
rect 8092 62580 8148 63084
rect 12460 62916 12516 62926
rect 7980 62578 8148 62580
rect 7980 62526 7982 62578
rect 8034 62526 8148 62578
rect 7980 62524 8148 62526
rect 7980 62514 8036 62524
rect 7868 62302 7870 62354
rect 7922 62302 7924 62354
rect 7868 62244 7924 62302
rect 8092 62356 8148 62524
rect 12236 62860 12460 62916
rect 8540 62468 8596 62478
rect 8540 62374 8596 62412
rect 10892 62468 10948 62478
rect 10892 62374 10948 62412
rect 8092 62290 8148 62300
rect 8204 62356 8260 62366
rect 8428 62356 8484 62366
rect 8204 62354 8484 62356
rect 8204 62302 8206 62354
rect 8258 62302 8430 62354
rect 8482 62302 8484 62354
rect 8204 62300 8484 62302
rect 8204 62290 8260 62300
rect 8428 62290 8484 62300
rect 8764 62356 8820 62366
rect 9436 62356 9492 62366
rect 8764 62354 9492 62356
rect 8764 62302 8766 62354
rect 8818 62302 9438 62354
rect 9490 62302 9492 62354
rect 8764 62300 9492 62302
rect 8764 62290 8820 62300
rect 9436 62290 9492 62300
rect 10220 62356 10276 62366
rect 10220 62262 10276 62300
rect 7868 62178 7924 62188
rect 10556 62244 10612 62254
rect 6860 61740 7588 61796
rect 7532 61684 7588 61740
rect 6748 61628 7028 61684
rect 6412 61460 6468 61470
rect 6748 61460 6804 61470
rect 6412 61458 6804 61460
rect 6412 61406 6414 61458
rect 6466 61406 6750 61458
rect 6802 61406 6804 61458
rect 6412 61404 6804 61406
rect 6412 61394 6468 61404
rect 6188 61348 6244 61358
rect 6188 60900 6244 61292
rect 6300 61346 6356 61358
rect 6300 61294 6302 61346
rect 6354 61294 6356 61346
rect 6300 61124 6356 61294
rect 6300 61068 6580 61124
rect 6300 60900 6356 60910
rect 6188 60898 6356 60900
rect 6188 60846 6302 60898
rect 6354 60846 6356 60898
rect 6188 60844 6356 60846
rect 6300 60676 6356 60844
rect 6300 60610 6356 60620
rect 5852 60062 5854 60114
rect 5906 60062 5908 60114
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4844 58772 4900 58782
rect 2828 58594 2884 58604
rect 4172 58604 4788 58660
rect 1820 57598 1822 57650
rect 1874 57598 1876 57650
rect 1820 54514 1876 57598
rect 1820 54462 1822 54514
rect 1874 54462 1876 54514
rect 1820 54450 1876 54462
rect 2268 58434 2324 58446
rect 2268 58382 2270 58434
rect 2322 58382 2324 58434
rect 1820 50594 1876 50606
rect 1820 50542 1822 50594
rect 1874 50542 1876 50594
rect 1820 47572 1876 50542
rect 1820 47458 1876 47516
rect 1820 47406 1822 47458
rect 1874 47406 1876 47458
rect 1820 47394 1876 47406
rect 2268 43708 2324 58382
rect 4172 58434 4228 58604
rect 4172 58382 4174 58434
rect 4226 58382 4228 58434
rect 4172 58370 4228 58382
rect 4284 58434 4340 58446
rect 4284 58382 4286 58434
rect 4338 58382 4340 58434
rect 3836 58324 3892 58334
rect 3836 58230 3892 58268
rect 4060 58324 4116 58334
rect 2492 58212 2548 58222
rect 2492 57762 2548 58156
rect 3948 58212 4004 58222
rect 3948 58118 4004 58156
rect 4060 58100 4116 58268
rect 4060 58044 4228 58100
rect 2492 57710 2494 57762
rect 2546 57710 2548 57762
rect 2492 57698 2548 57710
rect 4172 56756 4228 58044
rect 4284 56980 4340 58382
rect 4620 57540 4676 57550
rect 4620 57446 4676 57484
rect 4732 57428 4788 58604
rect 4844 58546 4900 58716
rect 5852 58772 5908 60062
rect 6524 60002 6580 61068
rect 6524 59950 6526 60002
rect 6578 59950 6580 60002
rect 6524 59938 6580 59950
rect 6748 60786 6804 61404
rect 6860 61348 6916 61358
rect 6860 61254 6916 61292
rect 6748 60734 6750 60786
rect 6802 60734 6804 60786
rect 5852 58706 5908 58716
rect 6636 58772 6692 58782
rect 4844 58494 4846 58546
rect 4898 58494 4900 58546
rect 4844 58482 4900 58494
rect 5628 58436 5684 58446
rect 5628 58434 5908 58436
rect 5628 58382 5630 58434
rect 5682 58382 5908 58434
rect 5628 58380 5908 58382
rect 5628 58370 5684 58380
rect 4956 58324 5012 58334
rect 4956 57762 5012 58268
rect 5740 58210 5796 58222
rect 5740 58158 5742 58210
rect 5794 58158 5796 58210
rect 5740 57764 5796 58158
rect 4956 57710 4958 57762
rect 5010 57710 5012 57762
rect 4956 57698 5012 57710
rect 5628 57708 5796 57764
rect 5628 57650 5684 57708
rect 5628 57598 5630 57650
rect 5682 57598 5684 57650
rect 5628 57540 5684 57598
rect 4732 57372 4900 57428
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4508 56980 4564 56990
rect 4844 56980 4900 57372
rect 4284 56978 4564 56980
rect 4284 56926 4510 56978
rect 4562 56926 4564 56978
rect 4284 56924 4564 56926
rect 4508 56914 4564 56924
rect 4620 56924 4844 56980
rect 4620 56866 4676 56924
rect 4620 56814 4622 56866
rect 4674 56814 4676 56866
rect 4620 56802 4676 56814
rect 4396 56756 4452 56766
rect 4172 56754 4452 56756
rect 4172 56702 4398 56754
rect 4450 56702 4452 56754
rect 4172 56700 4452 56702
rect 4396 56690 4452 56700
rect 4732 56420 4788 56924
rect 4844 56886 4900 56924
rect 5516 56980 5572 56990
rect 5068 56866 5124 56878
rect 5068 56814 5070 56866
rect 5122 56814 5124 56866
rect 4732 56364 4900 56420
rect 4620 55972 4676 55982
rect 4284 55916 4620 55972
rect 4284 55468 4340 55916
rect 4620 55878 4676 55916
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4844 55522 4900 56364
rect 5068 55972 5124 56814
rect 5292 56868 5348 56878
rect 5180 55972 5236 55982
rect 5068 55916 5180 55972
rect 5180 55878 5236 55916
rect 4844 55470 4846 55522
rect 4898 55470 4900 55522
rect 4284 55412 4564 55468
rect 4844 55458 4900 55470
rect 2940 55300 2996 55310
rect 3500 55300 3556 55310
rect 3948 55300 4004 55310
rect 2940 55298 3220 55300
rect 2940 55246 2942 55298
rect 2994 55246 3220 55298
rect 2940 55244 3220 55246
rect 2940 55234 2996 55244
rect 3052 55074 3108 55086
rect 3052 55022 3054 55074
rect 3106 55022 3108 55074
rect 3052 54740 3108 55022
rect 2492 54684 3108 54740
rect 3164 55076 3220 55244
rect 3500 55298 4004 55300
rect 3500 55246 3502 55298
rect 3554 55246 3950 55298
rect 4002 55246 4004 55298
rect 3500 55244 4004 55246
rect 3500 55234 3556 55244
rect 3948 55234 4004 55244
rect 4508 55298 4564 55412
rect 4508 55246 4510 55298
rect 4562 55246 4564 55298
rect 4508 55234 4564 55246
rect 2492 54626 2548 54684
rect 3164 54628 3220 55020
rect 2492 54574 2494 54626
rect 2546 54574 2548 54626
rect 2492 54562 2548 54574
rect 2940 54572 3220 54628
rect 3276 55186 3332 55198
rect 3276 55134 3278 55186
rect 3330 55134 3332 55186
rect 3276 54628 3332 55134
rect 4956 55188 5012 55198
rect 4956 55186 5124 55188
rect 4956 55134 4958 55186
rect 5010 55134 5124 55186
rect 4956 55132 5124 55134
rect 4956 55122 5012 55132
rect 3836 55076 3892 55086
rect 3836 54982 3892 55020
rect 4060 55074 4116 55086
rect 4060 55022 4062 55074
rect 4114 55022 4116 55074
rect 2940 53842 2996 54572
rect 3276 54562 3332 54572
rect 4060 54628 4116 55022
rect 4060 54562 4116 54572
rect 4844 55074 4900 55086
rect 4844 55022 4846 55074
rect 4898 55022 4900 55074
rect 4620 54516 4676 54526
rect 4620 54404 4676 54460
rect 4284 54402 4676 54404
rect 4284 54350 4622 54402
rect 4674 54350 4676 54402
rect 4284 54348 4676 54350
rect 2940 53790 2942 53842
rect 2994 53790 2996 53842
rect 2940 53778 2996 53790
rect 3388 53956 3444 53966
rect 3388 53730 3444 53900
rect 4284 53956 4340 54348
rect 4620 54338 4676 54348
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4844 53956 4900 55022
rect 5068 54738 5124 55132
rect 5068 54686 5070 54738
rect 5122 54686 5124 54738
rect 5068 54674 5124 54686
rect 4340 53900 4452 53956
rect 4284 53862 4340 53900
rect 3388 53678 3390 53730
rect 3442 53678 3444 53730
rect 3388 53666 3444 53678
rect 3836 53730 3892 53742
rect 3836 53678 3838 53730
rect 3890 53678 3892 53730
rect 3836 53620 3892 53678
rect 4284 53620 4340 53630
rect 3836 53618 4340 53620
rect 3836 53566 4286 53618
rect 4338 53566 4340 53618
rect 3836 53564 4340 53566
rect 4284 53060 4340 53564
rect 4396 53618 4452 53900
rect 4620 53900 4900 53956
rect 4956 54514 5012 54526
rect 4956 54462 4958 54514
rect 5010 54462 5012 54514
rect 4620 53730 4676 53900
rect 4620 53678 4622 53730
rect 4674 53678 4676 53730
rect 4620 53666 4676 53678
rect 4396 53566 4398 53618
rect 4450 53566 4452 53618
rect 4396 53554 4452 53566
rect 4284 52994 4340 53004
rect 4956 53060 5012 54462
rect 5180 54516 5236 54526
rect 5180 54422 5236 54460
rect 5292 54180 5348 56812
rect 5516 56866 5572 56924
rect 5516 56814 5518 56866
rect 5570 56814 5572 56866
rect 5516 56802 5572 56814
rect 5628 56868 5684 57484
rect 5852 57538 5908 58380
rect 5964 58212 6020 58222
rect 5964 58210 6356 58212
rect 5964 58158 5966 58210
rect 6018 58158 6356 58210
rect 5964 58156 6356 58158
rect 5964 58146 6020 58156
rect 6300 57650 6356 58156
rect 6300 57598 6302 57650
rect 6354 57598 6356 57650
rect 6300 57586 6356 57598
rect 5852 57486 5854 57538
rect 5906 57486 5908 57538
rect 5852 57092 5908 57486
rect 6524 57428 6580 57438
rect 5852 57026 5908 57036
rect 6076 57426 6580 57428
rect 6076 57374 6526 57426
rect 6578 57374 6580 57426
rect 6076 57372 6580 57374
rect 6076 56978 6132 57372
rect 6524 57362 6580 57372
rect 6076 56926 6078 56978
rect 6130 56926 6132 56978
rect 6076 56914 6132 56926
rect 6188 57092 6244 57102
rect 5964 56868 6020 56878
rect 5628 56866 6020 56868
rect 5628 56814 5966 56866
rect 6018 56814 6020 56866
rect 5628 56812 6020 56814
rect 5964 56802 6020 56812
rect 6188 56642 6244 57036
rect 6636 56868 6692 58716
rect 6748 57652 6804 60734
rect 6972 60226 7028 61628
rect 7532 61682 7700 61684
rect 7532 61630 7534 61682
rect 7586 61630 7700 61682
rect 7532 61628 7700 61630
rect 7532 61618 7588 61628
rect 7084 61348 7140 61358
rect 7084 61346 7476 61348
rect 7084 61294 7086 61346
rect 7138 61294 7476 61346
rect 7084 61292 7476 61294
rect 7084 61282 7140 61292
rect 6972 60174 6974 60226
rect 7026 60174 7028 60226
rect 6972 60162 7028 60174
rect 7084 60002 7140 60014
rect 7084 59950 7086 60002
rect 7138 59950 7140 60002
rect 7084 59780 7140 59950
rect 7420 60002 7476 61292
rect 7420 59950 7422 60002
rect 7474 59950 7476 60002
rect 7420 59938 7476 59950
rect 7532 60786 7588 60798
rect 7532 60734 7534 60786
rect 7586 60734 7588 60786
rect 7532 59780 7588 60734
rect 6860 59724 7588 59780
rect 6860 57874 6916 59724
rect 7644 59668 7700 61628
rect 6860 57822 6862 57874
rect 6914 57822 6916 57874
rect 6860 57810 6916 57822
rect 7196 59612 7700 59668
rect 7868 61010 7924 61022
rect 7868 60958 7870 61010
rect 7922 60958 7924 61010
rect 6748 57596 6916 57652
rect 6748 56868 6804 56878
rect 6636 56812 6748 56868
rect 6748 56774 6804 56812
rect 6860 56756 6916 57596
rect 6860 56690 6916 56700
rect 6188 56590 6190 56642
rect 6242 56590 6244 56642
rect 6188 55524 6244 56590
rect 6188 55458 6244 55468
rect 6636 55972 6692 55982
rect 6636 55468 6692 55916
rect 7196 55468 7252 59612
rect 7644 59444 7700 59454
rect 7644 59350 7700 59388
rect 7532 59332 7588 59342
rect 7532 59238 7588 59276
rect 7756 59332 7812 59342
rect 7868 59332 7924 60958
rect 10220 60788 10276 60798
rect 9100 60116 9156 60126
rect 9100 60022 9156 60060
rect 8428 60004 8484 60014
rect 8428 59910 8484 59948
rect 8652 60004 8708 60014
rect 7756 59330 7924 59332
rect 7756 59278 7758 59330
rect 7810 59278 7924 59330
rect 7756 59276 7924 59278
rect 8204 59332 8260 59342
rect 7756 59266 7812 59276
rect 8204 59238 8260 59276
rect 7980 57708 8260 57764
rect 7980 57650 8036 57708
rect 7980 57598 7982 57650
rect 8034 57598 8036 57650
rect 7980 57586 8036 57598
rect 8092 57538 8148 57550
rect 8092 57486 8094 57538
rect 8146 57486 8148 57538
rect 8092 57204 8148 57486
rect 7420 57148 8148 57204
rect 7420 56978 7476 57148
rect 7420 56926 7422 56978
rect 7474 56926 7476 56978
rect 7420 56914 7476 56926
rect 8204 56308 8260 57708
rect 8316 57652 8372 57662
rect 8428 57652 8484 57662
rect 8316 57650 8428 57652
rect 8316 57598 8318 57650
rect 8370 57598 8428 57650
rect 8316 57596 8428 57598
rect 8316 57586 8372 57596
rect 8204 56242 8260 56252
rect 8316 56196 8372 56206
rect 8316 56102 8372 56140
rect 8428 56084 8484 57596
rect 8540 57650 8596 57662
rect 8540 57598 8542 57650
rect 8594 57598 8596 57650
rect 8540 56308 8596 57598
rect 8652 56868 8708 59948
rect 10220 58548 10276 60732
rect 10556 60228 10612 62188
rect 12236 61684 12292 62860
rect 12460 62822 12516 62860
rect 12572 62132 12628 63084
rect 12908 62354 12964 64428
rect 13020 64418 13076 64428
rect 13468 64484 13524 64654
rect 13804 64596 13860 64606
rect 13468 64418 13524 64428
rect 13692 64482 13748 64494
rect 13692 64430 13694 64482
rect 13746 64430 13748 64482
rect 13580 63924 13636 63934
rect 13580 63830 13636 63868
rect 13692 63364 13748 64430
rect 13804 63476 13860 64540
rect 17612 64146 17668 65324
rect 19516 65380 19572 65390
rect 19516 65286 19572 65324
rect 17948 64708 18004 64718
rect 17948 64614 18004 64652
rect 20188 64708 20244 65436
rect 20860 65492 20916 65502
rect 20860 65378 20916 65436
rect 20860 65326 20862 65378
rect 20914 65326 20916 65378
rect 18620 64596 18676 64606
rect 18620 64594 19684 64596
rect 18620 64542 18622 64594
rect 18674 64542 19684 64594
rect 18620 64540 19684 64542
rect 18620 64530 18676 64540
rect 17612 64094 17614 64146
rect 17666 64094 17668 64146
rect 17612 64082 17668 64094
rect 16716 64036 16772 64046
rect 14252 63812 14308 63822
rect 14252 63810 14980 63812
rect 14252 63758 14254 63810
rect 14306 63758 14980 63810
rect 14252 63756 14980 63758
rect 14252 63746 14308 63756
rect 13804 63420 14084 63476
rect 13692 63308 13860 63364
rect 13692 62916 13748 62926
rect 12908 62302 12910 62354
rect 12962 62302 12964 62354
rect 12908 62290 12964 62302
rect 13132 62466 13188 62478
rect 13132 62414 13134 62466
rect 13186 62414 13188 62466
rect 13132 62132 13188 62414
rect 13692 62356 13748 62860
rect 13692 62290 13748 62300
rect 13804 62354 13860 63308
rect 13916 63140 13972 63150
rect 13916 62578 13972 63084
rect 13916 62526 13918 62578
rect 13970 62526 13972 62578
rect 13916 62514 13972 62526
rect 13804 62302 13806 62354
rect 13858 62302 13860 62354
rect 13804 62290 13860 62302
rect 14028 62132 14084 63420
rect 14812 63026 14868 63038
rect 14812 62974 14814 63026
rect 14866 62974 14868 63026
rect 14812 62466 14868 62974
rect 14924 62578 14980 63756
rect 16380 63810 16436 63822
rect 16380 63758 16382 63810
rect 16434 63758 16436 63810
rect 15484 63140 15540 63150
rect 15484 63046 15540 63084
rect 16268 63138 16324 63150
rect 16268 63086 16270 63138
rect 16322 63086 16324 63138
rect 14924 62526 14926 62578
rect 14978 62526 14980 62578
rect 14924 62514 14980 62526
rect 16268 62916 16324 63086
rect 14812 62414 14814 62466
rect 14866 62414 14868 62466
rect 14812 62402 14868 62414
rect 15148 62356 15204 62366
rect 16268 62356 16324 62860
rect 16380 63028 16436 63758
rect 16380 62580 16436 62972
rect 16492 62580 16548 62590
rect 16380 62578 16548 62580
rect 16380 62526 16494 62578
rect 16546 62526 16548 62578
rect 16380 62524 16548 62526
rect 16492 62514 16548 62524
rect 16716 62578 16772 63980
rect 17724 64036 17780 64046
rect 17724 63942 17780 63980
rect 16828 63924 16884 63934
rect 16828 63830 16884 63868
rect 17276 63922 17332 63934
rect 17276 63870 17278 63922
rect 17330 63870 17332 63922
rect 17276 63140 17332 63870
rect 17836 63922 17892 63934
rect 17836 63870 17838 63922
rect 17890 63870 17892 63922
rect 17836 63476 17892 63870
rect 17500 63420 17892 63476
rect 17500 63250 17556 63420
rect 19628 63362 19684 64540
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 20188 63922 20244 64652
rect 20748 64818 20804 64830
rect 20748 64766 20750 64818
rect 20802 64766 20804 64818
rect 20748 64036 20804 64766
rect 20860 64484 20916 65326
rect 20860 64418 20916 64428
rect 20748 63980 21028 64036
rect 20188 63870 20190 63922
rect 20242 63870 20244 63922
rect 20188 63858 20244 63870
rect 19628 63310 19630 63362
rect 19682 63310 19684 63362
rect 19628 63298 19684 63310
rect 20860 63810 20916 63822
rect 20860 63758 20862 63810
rect 20914 63758 20916 63810
rect 17500 63198 17502 63250
rect 17554 63198 17556 63250
rect 17500 63186 17556 63198
rect 19628 63140 19684 63150
rect 17276 63074 17332 63084
rect 19404 63138 19684 63140
rect 19404 63086 19630 63138
rect 19682 63086 19684 63138
rect 19404 63084 19684 63086
rect 17612 63028 17668 63038
rect 17612 62934 17668 62972
rect 16716 62526 16718 62578
rect 16770 62526 16772 62578
rect 16716 62514 16772 62526
rect 17388 62916 17444 62926
rect 16380 62356 16436 62366
rect 16268 62354 16436 62356
rect 16268 62302 16382 62354
rect 16434 62302 16436 62354
rect 16268 62300 16436 62302
rect 15148 62244 15204 62300
rect 15596 62244 15652 62254
rect 15148 62242 15652 62244
rect 15148 62190 15598 62242
rect 15650 62190 15652 62242
rect 15148 62188 15652 62190
rect 12572 62076 13188 62132
rect 11788 61682 12292 61684
rect 11788 61630 12238 61682
rect 12290 61630 12292 61682
rect 11788 61628 12292 61630
rect 11004 60900 11060 60910
rect 10780 60788 10836 60798
rect 10780 60694 10836 60732
rect 10556 60162 10612 60172
rect 11004 60004 11060 60844
rect 11564 60788 11620 60798
rect 11116 60786 11620 60788
rect 11116 60734 11566 60786
rect 11618 60734 11620 60786
rect 11116 60732 11620 60734
rect 11116 60674 11172 60732
rect 11564 60722 11620 60732
rect 11116 60622 11118 60674
rect 11170 60622 11172 60674
rect 11116 60610 11172 60622
rect 11788 60452 11844 61628
rect 12236 61618 12292 61628
rect 13020 60900 13076 60910
rect 12572 60898 13076 60900
rect 12572 60846 13022 60898
rect 13074 60846 13076 60898
rect 12572 60844 13076 60846
rect 11676 60396 11844 60452
rect 11900 60786 11956 60798
rect 11900 60734 11902 60786
rect 11954 60734 11956 60786
rect 11228 60114 11284 60126
rect 11228 60062 11230 60114
rect 11282 60062 11284 60114
rect 11228 60004 11284 60062
rect 10668 59948 11284 60004
rect 11340 60004 11396 60014
rect 10220 58546 10612 58548
rect 10220 58494 10222 58546
rect 10274 58494 10612 58546
rect 10220 58492 10612 58494
rect 10220 58482 10276 58492
rect 10556 58100 10612 58492
rect 10668 58322 10724 59948
rect 11340 59442 11396 59948
rect 11676 60002 11732 60396
rect 11788 60116 11844 60126
rect 11788 60022 11844 60060
rect 11676 59950 11678 60002
rect 11730 59950 11732 60002
rect 11676 59938 11732 59950
rect 11340 59390 11342 59442
rect 11394 59390 11396 59442
rect 11340 59332 11396 59390
rect 11340 59266 11396 59276
rect 11900 58884 11956 60734
rect 12572 60786 12628 60844
rect 13020 60834 13076 60844
rect 12572 60734 12574 60786
rect 12626 60734 12628 60786
rect 12572 60722 12628 60734
rect 12684 60676 12740 60686
rect 13132 60676 13188 62076
rect 13804 62076 14084 62132
rect 13244 60900 13300 60910
rect 13244 60806 13300 60844
rect 13356 60788 13412 60798
rect 13356 60694 13412 60732
rect 12684 60674 13188 60676
rect 12684 60622 12686 60674
rect 12738 60622 13188 60674
rect 12684 60620 13188 60622
rect 12684 60610 12740 60620
rect 12460 60002 12516 60014
rect 12460 59950 12462 60002
rect 12514 59950 12516 60002
rect 12012 59892 12068 59902
rect 12012 59890 12292 59892
rect 12012 59838 12014 59890
rect 12066 59838 12292 59890
rect 12012 59836 12292 59838
rect 12012 59826 12068 59836
rect 12236 59444 12292 59836
rect 12460 59780 12516 59950
rect 12908 60004 12964 60014
rect 12908 59910 12964 59948
rect 13804 59892 13860 62076
rect 14588 60788 14644 60798
rect 13916 60676 13972 60686
rect 14252 60676 14308 60686
rect 13916 60674 14308 60676
rect 13916 60622 13918 60674
rect 13970 60622 14254 60674
rect 14306 60622 14308 60674
rect 13916 60620 14308 60622
rect 13916 60610 13972 60620
rect 12460 59714 12516 59724
rect 13692 59890 13860 59892
rect 13692 59838 13806 59890
rect 13858 59838 13860 59890
rect 13692 59836 13860 59838
rect 12236 59388 12404 59444
rect 11788 58828 11956 58884
rect 12236 59218 12292 59230
rect 12236 59166 12238 59218
rect 12290 59166 12292 59218
rect 11788 58434 11844 58828
rect 12236 58772 12292 59166
rect 11788 58382 11790 58434
rect 11842 58382 11844 58434
rect 10668 58270 10670 58322
rect 10722 58270 10724 58322
rect 10668 58258 10724 58270
rect 11004 58324 11060 58334
rect 10556 58044 10836 58100
rect 9884 57876 9940 57886
rect 10556 57876 10612 57886
rect 9548 57874 10612 57876
rect 9548 57822 9886 57874
rect 9938 57822 10558 57874
rect 10610 57822 10612 57874
rect 9548 57820 10612 57822
rect 9436 57652 9492 57662
rect 9436 57558 9492 57596
rect 9548 56978 9604 57820
rect 9884 57810 9940 57820
rect 10108 57652 10164 57662
rect 10332 57652 10388 57662
rect 10108 57558 10164 57596
rect 10220 57650 10388 57652
rect 10220 57598 10334 57650
rect 10386 57598 10388 57650
rect 10220 57596 10388 57598
rect 9996 57538 10052 57550
rect 9996 57486 9998 57538
rect 10050 57486 10052 57538
rect 9996 57092 10052 57486
rect 9996 57026 10052 57036
rect 9548 56926 9550 56978
rect 9602 56926 9604 56978
rect 9548 56914 9604 56926
rect 8652 56802 8708 56812
rect 9772 56868 9828 56878
rect 8764 56756 8820 56766
rect 8652 56308 8708 56318
rect 8540 56306 8708 56308
rect 8540 56254 8654 56306
rect 8706 56254 8708 56306
rect 8540 56252 8708 56254
rect 8652 56242 8708 56252
rect 8764 56308 8820 56700
rect 8764 56214 8820 56252
rect 9772 56306 9828 56812
rect 9884 56756 9940 56766
rect 9884 56662 9940 56700
rect 9772 56254 9774 56306
rect 9826 56254 9828 56306
rect 9772 56242 9828 56254
rect 9212 56196 9268 56206
rect 8540 56084 8596 56094
rect 8428 56082 9044 56084
rect 8428 56030 8542 56082
rect 8594 56030 9044 56082
rect 8428 56028 9044 56030
rect 8540 56018 8596 56028
rect 6636 55412 7252 55468
rect 5068 54124 5348 54180
rect 5404 54628 5460 54638
rect 5068 53730 5124 54124
rect 5068 53678 5070 53730
rect 5122 53678 5124 53730
rect 5068 53666 5124 53678
rect 4956 52994 5012 53004
rect 5180 52946 5236 52958
rect 5180 52894 5182 52946
rect 5234 52894 5236 52946
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 3836 52164 3892 52174
rect 3388 51490 3444 51502
rect 3388 51438 3390 51490
rect 3442 51438 3444 51490
rect 3276 51378 3332 51390
rect 3276 51326 3278 51378
rect 3330 51326 3332 51378
rect 3276 51268 3332 51326
rect 3276 51202 3332 51212
rect 3388 51380 3444 51438
rect 2492 50482 2548 50494
rect 2492 50430 2494 50482
rect 2546 50430 2548 50482
rect 2492 50036 2548 50430
rect 2492 49970 2548 49980
rect 3388 49810 3444 51324
rect 3612 51378 3668 51390
rect 3612 51326 3614 51378
rect 3666 51326 3668 51378
rect 3612 50596 3668 51326
rect 3612 50530 3668 50540
rect 3836 51378 3892 52108
rect 4620 52164 4676 52174
rect 4620 52070 4676 52108
rect 4172 51380 4228 51390
rect 3836 51326 3838 51378
rect 3890 51326 3892 51378
rect 3388 49758 3390 49810
rect 3442 49758 3444 49810
rect 3388 49746 3444 49758
rect 2492 47348 2548 47358
rect 2492 47346 2660 47348
rect 2492 47294 2494 47346
rect 2546 47294 2660 47346
rect 2492 47292 2660 47294
rect 2492 47282 2548 47292
rect 2604 46898 2660 47292
rect 2604 46846 2606 46898
rect 2658 46846 2660 46898
rect 2604 46834 2660 46846
rect 2492 46786 2548 46798
rect 2492 46734 2494 46786
rect 2546 46734 2548 46786
rect 2492 46340 2548 46734
rect 2716 46564 2772 46574
rect 3164 46564 3220 46574
rect 2716 46470 2772 46508
rect 2828 46562 3220 46564
rect 2828 46510 3166 46562
rect 3218 46510 3220 46562
rect 2828 46508 3220 46510
rect 2828 46340 2884 46508
rect 2492 46284 2884 46340
rect 2492 44324 2548 46284
rect 3052 45330 3108 46508
rect 3164 46498 3220 46508
rect 3500 46564 3556 46574
rect 3500 46470 3556 46508
rect 3052 45278 3054 45330
rect 3106 45278 3108 45330
rect 3052 45266 3108 45278
rect 3500 44546 3556 44558
rect 3500 44494 3502 44546
rect 3554 44494 3556 44546
rect 2156 43652 2324 43708
rect 2380 44322 2548 44324
rect 2380 44270 2494 44322
rect 2546 44270 2548 44322
rect 2380 44268 2548 44270
rect 2380 43764 2436 44268
rect 2492 44258 2548 44268
rect 3388 44436 3444 44446
rect 3500 44436 3556 44494
rect 3836 44436 3892 51326
rect 4060 51378 4228 51380
rect 4060 51326 4174 51378
rect 4226 51326 4228 51378
rect 4060 51324 4228 51326
rect 3948 51268 4004 51278
rect 3948 49810 4004 51212
rect 4060 50484 4116 51324
rect 4172 51314 4228 51324
rect 4396 51378 4452 51390
rect 4396 51326 4398 51378
rect 4450 51326 4452 51378
rect 4284 51266 4340 51278
rect 4284 51214 4286 51266
rect 4338 51214 4340 51266
rect 4284 51156 4340 51214
rect 4172 51100 4340 51156
rect 4396 51156 4452 51326
rect 4172 50596 4228 51100
rect 4396 51090 4452 51100
rect 5068 51380 5124 51390
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 5068 50818 5124 51324
rect 5068 50766 5070 50818
rect 5122 50766 5124 50818
rect 5068 50754 5124 50766
rect 4620 50708 4676 50718
rect 4620 50706 5012 50708
rect 4620 50654 4622 50706
rect 4674 50654 5012 50706
rect 4620 50652 5012 50654
rect 4620 50642 4676 50652
rect 4172 50540 4564 50596
rect 4508 50484 4564 50540
rect 4956 50594 5012 50652
rect 4956 50542 4958 50594
rect 5010 50542 5012 50594
rect 4956 50530 5012 50542
rect 4508 50428 4900 50484
rect 4060 50418 4116 50428
rect 4284 50372 4340 50382
rect 4060 49924 4116 49934
rect 4284 49924 4340 50316
rect 4732 50260 4788 50270
rect 4508 50036 4564 50046
rect 4508 49942 4564 49980
rect 4060 49922 4340 49924
rect 4060 49870 4062 49922
rect 4114 49870 4340 49922
rect 4060 49868 4340 49870
rect 4060 49858 4116 49868
rect 3948 49758 3950 49810
rect 4002 49758 4004 49810
rect 3948 49746 4004 49758
rect 4284 49810 4340 49868
rect 4284 49758 4286 49810
rect 4338 49758 4340 49810
rect 4284 49746 4340 49758
rect 4732 49810 4788 50204
rect 4732 49758 4734 49810
rect 4786 49758 4788 49810
rect 4732 49588 4788 49758
rect 4844 49810 4900 50428
rect 5180 50428 5236 52894
rect 5404 51490 5460 54572
rect 5964 53508 6020 53518
rect 5964 53058 6020 53452
rect 5964 53006 5966 53058
rect 6018 53006 6020 53058
rect 5964 52994 6020 53006
rect 5404 51438 5406 51490
rect 5458 51438 5460 51490
rect 5404 51426 5460 51438
rect 5740 51378 5796 51390
rect 5740 51326 5742 51378
rect 5794 51326 5796 51378
rect 5516 51268 5572 51278
rect 5516 50708 5572 51212
rect 5740 50818 5796 51326
rect 5740 50766 5742 50818
rect 5794 50766 5796 50818
rect 5740 50754 5796 50766
rect 5516 50642 5572 50652
rect 5628 50596 5684 50606
rect 5628 50502 5684 50540
rect 5740 50484 5796 50494
rect 5180 50372 5460 50428
rect 5740 50390 5796 50428
rect 4844 49758 4846 49810
rect 4898 49758 4900 49810
rect 4844 49746 4900 49758
rect 5404 49698 5460 50372
rect 5404 49646 5406 49698
rect 5458 49646 5460 49698
rect 4732 49532 4900 49588
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4844 48354 4900 49532
rect 5404 49028 5460 49646
rect 4844 48302 4846 48354
rect 4898 48302 4900 48354
rect 4844 48290 4900 48302
rect 5068 48972 5404 49028
rect 4732 48242 4788 48254
rect 4732 48190 4734 48242
rect 4786 48190 4788 48242
rect 4732 48020 4788 48190
rect 4284 47964 4788 48020
rect 4172 46676 4228 46686
rect 4284 46676 4340 47964
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4620 47570 4676 47582
rect 4620 47518 4622 47570
rect 4674 47518 4676 47570
rect 4620 47348 4676 47518
rect 5068 47572 5124 48972
rect 5404 48962 5460 48972
rect 6076 49028 6132 49038
rect 6076 48934 6132 48972
rect 6188 48356 6244 48366
rect 6076 48354 6244 48356
rect 6076 48302 6190 48354
rect 6242 48302 6244 48354
rect 6076 48300 6244 48302
rect 5740 48244 5796 48254
rect 5964 48244 6020 48254
rect 5740 48242 6020 48244
rect 5740 48190 5742 48242
rect 5794 48190 5966 48242
rect 6018 48190 6020 48242
rect 5740 48188 6020 48190
rect 5740 48178 5796 48188
rect 5964 48178 6020 48188
rect 5180 48130 5236 48142
rect 5180 48078 5182 48130
rect 5234 48078 5236 48130
rect 5180 47684 5236 48078
rect 5628 47684 5684 47694
rect 5180 47682 5684 47684
rect 5180 47630 5630 47682
rect 5682 47630 5684 47682
rect 5180 47628 5684 47630
rect 5628 47618 5684 47628
rect 6076 47572 6132 48300
rect 6188 48290 6244 48300
rect 5124 47516 5460 47572
rect 5068 47478 5124 47516
rect 4620 47282 4676 47292
rect 5292 47348 5348 47358
rect 5292 46786 5348 47292
rect 5292 46734 5294 46786
rect 5346 46734 5348 46786
rect 5292 46722 5348 46734
rect 4172 46674 4340 46676
rect 4172 46622 4174 46674
rect 4226 46622 4340 46674
rect 4172 46620 4340 46622
rect 3500 44380 3780 44436
rect 3836 44380 4116 44436
rect 2828 44210 2884 44222
rect 2828 44158 2830 44210
rect 2882 44158 2884 44210
rect 2716 44100 2772 44110
rect 2380 43698 2436 43708
rect 2492 44098 2772 44100
rect 2492 44046 2718 44098
rect 2770 44046 2772 44098
rect 2492 44044 2772 44046
rect 1820 43538 1876 43550
rect 1820 43486 1822 43538
rect 1874 43486 1876 43538
rect 1820 42084 1876 43486
rect 1820 40402 1876 42028
rect 1820 40350 1822 40402
rect 1874 40350 1876 40402
rect 1820 40338 1876 40350
rect 1820 37492 1876 37502
rect 1820 36482 1876 37436
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1820 36418 1876 36430
rect 1820 35698 1876 35710
rect 1820 35646 1822 35698
rect 1874 35646 1876 35698
rect 1820 35028 1876 35646
rect 1820 34934 1876 34972
rect 2156 31948 2212 43652
rect 2492 43650 2548 44044
rect 2716 44034 2772 44044
rect 2492 43598 2494 43650
rect 2546 43598 2548 43650
rect 2492 43586 2548 43598
rect 2604 43764 2660 43774
rect 2604 41972 2660 43708
rect 2828 42868 2884 44158
rect 3388 44212 3444 44380
rect 3500 44212 3556 44222
rect 3388 44210 3556 44212
rect 3388 44158 3502 44210
rect 3554 44158 3556 44210
rect 3388 44156 3556 44158
rect 3500 44146 3556 44156
rect 3612 44210 3668 44222
rect 3612 44158 3614 44210
rect 3666 44158 3668 44210
rect 3612 43652 3668 44158
rect 3612 43586 3668 43596
rect 2940 42868 2996 42878
rect 2828 42866 2996 42868
rect 2828 42814 2942 42866
rect 2994 42814 2996 42866
rect 2828 42812 2996 42814
rect 2940 42802 2996 42812
rect 3724 42866 3780 44380
rect 3724 42814 3726 42866
rect 3778 42814 3780 42866
rect 3724 42802 3780 42814
rect 3948 44210 4004 44222
rect 3948 44158 3950 44210
rect 4002 44158 4004 44210
rect 3612 42754 3668 42766
rect 3612 42702 3614 42754
rect 3666 42702 3668 42754
rect 3612 42644 3668 42702
rect 3948 42644 4004 44158
rect 3612 42588 4004 42644
rect 2604 41916 2884 41972
rect 2828 41412 2884 41916
rect 2716 41300 2772 41310
rect 2492 41298 2772 41300
rect 2492 41246 2718 41298
rect 2770 41246 2772 41298
rect 2492 41244 2772 41246
rect 2492 40514 2548 41244
rect 2716 41234 2772 41244
rect 2828 41074 2884 41356
rect 3276 41858 3332 41870
rect 3276 41806 3278 41858
rect 3330 41806 3332 41858
rect 3276 41412 3332 41806
rect 3276 41346 3332 41356
rect 3052 41076 3108 41086
rect 2828 41022 2830 41074
rect 2882 41022 2884 41074
rect 2828 41010 2884 41022
rect 2940 41074 3108 41076
rect 2940 41022 3054 41074
rect 3106 41022 3108 41074
rect 2940 41020 3108 41022
rect 3612 41076 3668 42588
rect 4060 41412 4116 44380
rect 4172 44434 4228 46620
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4956 45220 5012 45230
rect 4844 45218 5012 45220
rect 4844 45166 4958 45218
rect 5010 45166 5012 45218
rect 4844 45164 5012 45166
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4172 44382 4174 44434
rect 4226 44382 4228 44434
rect 4172 44370 4228 44382
rect 4508 44436 4564 44446
rect 4508 44322 4564 44380
rect 4508 44270 4510 44322
rect 4562 44270 4564 44322
rect 4508 44258 4564 44270
rect 4844 44324 4900 45164
rect 4956 45154 5012 45164
rect 5068 45108 5124 45118
rect 5068 45106 5236 45108
rect 5068 45054 5070 45106
rect 5122 45054 5236 45106
rect 5068 45052 5236 45054
rect 5068 45042 5124 45052
rect 4956 44882 5012 44894
rect 4956 44830 4958 44882
rect 5010 44830 5012 44882
rect 4956 44548 5012 44830
rect 5180 44548 5236 45052
rect 5292 44548 5348 44558
rect 4956 44492 5124 44548
rect 5180 44492 5292 44548
rect 4620 43428 4676 43438
rect 4844 43428 4900 44268
rect 4956 44322 5012 44334
rect 4956 44270 4958 44322
rect 5010 44270 5012 44322
rect 4956 43762 5012 44270
rect 4956 43710 4958 43762
rect 5010 43710 5012 43762
rect 4956 43698 5012 43710
rect 5068 43652 5124 44492
rect 5292 44482 5348 44492
rect 5068 43558 5124 43596
rect 5404 43652 5460 47516
rect 5740 47516 6132 47572
rect 6300 48242 6356 48254
rect 6300 48190 6302 48242
rect 6354 48190 6356 48242
rect 5740 47348 5796 47516
rect 5740 47254 5796 47292
rect 5964 47348 6020 47358
rect 6300 47348 6356 48190
rect 5964 47346 6356 47348
rect 5964 47294 5966 47346
rect 6018 47294 6356 47346
rect 5964 47292 6356 47294
rect 5964 47282 6020 47292
rect 5516 47012 5572 47022
rect 5516 46562 5572 46956
rect 6300 47012 6356 47292
rect 6300 46946 6356 46956
rect 5516 46510 5518 46562
rect 5570 46510 5572 46562
rect 5516 46498 5572 46510
rect 6076 45108 6132 45118
rect 6076 45014 6132 45052
rect 5964 44548 6020 44558
rect 5964 44454 6020 44492
rect 5628 44436 5684 44446
rect 5628 44342 5684 44380
rect 6188 44324 6244 44334
rect 6188 44230 6244 44268
rect 5516 43652 5572 43662
rect 5404 43596 5516 43652
rect 4620 43426 4900 43428
rect 4620 43374 4622 43426
rect 4674 43374 4900 43426
rect 4620 43372 4900 43374
rect 4620 43362 4676 43372
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 5068 42084 5124 42094
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 3836 41356 4116 41412
rect 3724 41076 3780 41086
rect 3612 41074 3780 41076
rect 3612 41022 3726 41074
rect 3778 41022 3780 41074
rect 3612 41020 3780 41022
rect 2492 40462 2494 40514
rect 2546 40462 2548 40514
rect 2492 40450 2548 40462
rect 2828 39396 2884 39406
rect 2940 39396 2996 41020
rect 3052 41010 3108 41020
rect 3724 41010 3780 41020
rect 3836 39732 3892 41356
rect 4172 41298 4228 41310
rect 4172 41246 4174 41298
rect 4226 41246 4228 41298
rect 4060 41188 4116 41198
rect 3836 39666 3892 39676
rect 3948 41186 4116 41188
rect 3948 41134 4062 41186
rect 4114 41134 4116 41186
rect 3948 41132 4116 41134
rect 3164 39620 3220 39630
rect 3164 39526 3220 39564
rect 3948 39620 4004 41132
rect 4060 41122 4116 41132
rect 4172 39844 4228 41246
rect 5068 40626 5124 42028
rect 5404 42084 5460 43596
rect 5516 43558 5572 43596
rect 5404 41970 5460 42028
rect 5404 41918 5406 41970
rect 5458 41918 5460 41970
rect 5404 41906 5460 41918
rect 6076 41860 6132 41870
rect 6076 41766 6132 41804
rect 5180 41188 5236 41198
rect 5516 41188 5572 41198
rect 5180 41186 5572 41188
rect 5180 41134 5182 41186
rect 5234 41134 5518 41186
rect 5570 41134 5572 41186
rect 5180 41132 5572 41134
rect 5180 41122 5236 41132
rect 5516 41122 5572 41132
rect 5852 41074 5908 41086
rect 5852 41022 5854 41074
rect 5906 41022 5908 41074
rect 5068 40574 5070 40626
rect 5122 40574 5124 40626
rect 4620 40292 4676 40302
rect 4172 39778 4228 39788
rect 4284 40236 4620 40292
rect 2828 39394 2996 39396
rect 2828 39342 2830 39394
rect 2882 39342 2996 39394
rect 2828 39340 2996 39342
rect 2828 39330 2884 39340
rect 3948 38274 4004 39564
rect 4284 39506 4340 40236
rect 4620 40198 4676 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4284 39454 4286 39506
rect 4338 39454 4340 39506
rect 4284 39442 4340 39454
rect 4396 39732 4452 39742
rect 4396 38724 4452 39676
rect 4620 39732 4676 39742
rect 4620 39638 4676 39676
rect 4396 38612 4452 38668
rect 3948 38222 3950 38274
rect 4002 38222 4004 38274
rect 3948 38210 4004 38222
rect 4284 38556 4452 38612
rect 4284 38276 4340 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4284 38220 4564 38276
rect 4060 38052 4116 38062
rect 3612 37996 4060 38052
rect 2716 37604 2772 37614
rect 2716 37378 2772 37548
rect 3612 37604 3668 37996
rect 4060 37958 4116 37996
rect 3612 37490 3668 37548
rect 3612 37438 3614 37490
rect 3666 37438 3668 37490
rect 3612 37426 3668 37438
rect 3948 37826 4004 37838
rect 3948 37774 3950 37826
rect 4002 37774 4004 37826
rect 2716 37326 2718 37378
rect 2770 37326 2772 37378
rect 2716 37314 2772 37326
rect 3052 37380 3108 37390
rect 3052 37286 3108 37324
rect 3948 37380 4004 37774
rect 3164 37268 3220 37278
rect 3164 37174 3220 37212
rect 3724 37268 3780 37278
rect 3724 37174 3780 37212
rect 3836 37268 3892 37278
rect 3948 37268 4004 37324
rect 3836 37266 4004 37268
rect 3836 37214 3838 37266
rect 3890 37214 4004 37266
rect 3836 37212 4004 37214
rect 4284 37266 4340 38220
rect 4508 38162 4564 38220
rect 4508 38110 4510 38162
rect 4562 38110 4564 38162
rect 4508 38098 4564 38110
rect 4284 37214 4286 37266
rect 4338 37214 4340 37266
rect 2828 37154 2884 37166
rect 2828 37102 2830 37154
rect 2882 37102 2884 37154
rect 2828 36820 2884 37102
rect 2492 36764 2884 36820
rect 2492 36594 2548 36764
rect 2492 36542 2494 36594
rect 2546 36542 2548 36594
rect 2492 36530 2548 36542
rect 3836 36596 3892 37212
rect 4284 37202 4340 37214
rect 4620 37492 4676 37502
rect 4620 37266 4676 37436
rect 4620 37214 4622 37266
rect 4674 37214 4676 37266
rect 4620 37202 4676 37214
rect 5068 37492 5124 40574
rect 5740 40962 5796 40974
rect 5740 40910 5742 40962
rect 5794 40910 5796 40962
rect 5740 40292 5796 40910
rect 5852 40964 5908 41022
rect 6524 40964 6580 40974
rect 5908 40908 6020 40964
rect 5852 40898 5908 40908
rect 5628 39844 5684 39854
rect 5628 39750 5684 39788
rect 5740 39506 5796 40236
rect 5964 39842 6020 40908
rect 5964 39790 5966 39842
rect 6018 39790 6020 39842
rect 5964 39778 6020 39790
rect 6188 40514 6244 40526
rect 6188 40462 6190 40514
rect 6242 40462 6244 40514
rect 6188 39732 6244 40462
rect 6524 40514 6580 40908
rect 6524 40462 6526 40514
rect 6578 40462 6580 40514
rect 6524 40450 6580 40462
rect 6636 39732 6692 55412
rect 6748 54404 6804 54414
rect 6748 52164 6804 54348
rect 8988 53954 9044 56028
rect 8988 53902 8990 53954
rect 9042 53902 9044 53954
rect 8988 53890 9044 53902
rect 7868 53730 7924 53742
rect 7868 53678 7870 53730
rect 7922 53678 7924 53730
rect 7084 53618 7140 53630
rect 7084 53566 7086 53618
rect 7138 53566 7140 53618
rect 7084 52836 7140 53566
rect 7420 53620 7476 53630
rect 7420 53526 7476 53564
rect 7644 53618 7700 53630
rect 7644 53566 7646 53618
rect 7698 53566 7700 53618
rect 7196 53508 7252 53518
rect 7196 53414 7252 53452
rect 7644 53172 7700 53566
rect 7868 53620 7924 53678
rect 8428 53732 8484 53742
rect 8876 53732 8932 53742
rect 8428 53730 8932 53732
rect 8428 53678 8430 53730
rect 8482 53678 8878 53730
rect 8930 53678 8932 53730
rect 8428 53676 8932 53678
rect 8428 53666 8484 53676
rect 8876 53666 8932 53676
rect 7868 53554 7924 53564
rect 9100 53620 9156 53630
rect 8316 53508 8372 53518
rect 7644 53106 7700 53116
rect 8092 53506 8372 53508
rect 8092 53454 8318 53506
rect 8370 53454 8372 53506
rect 8092 53452 8372 53454
rect 7308 52836 7364 52846
rect 7084 52780 7308 52836
rect 7308 52274 7364 52780
rect 7308 52222 7310 52274
rect 7362 52222 7364 52274
rect 7308 52210 7364 52222
rect 8092 52834 8148 53452
rect 8316 53442 8372 53452
rect 8540 53506 8596 53518
rect 8540 53454 8542 53506
rect 8594 53454 8596 53506
rect 8540 53284 8596 53454
rect 8092 52782 8094 52834
rect 8146 52782 8148 52834
rect 6748 52098 6804 52108
rect 7980 52164 8036 52174
rect 8092 52164 8148 52782
rect 8204 53228 8596 53284
rect 8988 53506 9044 53518
rect 8988 53454 8990 53506
rect 9042 53454 9044 53506
rect 8204 52276 8260 53228
rect 8652 53172 8708 53182
rect 8988 53172 9044 53454
rect 8540 53116 8652 53172
rect 8540 53058 8596 53116
rect 8652 53106 8708 53116
rect 8764 53116 9044 53172
rect 8540 53006 8542 53058
rect 8594 53006 8596 53058
rect 8540 52994 8596 53006
rect 8428 52948 8484 52958
rect 8428 52854 8484 52892
rect 8652 52948 8708 52958
rect 8652 52500 8708 52892
rect 8204 52182 8260 52220
rect 8540 52444 8708 52500
rect 7980 52162 8148 52164
rect 7980 52110 7982 52162
rect 8034 52110 8148 52162
rect 7980 52108 8148 52110
rect 7980 52052 8036 52108
rect 7980 51986 8036 51996
rect 7644 51156 7700 51166
rect 6748 48916 6804 48926
rect 6748 48822 6804 48860
rect 7532 45220 7588 45230
rect 6748 44996 6804 45006
rect 6748 44994 7364 44996
rect 6748 44942 6750 44994
rect 6802 44942 7364 44994
rect 6748 44940 7364 44942
rect 6748 44930 6804 44940
rect 7196 44436 7252 44446
rect 7196 44322 7252 44380
rect 7308 44434 7364 44940
rect 7308 44382 7310 44434
rect 7362 44382 7364 44434
rect 7308 44370 7364 44382
rect 7196 44270 7198 44322
rect 7250 44270 7252 44322
rect 7196 44258 7252 44270
rect 7532 44322 7588 45164
rect 7532 44270 7534 44322
rect 7586 44270 7588 44322
rect 7532 44258 7588 44270
rect 7084 40404 7140 40414
rect 6860 39732 6916 39742
rect 6636 39730 6916 39732
rect 6636 39678 6862 39730
rect 6914 39678 6916 39730
rect 6636 39676 6916 39678
rect 6188 39666 6244 39676
rect 5740 39454 5742 39506
rect 5794 39454 5796 39506
rect 5740 39442 5796 39454
rect 6188 39060 6244 39070
rect 6188 38966 6244 39004
rect 6860 39060 6916 39676
rect 5852 38836 5908 38846
rect 5852 38050 5908 38780
rect 6412 38834 6468 38846
rect 6412 38782 6414 38834
rect 6466 38782 6468 38834
rect 6412 38612 6468 38782
rect 6636 38836 6692 38846
rect 6636 38742 6692 38780
rect 5852 37998 5854 38050
rect 5906 37998 5908 38050
rect 5852 37986 5908 37998
rect 6188 38556 6412 38612
rect 6188 38050 6244 38556
rect 6412 38546 6468 38556
rect 6524 38722 6580 38734
rect 6524 38670 6526 38722
rect 6578 38670 6580 38722
rect 6188 37998 6190 38050
rect 6242 37998 6244 38050
rect 6188 37986 6244 37998
rect 6412 38052 6468 38062
rect 6524 38052 6580 38670
rect 6860 38162 6916 39004
rect 7084 38836 7140 40348
rect 7084 38834 7252 38836
rect 7084 38782 7086 38834
rect 7138 38782 7252 38834
rect 7084 38780 7252 38782
rect 7084 38770 7140 38780
rect 6860 38110 6862 38162
rect 6914 38110 6916 38162
rect 6860 38098 6916 38110
rect 7084 38612 7140 38622
rect 6412 38050 6580 38052
rect 6412 37998 6414 38050
rect 6466 37998 6580 38050
rect 6412 37996 6580 37998
rect 6412 37986 6468 37996
rect 5964 37826 6020 37838
rect 5964 37774 5966 37826
rect 6018 37774 6020 37826
rect 5964 37604 6020 37774
rect 7084 37828 7140 38556
rect 7196 38164 7252 38780
rect 7420 38724 7476 38762
rect 7420 38658 7476 38668
rect 7644 38388 7700 51100
rect 8540 50484 8596 52444
rect 8764 52386 8820 53116
rect 8764 52334 8766 52386
rect 8818 52334 8820 52386
rect 8764 52322 8820 52334
rect 8988 52946 9044 52958
rect 8988 52894 8990 52946
rect 9042 52894 9044 52946
rect 8988 52724 9044 52894
rect 9100 52948 9156 53564
rect 9100 52882 9156 52892
rect 9212 52724 9268 56140
rect 10220 56082 10276 57596
rect 10332 57586 10388 57596
rect 10220 56030 10222 56082
rect 10274 56030 10276 56082
rect 10220 56018 10276 56030
rect 10444 57092 10500 57102
rect 10444 56082 10500 57036
rect 10556 56866 10612 57820
rect 10556 56814 10558 56866
rect 10610 56814 10612 56866
rect 10556 56802 10612 56814
rect 10668 57652 10724 57662
rect 10668 56978 10724 57596
rect 10780 57092 10836 58044
rect 10780 57026 10836 57036
rect 10668 56926 10670 56978
rect 10722 56926 10724 56978
rect 10444 56030 10446 56082
rect 10498 56030 10500 56082
rect 10444 56018 10500 56030
rect 10332 55524 10388 55534
rect 10332 53618 10388 55468
rect 10668 55468 10724 56926
rect 10780 56308 10836 56318
rect 11004 56308 11060 58268
rect 11788 58324 11844 58382
rect 11788 58258 11844 58268
rect 11900 58716 12236 58772
rect 10780 56306 11060 56308
rect 10780 56254 10782 56306
rect 10834 56254 11060 56306
rect 10780 56252 11060 56254
rect 11228 56644 11284 56654
rect 11228 56306 11284 56588
rect 11228 56254 11230 56306
rect 11282 56254 11284 56306
rect 10780 56242 10836 56252
rect 11228 56242 11284 56254
rect 11564 56084 11620 56094
rect 11788 56084 11844 56094
rect 11564 56082 11788 56084
rect 11564 56030 11566 56082
rect 11618 56030 11788 56082
rect 11564 56028 11788 56030
rect 11564 56018 11620 56028
rect 11004 55524 11060 55534
rect 10668 55412 10948 55468
rect 10892 55076 10948 55412
rect 11004 55298 11060 55468
rect 11788 55410 11844 56028
rect 11788 55358 11790 55410
rect 11842 55358 11844 55410
rect 11788 55346 11844 55358
rect 11004 55246 11006 55298
rect 11058 55246 11060 55298
rect 11004 55234 11060 55246
rect 11340 55300 11396 55310
rect 11340 55206 11396 55244
rect 11116 55076 11172 55086
rect 10892 55074 11172 55076
rect 10892 55022 11118 55074
rect 11170 55022 11172 55074
rect 10892 55020 11172 55022
rect 11004 54738 11060 55020
rect 11116 55010 11172 55020
rect 11004 54686 11006 54738
rect 11058 54686 11060 54738
rect 11004 54674 11060 54686
rect 10332 53566 10334 53618
rect 10386 53566 10388 53618
rect 10332 53554 10388 53566
rect 11340 54514 11396 54526
rect 11340 54462 11342 54514
rect 11394 54462 11396 54514
rect 10668 53508 10724 53518
rect 10668 53506 10836 53508
rect 10668 53454 10670 53506
rect 10722 53454 10836 53506
rect 10668 53452 10836 53454
rect 10668 53442 10724 53452
rect 9996 53060 10052 53070
rect 8988 52668 9268 52724
rect 9772 52834 9828 52846
rect 9772 52782 9774 52834
rect 9826 52782 9828 52834
rect 8652 52276 8708 52286
rect 8652 52162 8708 52220
rect 8652 52110 8654 52162
rect 8706 52110 8708 52162
rect 8652 52098 8708 52110
rect 8764 52052 8820 52062
rect 8764 51958 8820 51996
rect 8876 50484 8932 50494
rect 8540 50482 8932 50484
rect 8540 50430 8878 50482
rect 8930 50430 8932 50482
rect 8540 50428 8932 50430
rect 8876 50418 8932 50428
rect 8652 49924 8708 49934
rect 8652 49810 8708 49868
rect 8652 49758 8654 49810
rect 8706 49758 8708 49810
rect 7980 49700 8036 49710
rect 7980 49698 8372 49700
rect 7980 49646 7982 49698
rect 8034 49646 8372 49698
rect 7980 49644 8372 49646
rect 7980 49634 8036 49644
rect 8316 49028 8372 49644
rect 8540 49140 8596 49150
rect 8540 49028 8596 49084
rect 8316 48972 8596 49028
rect 8428 48804 8484 48814
rect 8316 48468 8372 48478
rect 8316 48374 8372 48412
rect 8428 48466 8484 48748
rect 8428 48414 8430 48466
rect 8482 48414 8484 48466
rect 8428 48402 8484 48414
rect 8540 48466 8596 48972
rect 8540 48414 8542 48466
rect 8594 48414 8596 48466
rect 8540 48402 8596 48414
rect 8092 48356 8148 48366
rect 8092 46228 8148 48300
rect 8652 48132 8708 49758
rect 8876 49812 8932 49822
rect 8876 49718 8932 49756
rect 8988 49588 9044 52668
rect 9660 52164 9716 52174
rect 9660 50932 9716 52108
rect 8764 49532 9044 49588
rect 9100 50876 9716 50932
rect 8764 48356 8820 49532
rect 9100 49364 9156 50876
rect 9772 50820 9828 52782
rect 9996 52050 10052 53004
rect 10332 53060 10388 53070
rect 10332 52946 10388 53004
rect 10332 52894 10334 52946
rect 10386 52894 10388 52946
rect 10332 52882 10388 52894
rect 10108 52834 10164 52846
rect 10108 52782 10110 52834
rect 10162 52782 10164 52834
rect 10108 52276 10164 52782
rect 10668 52836 10724 52846
rect 10780 52836 10836 53452
rect 11340 52948 11396 54462
rect 11564 52948 11620 52958
rect 11340 52946 11620 52948
rect 11340 52894 11566 52946
rect 11618 52894 11620 52946
rect 11340 52892 11620 52894
rect 11116 52836 11172 52846
rect 10780 52834 11172 52836
rect 10780 52782 11118 52834
rect 11170 52782 11172 52834
rect 10780 52780 11172 52782
rect 10668 52742 10724 52780
rect 10108 52210 10164 52220
rect 10220 52164 10276 52174
rect 10220 52070 10276 52108
rect 9996 51998 9998 52050
rect 10050 51998 10052 52050
rect 9996 51986 10052 51998
rect 11116 51156 11172 52780
rect 11452 52276 11508 52286
rect 11452 52050 11508 52220
rect 11452 51998 11454 52050
rect 11506 51998 11508 52050
rect 11452 51986 11508 51998
rect 11116 51090 11172 51100
rect 11564 50932 11620 52892
rect 11788 51938 11844 51950
rect 11788 51886 11790 51938
rect 11842 51886 11844 51938
rect 11788 51604 11844 51886
rect 11788 51538 11844 51548
rect 11564 50866 11620 50876
rect 9772 50764 10052 50820
rect 9324 50706 9380 50718
rect 9324 50654 9326 50706
rect 9378 50654 9380 50706
rect 9212 50594 9268 50606
rect 9212 50542 9214 50594
rect 9266 50542 9268 50594
rect 9212 49924 9268 50542
rect 9212 49858 9268 49868
rect 9324 49812 9380 50654
rect 9884 50594 9940 50606
rect 9884 50542 9886 50594
rect 9938 50542 9940 50594
rect 9884 50428 9940 50542
rect 9436 50372 9940 50428
rect 9996 50428 10052 50764
rect 11564 50708 11620 50718
rect 11564 50614 11620 50652
rect 10780 50484 10836 50494
rect 11116 50484 11172 50494
rect 10668 50482 11172 50484
rect 10668 50430 10782 50482
rect 10834 50430 11118 50482
rect 11170 50430 11172 50482
rect 10668 50428 11172 50430
rect 9996 50372 10164 50428
rect 10668 50372 10836 50428
rect 11116 50418 11172 50428
rect 9436 50034 9492 50372
rect 9436 49982 9438 50034
rect 9490 49982 9492 50034
rect 9436 49970 9492 49982
rect 9660 49924 9716 49934
rect 9324 49746 9380 49756
rect 9548 49922 9716 49924
rect 9548 49870 9662 49922
rect 9714 49870 9716 49922
rect 9548 49868 9716 49870
rect 9100 49308 9268 49364
rect 8764 48290 8820 48300
rect 8876 49138 8932 49150
rect 8876 49086 8878 49138
rect 8930 49086 8932 49138
rect 8876 48354 8932 49086
rect 9100 49140 9156 49150
rect 9100 49026 9156 49084
rect 9100 48974 9102 49026
rect 9154 48974 9156 49026
rect 9100 48962 9156 48974
rect 8876 48302 8878 48354
rect 8930 48302 8932 48354
rect 8876 48290 8932 48302
rect 8988 48132 9044 48142
rect 8652 48130 9044 48132
rect 8652 48078 8990 48130
rect 9042 48078 9044 48130
rect 8652 48076 9044 48078
rect 8988 48066 9044 48076
rect 8876 46786 8932 46798
rect 8876 46734 8878 46786
rect 8930 46734 8932 46786
rect 8764 46674 8820 46686
rect 8764 46622 8766 46674
rect 8818 46622 8820 46674
rect 8092 46172 8484 46228
rect 8092 45666 8148 45678
rect 8092 45614 8094 45666
rect 8146 45614 8148 45666
rect 8092 44436 8148 45614
rect 8092 44342 8148 44380
rect 8204 45666 8260 45678
rect 8204 45614 8206 45666
rect 8258 45614 8260 45666
rect 7756 44212 7812 44222
rect 8204 44212 8260 45614
rect 8316 45666 8372 45678
rect 8316 45614 8318 45666
rect 8370 45614 8372 45666
rect 8316 45332 8372 45614
rect 8316 45266 8372 45276
rect 8428 45668 8484 46172
rect 8540 45668 8596 45678
rect 8428 45666 8596 45668
rect 8428 45614 8542 45666
rect 8594 45614 8596 45666
rect 8428 45612 8596 45614
rect 8428 45108 8484 45612
rect 8540 45602 8596 45612
rect 8764 45668 8820 46622
rect 8764 45602 8820 45612
rect 7756 44210 8260 44212
rect 7756 44158 7758 44210
rect 7810 44158 8260 44210
rect 7756 44156 8260 44158
rect 8316 45052 8484 45108
rect 8876 45332 8932 46734
rect 9100 46674 9156 46686
rect 9100 46622 9102 46674
rect 9154 46622 9156 46674
rect 9100 46002 9156 46622
rect 9100 45950 9102 46002
rect 9154 45950 9156 46002
rect 9100 45938 9156 45950
rect 7756 44146 7812 44156
rect 8316 44100 8372 45052
rect 8876 44996 8932 45276
rect 8764 44994 8932 44996
rect 8764 44942 8878 44994
rect 8930 44942 8932 44994
rect 8764 44940 8932 44942
rect 8764 44322 8820 44940
rect 8876 44930 8932 44940
rect 8988 45668 9044 45678
rect 8988 44434 9044 45612
rect 8988 44382 8990 44434
rect 9042 44382 9044 44434
rect 8988 44370 9044 44382
rect 8764 44270 8766 44322
rect 8818 44270 8820 44322
rect 8764 44258 8820 44270
rect 8092 44044 8372 44100
rect 8092 40626 8148 44044
rect 8428 43652 8484 43662
rect 8428 42866 8484 43596
rect 8428 42814 8430 42866
rect 8482 42814 8484 42866
rect 8428 42802 8484 42814
rect 8876 42756 8932 42766
rect 8876 42662 8932 42700
rect 8764 42642 8820 42654
rect 8764 42590 8766 42642
rect 8818 42590 8820 42642
rect 8764 42532 8820 42590
rect 8988 42532 9044 42542
rect 8764 42466 8820 42476
rect 8876 42530 9044 42532
rect 8876 42478 8990 42530
rect 9042 42478 9044 42530
rect 8876 42476 9044 42478
rect 8204 41972 8260 41982
rect 8204 41858 8260 41916
rect 8876 41972 8932 42476
rect 8988 42466 9044 42476
rect 8876 41906 8932 41916
rect 8988 41970 9044 41982
rect 8988 41918 8990 41970
rect 9042 41918 9044 41970
rect 8204 41806 8206 41858
rect 8258 41806 8260 41858
rect 8204 41794 8260 41806
rect 8764 41860 8820 41870
rect 8764 41766 8820 41804
rect 8988 41860 9044 41918
rect 8988 41794 9044 41804
rect 8652 41746 8708 41758
rect 8652 41694 8654 41746
rect 8706 41694 8708 41746
rect 8540 41188 8596 41198
rect 8092 40574 8094 40626
rect 8146 40574 8148 40626
rect 8092 40562 8148 40574
rect 8204 41132 8540 41188
rect 7868 40404 7924 40414
rect 7868 40310 7924 40348
rect 8204 39058 8260 41132
rect 8540 41094 8596 41132
rect 8316 40964 8372 40974
rect 8652 40964 8708 41694
rect 8316 40962 8708 40964
rect 8316 40910 8318 40962
rect 8370 40910 8708 40962
rect 8316 40908 8708 40910
rect 8316 40898 8372 40908
rect 8204 39006 8206 39058
rect 8258 39006 8260 39058
rect 8204 38994 8260 39006
rect 8540 40404 8596 40414
rect 8540 40290 8596 40348
rect 8540 40238 8542 40290
rect 8594 40238 8596 40290
rect 8540 39172 8596 40238
rect 8540 39058 8596 39116
rect 8540 39006 8542 39058
rect 8594 39006 8596 39058
rect 8540 38994 8596 39006
rect 7980 38946 8036 38958
rect 7980 38894 7982 38946
rect 8034 38894 8036 38946
rect 7868 38836 7924 38846
rect 7868 38742 7924 38780
rect 7980 38612 8036 38894
rect 9212 38668 9268 49308
rect 9324 48916 9380 48926
rect 9324 48822 9380 48860
rect 9548 48914 9604 49868
rect 9660 49858 9716 49868
rect 9772 49812 9828 49822
rect 9996 49812 10052 49822
rect 9772 49810 10052 49812
rect 9772 49758 9774 49810
rect 9826 49758 9998 49810
rect 10050 49758 10052 49810
rect 9772 49756 10052 49758
rect 9772 49746 9828 49756
rect 9996 49746 10052 49756
rect 10108 49140 10164 50372
rect 10220 49924 10276 49934
rect 10220 49830 10276 49868
rect 10332 49812 10388 49822
rect 10332 49718 10388 49756
rect 10780 49700 10836 50372
rect 10220 49140 10276 49150
rect 10108 49138 10276 49140
rect 10108 49086 10222 49138
rect 10274 49086 10276 49138
rect 10108 49084 10276 49086
rect 9548 48862 9550 48914
rect 9602 48862 9604 48914
rect 9548 48468 9604 48862
rect 9660 49026 9716 49038
rect 9660 48974 9662 49026
rect 9714 48974 9716 49026
rect 9660 48804 9716 48974
rect 9660 48738 9716 48748
rect 10108 49028 10164 49084
rect 10220 49074 10276 49084
rect 9548 47684 9604 48412
rect 9548 47618 9604 47628
rect 9996 48356 10052 48366
rect 9660 47460 9716 47470
rect 9660 46114 9716 47404
rect 9660 46062 9662 46114
rect 9714 46062 9716 46114
rect 9660 46050 9716 46062
rect 9996 46002 10052 48300
rect 10108 46562 10164 48972
rect 10556 48356 10612 48366
rect 10556 48262 10612 48300
rect 10108 46510 10110 46562
rect 10162 46510 10164 46562
rect 10108 46498 10164 46510
rect 9996 45950 9998 46002
rect 10050 45950 10052 46002
rect 9996 45938 10052 45950
rect 9324 45892 9380 45902
rect 9324 45890 9604 45892
rect 9324 45838 9326 45890
rect 9378 45838 9604 45890
rect 9324 45836 9604 45838
rect 9324 45826 9380 45836
rect 9436 45444 9492 45454
rect 9436 45108 9492 45388
rect 9548 45332 9604 45836
rect 9996 45668 10052 45678
rect 9884 45612 9996 45668
rect 9660 45332 9716 45342
rect 9548 45330 9716 45332
rect 9548 45278 9662 45330
rect 9714 45278 9716 45330
rect 9548 45276 9716 45278
rect 9660 45266 9716 45276
rect 9772 45332 9828 45342
rect 9772 45238 9828 45276
rect 9436 44436 9492 45052
rect 9548 45108 9604 45118
rect 9884 45108 9940 45612
rect 9996 45602 10052 45612
rect 9548 45106 9940 45108
rect 9548 45054 9550 45106
rect 9602 45054 9940 45106
rect 9548 45052 9940 45054
rect 10108 45220 10164 45230
rect 10108 45106 10164 45164
rect 10108 45054 10110 45106
rect 10162 45054 10164 45106
rect 9548 45042 9604 45052
rect 9548 44436 9604 44446
rect 9436 44434 9604 44436
rect 9436 44382 9550 44434
rect 9602 44382 9604 44434
rect 9436 44380 9604 44382
rect 9548 44370 9604 44380
rect 10108 42978 10164 45054
rect 10108 42926 10110 42978
rect 10162 42926 10164 42978
rect 10108 42914 10164 42926
rect 9660 42756 9716 42766
rect 9660 42662 9716 42700
rect 10108 42754 10164 42766
rect 10108 42702 10110 42754
rect 10162 42702 10164 42754
rect 9772 42532 9828 42542
rect 9660 42196 9716 42206
rect 9436 42194 9716 42196
rect 9436 42142 9662 42194
rect 9714 42142 9716 42194
rect 9436 42140 9716 42142
rect 9436 41972 9492 42140
rect 9660 42130 9716 42140
rect 9436 40964 9492 41916
rect 9548 41972 9604 41982
rect 9772 41972 9828 42476
rect 9548 41970 9828 41972
rect 9548 41918 9550 41970
rect 9602 41918 9828 41970
rect 9548 41916 9828 41918
rect 9884 42196 9940 42206
rect 9884 41970 9940 42140
rect 9884 41918 9886 41970
rect 9938 41918 9940 41970
rect 9548 41186 9604 41916
rect 9884 41906 9940 41918
rect 9548 41134 9550 41186
rect 9602 41134 9604 41186
rect 9548 41122 9604 41134
rect 10108 41188 10164 42702
rect 10556 42754 10612 42766
rect 10556 42702 10558 42754
rect 10610 42702 10612 42754
rect 10556 42196 10612 42702
rect 10556 42130 10612 42140
rect 10332 41860 10388 41870
rect 10332 41766 10388 41804
rect 10108 41122 10164 41132
rect 9660 41074 9716 41086
rect 9660 41022 9662 41074
rect 9714 41022 9716 41074
rect 9660 40964 9716 41022
rect 9436 40908 9716 40964
rect 9884 38724 9940 38734
rect 9212 38612 9828 38668
rect 7980 38546 8036 38556
rect 7644 38332 8036 38388
rect 7756 38164 7812 38174
rect 7196 38162 7812 38164
rect 7196 38110 7758 38162
rect 7810 38110 7812 38162
rect 7196 38108 7812 38110
rect 7196 38050 7252 38108
rect 7756 38098 7812 38108
rect 7196 37998 7198 38050
rect 7250 37998 7252 38050
rect 7196 37986 7252 37998
rect 7084 37772 7476 37828
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36596 4676 36606
rect 3836 36594 4676 36596
rect 3836 36542 4622 36594
rect 4674 36542 4676 36594
rect 3836 36540 4676 36542
rect 5068 36596 5124 37436
rect 5292 37548 6020 37604
rect 5292 37378 5348 37548
rect 5292 37326 5294 37378
rect 5346 37326 5348 37378
rect 5292 37314 5348 37326
rect 7420 37154 7476 37772
rect 7868 37492 7924 37502
rect 7868 37398 7924 37436
rect 7420 37102 7422 37154
rect 7474 37102 7476 37154
rect 7420 37090 7476 37102
rect 7980 37044 8036 38332
rect 9772 38274 9828 38612
rect 9772 38222 9774 38274
rect 9826 38222 9828 38274
rect 9772 38210 9828 38222
rect 8540 38108 8820 38164
rect 8428 37380 8484 37390
rect 8428 37286 8484 37324
rect 7980 36978 8036 36988
rect 5180 36596 5236 36606
rect 5068 36594 5236 36596
rect 5068 36542 5182 36594
rect 5234 36542 5236 36594
rect 5068 36540 5236 36542
rect 4620 36530 4676 36540
rect 5180 36530 5236 36540
rect 8204 36484 8260 36494
rect 2268 35812 2324 35822
rect 2268 35718 2324 35756
rect 7868 35700 7924 35710
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 5852 34916 5908 34926
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 2156 31892 2324 31948
rect 2268 26292 2324 31892
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 29426 4340 29438
rect 4284 29374 4286 29426
rect 4338 29374 4340 29426
rect 4284 28644 4340 29374
rect 5068 29314 5124 29326
rect 5068 29262 5070 29314
rect 5122 29262 5124 29314
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 5068 28980 5124 29262
rect 5068 28914 5124 28924
rect 4284 28578 4340 28588
rect 4732 28644 4788 28654
rect 4732 27858 4788 28588
rect 4732 27806 4734 27858
rect 4786 27806 4788 27858
rect 4732 27794 4788 27806
rect 5404 27748 5460 27758
rect 5404 27654 5460 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 2268 26226 2324 26236
rect 5628 27076 5684 27086
rect 5628 26178 5684 27020
rect 5628 26126 5630 26178
rect 5682 26126 5684 26178
rect 5628 26114 5684 26126
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 5852 11732 5908 34860
rect 7308 34914 7364 34926
rect 7308 34862 7310 34914
rect 7362 34862 7364 34914
rect 7308 34132 7364 34862
rect 7532 34804 7588 34814
rect 7532 34710 7588 34748
rect 7868 34354 7924 35644
rect 8092 35476 8148 35486
rect 7868 34302 7870 34354
rect 7922 34302 7924 34354
rect 7756 34132 7812 34142
rect 7196 34130 7812 34132
rect 7196 34078 7758 34130
rect 7810 34078 7812 34130
rect 7196 34076 7812 34078
rect 7196 31948 7252 34076
rect 7756 34066 7812 34076
rect 7084 31892 7252 31948
rect 7420 33908 7476 33918
rect 7308 31892 7364 31902
rect 6972 28644 7028 28654
rect 6972 28550 7028 28588
rect 6748 27076 6804 27086
rect 6748 26982 6804 27020
rect 6972 26964 7028 26974
rect 7084 26964 7140 31892
rect 7308 31798 7364 31836
rect 7196 31778 7252 31790
rect 7196 31726 7198 31778
rect 7250 31726 7252 31778
rect 7196 30994 7252 31726
rect 7196 30942 7198 30994
rect 7250 30942 7252 30994
rect 7196 29428 7252 30942
rect 7196 29314 7252 29372
rect 7196 29262 7198 29314
rect 7250 29262 7252 29314
rect 7196 29250 7252 29262
rect 7308 28642 7364 28654
rect 7308 28590 7310 28642
rect 7362 28590 7364 28642
rect 7308 28196 7364 28590
rect 7420 28418 7476 33852
rect 7868 31892 7924 34302
rect 7980 34914 8036 34926
rect 7980 34862 7982 34914
rect 8034 34862 8036 34914
rect 7980 33908 8036 34862
rect 8092 34690 8148 35420
rect 8092 34638 8094 34690
rect 8146 34638 8148 34690
rect 8092 34626 8148 34638
rect 8092 34356 8148 34366
rect 8204 34356 8260 36428
rect 8540 36482 8596 38108
rect 8764 38050 8820 38108
rect 8764 37998 8766 38050
rect 8818 37998 8820 38050
rect 8764 37986 8820 37998
rect 9436 38050 9492 38062
rect 9436 37998 9438 38050
rect 9490 37998 9492 38050
rect 8540 36430 8542 36482
rect 8594 36430 8596 36482
rect 8540 36418 8596 36430
rect 8652 37938 8708 37950
rect 8652 37886 8654 37938
rect 8706 37886 8708 37938
rect 8652 37378 8708 37886
rect 8988 37492 9044 37502
rect 8988 37398 9044 37436
rect 9436 37492 9492 37998
rect 9436 37426 9492 37436
rect 8652 37326 8654 37378
rect 8706 37326 8708 37378
rect 8092 34354 8260 34356
rect 8092 34302 8094 34354
rect 8146 34302 8260 34354
rect 8092 34300 8260 34302
rect 8428 36260 8484 36270
rect 8092 34290 8148 34300
rect 8428 34242 8484 36204
rect 8652 35812 8708 37326
rect 8764 37378 8820 37390
rect 8764 37326 8766 37378
rect 8818 37326 8820 37378
rect 8764 36484 8820 37326
rect 9548 37380 9604 37390
rect 9436 37266 9492 37278
rect 9436 37214 9438 37266
rect 9490 37214 9492 37266
rect 8876 37156 8932 37166
rect 9436 37156 9492 37214
rect 8876 37154 9492 37156
rect 8876 37102 8878 37154
rect 8930 37102 9492 37154
rect 8876 37100 9492 37102
rect 8876 37090 8932 37100
rect 9324 36596 9380 36606
rect 9548 36596 9604 37324
rect 9660 37044 9716 37054
rect 9660 36950 9716 36988
rect 9324 36594 9604 36596
rect 9324 36542 9326 36594
rect 9378 36542 9604 36594
rect 9324 36540 9604 36542
rect 9324 36530 9380 36540
rect 8764 36418 8820 36428
rect 8876 36370 8932 36382
rect 8876 36318 8878 36370
rect 8930 36318 8932 36370
rect 8764 36260 8820 36270
rect 8876 36260 8932 36318
rect 8876 36204 9604 36260
rect 8764 36166 8820 36204
rect 8428 34190 8430 34242
rect 8482 34190 8484 34242
rect 8428 34178 8484 34190
rect 8540 35756 8708 35812
rect 8876 36036 8932 36046
rect 7980 33842 8036 33852
rect 7868 31332 7924 31836
rect 7868 31266 7924 31276
rect 7980 32564 8036 32574
rect 7756 30772 7812 30782
rect 7980 30772 8036 32508
rect 8540 31948 8596 35756
rect 8876 32788 8932 35980
rect 8988 34132 9044 34142
rect 8988 34130 9156 34132
rect 8988 34078 8990 34130
rect 9042 34078 9156 34130
rect 8988 34076 9156 34078
rect 8988 34066 9044 34076
rect 8988 32788 9044 32798
rect 8876 32786 9044 32788
rect 8876 32734 8990 32786
rect 9042 32734 9044 32786
rect 8876 32732 9044 32734
rect 8988 32722 9044 32732
rect 8428 31892 8596 31948
rect 8764 32562 8820 32574
rect 8764 32510 8766 32562
rect 8818 32510 8820 32562
rect 8764 31948 8820 32510
rect 9100 32116 9156 34076
rect 9548 34018 9604 36204
rect 9772 36258 9828 36270
rect 9772 36206 9774 36258
rect 9826 36206 9828 36258
rect 9772 36148 9828 36206
rect 9660 34356 9716 34366
rect 9772 34356 9828 36092
rect 9660 34354 9828 34356
rect 9660 34302 9662 34354
rect 9714 34302 9828 34354
rect 9660 34300 9828 34302
rect 9884 34914 9940 38668
rect 10668 37940 10724 37950
rect 10556 37938 10724 37940
rect 10556 37886 10670 37938
rect 10722 37886 10724 37938
rect 10556 37884 10724 37886
rect 9996 37492 10052 37502
rect 9996 37156 10052 37436
rect 10220 37268 10276 37278
rect 10556 37268 10612 37884
rect 10668 37874 10724 37884
rect 10780 37716 10836 49644
rect 11116 48914 11172 48926
rect 11116 48862 11118 48914
rect 11170 48862 11172 48914
rect 11116 48244 11172 48862
rect 11116 48150 11172 48188
rect 11228 48802 11284 48814
rect 11228 48750 11230 48802
rect 11282 48750 11284 48802
rect 11116 47684 11172 47694
rect 11116 47590 11172 47628
rect 11228 47570 11284 48750
rect 11228 47518 11230 47570
rect 11282 47518 11284 47570
rect 11228 47506 11284 47518
rect 11340 48802 11396 48814
rect 11340 48750 11342 48802
rect 11394 48750 11396 48802
rect 11340 48356 11396 48750
rect 11116 47460 11172 47470
rect 11116 47366 11172 47404
rect 11340 47348 11396 48300
rect 11788 48242 11844 48254
rect 11788 48190 11790 48242
rect 11842 48190 11844 48242
rect 11788 47460 11844 48190
rect 11788 47394 11844 47404
rect 11340 47282 11396 47292
rect 11788 46900 11844 46910
rect 11564 42084 11620 42094
rect 11564 41990 11620 42028
rect 11676 41970 11732 41982
rect 11676 41918 11678 41970
rect 11730 41918 11732 41970
rect 11676 41076 11732 41918
rect 11676 41010 11732 41020
rect 11452 39618 11508 39630
rect 11452 39566 11454 39618
rect 11506 39566 11508 39618
rect 11452 38948 11508 39566
rect 11340 38836 11396 38846
rect 11452 38836 11508 38892
rect 11340 38834 11508 38836
rect 11340 38782 11342 38834
rect 11394 38782 11508 38834
rect 11340 38780 11508 38782
rect 11564 39394 11620 39406
rect 11564 39342 11566 39394
rect 11618 39342 11620 39394
rect 11340 38770 11396 38780
rect 11564 38724 11620 39342
rect 11564 38658 11620 38668
rect 11004 38610 11060 38622
rect 11004 38558 11006 38610
rect 11058 38558 11060 38610
rect 11004 38052 11060 38558
rect 11788 38274 11844 46844
rect 11900 46676 11956 58716
rect 12236 58706 12292 58716
rect 12348 58546 12404 59388
rect 12796 59332 12852 59342
rect 12796 59106 12852 59276
rect 12796 59054 12798 59106
rect 12850 59054 12852 59106
rect 12796 58884 12852 59054
rect 12796 58818 12852 58828
rect 12348 58494 12350 58546
rect 12402 58494 12404 58546
rect 12348 58482 12404 58494
rect 13468 58324 13524 58334
rect 13692 58324 13748 59836
rect 13804 59826 13860 59836
rect 14028 60004 14084 60620
rect 14252 60610 14308 60620
rect 14140 60004 14196 60014
rect 14028 60002 14196 60004
rect 14028 59950 14142 60002
rect 14194 59950 14196 60002
rect 14028 59948 14196 59950
rect 13468 58322 13748 58324
rect 13468 58270 13470 58322
rect 13522 58270 13748 58322
rect 13468 58268 13748 58270
rect 14028 59780 14084 59948
rect 14140 59938 14196 59948
rect 13468 58258 13524 58268
rect 13804 58210 13860 58222
rect 13804 58158 13806 58210
rect 13858 58158 13860 58210
rect 13804 57764 13860 58158
rect 13804 57670 13860 57708
rect 13356 57652 13412 57662
rect 13356 57538 13412 57596
rect 13916 57652 13972 57662
rect 14028 57652 14084 59724
rect 14476 59220 14532 59230
rect 13972 57596 14084 57652
rect 14140 59218 14532 59220
rect 14140 59166 14478 59218
rect 14530 59166 14532 59218
rect 14140 59164 14532 59166
rect 13916 57558 13972 57596
rect 13356 57486 13358 57538
rect 13410 57486 13412 57538
rect 13356 57428 13412 57486
rect 13020 57372 13412 57428
rect 13804 57426 13860 57438
rect 13804 57374 13806 57426
rect 13858 57374 13860 57426
rect 12236 57092 12292 57102
rect 12124 57036 12236 57092
rect 12012 56754 12068 56766
rect 12012 56702 12014 56754
rect 12066 56702 12068 56754
rect 12012 56644 12068 56702
rect 12012 56578 12068 56588
rect 12124 56306 12180 57036
rect 12236 56998 12292 57036
rect 12572 56644 12628 56654
rect 12572 56550 12628 56588
rect 12124 56254 12126 56306
rect 12178 56254 12180 56306
rect 12124 56242 12180 56254
rect 12908 56194 12964 56206
rect 12908 56142 12910 56194
rect 12962 56142 12964 56194
rect 12460 56084 12516 56094
rect 12796 56084 12852 56094
rect 12460 56082 12852 56084
rect 12460 56030 12462 56082
rect 12514 56030 12798 56082
rect 12850 56030 12852 56082
rect 12460 56028 12852 56030
rect 12460 56018 12516 56028
rect 12684 55076 12740 56028
rect 12796 56018 12852 56028
rect 12908 56084 12964 56142
rect 12908 56018 12964 56028
rect 12684 54982 12740 55020
rect 12572 54516 12628 54526
rect 12572 53172 12628 54460
rect 13020 53284 13076 57372
rect 13692 56756 13748 56766
rect 13692 56306 13748 56700
rect 13804 56754 13860 57374
rect 14140 56978 14196 59164
rect 14476 59154 14532 59164
rect 14588 58772 14644 60732
rect 15596 60116 15652 62188
rect 16380 61684 16436 62300
rect 16044 61628 16436 61684
rect 15596 60050 15652 60060
rect 15708 60564 15764 60574
rect 15708 60114 15764 60508
rect 15708 60062 15710 60114
rect 15762 60062 15764 60114
rect 15708 60050 15764 60062
rect 15148 60004 15204 60014
rect 15036 59444 15092 59454
rect 15036 59350 15092 59388
rect 15148 59442 15204 59948
rect 15148 59390 15150 59442
rect 15202 59390 15204 59442
rect 15148 59378 15204 59390
rect 15260 60002 15316 60014
rect 15260 59950 15262 60002
rect 15314 59950 15316 60002
rect 14476 58548 14532 58558
rect 14588 58548 14644 58716
rect 14476 58546 14644 58548
rect 14476 58494 14478 58546
rect 14530 58494 14644 58546
rect 14476 58492 14644 58494
rect 14924 59218 14980 59230
rect 14924 59166 14926 59218
rect 14978 59166 14980 59218
rect 14476 58482 14532 58492
rect 14924 57764 14980 59166
rect 15260 58212 15316 59950
rect 15708 59444 15764 59454
rect 16044 59444 16100 61628
rect 17388 61124 17444 62860
rect 17836 62916 17892 62926
rect 17836 62822 17892 62860
rect 18508 62916 18564 62926
rect 18508 62822 18564 62860
rect 19404 62578 19460 63084
rect 19628 63074 19684 63084
rect 19964 63026 20020 63038
rect 19964 62974 19966 63026
rect 20018 62974 20020 63026
rect 19964 62916 20020 62974
rect 19404 62526 19406 62578
rect 19458 62526 19460 62578
rect 19404 62514 19460 62526
rect 19628 62860 20020 62916
rect 19628 62580 19684 62860
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19964 62580 20020 62590
rect 19628 62578 20020 62580
rect 19628 62526 19966 62578
rect 20018 62526 20020 62578
rect 19628 62524 20020 62526
rect 19964 62514 20020 62524
rect 18956 62468 19012 62478
rect 18732 62412 18956 62468
rect 20860 62468 20916 63758
rect 20972 63140 21028 63980
rect 21084 63364 21140 67172
rect 22876 66386 22932 69200
rect 24892 66500 24948 69200
rect 26908 67228 26964 69200
rect 28924 67228 28980 69200
rect 30940 67228 30996 69200
rect 32956 67228 33012 69200
rect 34972 67228 35028 69200
rect 26908 67172 27412 67228
rect 28924 67172 29204 67228
rect 30940 67172 31220 67228
rect 32956 67172 33236 67228
rect 34972 67172 35140 67228
rect 24892 66434 24948 66444
rect 26124 66500 26180 66510
rect 26124 66406 26180 66444
rect 22876 66334 22878 66386
rect 22930 66334 22932 66386
rect 22876 66322 22932 66334
rect 23548 66274 23604 66286
rect 25116 66276 25172 66286
rect 23548 66222 23550 66274
rect 23602 66222 23604 66274
rect 21868 65490 21924 65502
rect 23548 65492 23604 66222
rect 21868 65438 21870 65490
rect 21922 65438 21924 65490
rect 21420 64484 21476 64494
rect 21420 64390 21476 64428
rect 21868 64484 21924 65438
rect 22988 65436 23604 65492
rect 24668 66274 25172 66276
rect 24668 66222 25118 66274
rect 25170 66222 25172 66274
rect 24668 66220 25172 66222
rect 22540 65378 22596 65390
rect 22540 65326 22542 65378
rect 22594 65326 22596 65378
rect 22540 64932 22596 65326
rect 22540 64866 22596 64876
rect 21868 64418 21924 64428
rect 22988 63810 23044 65436
rect 24668 65378 24724 66220
rect 25116 66210 25172 66220
rect 24668 65326 24670 65378
rect 24722 65326 24724 65378
rect 24668 65314 24724 65326
rect 25452 65378 25508 65390
rect 25452 65326 25454 65378
rect 25506 65326 25508 65378
rect 23548 64932 23604 64942
rect 23548 64838 23604 64876
rect 23996 64706 24052 64718
rect 23996 64654 23998 64706
rect 24050 64654 24052 64706
rect 23660 64594 23716 64606
rect 23660 64542 23662 64594
rect 23714 64542 23716 64594
rect 23212 64484 23268 64494
rect 23212 63924 23268 64428
rect 23436 63924 23492 63934
rect 23660 63924 23716 64542
rect 23996 64484 24052 64654
rect 23996 64418 24052 64428
rect 24780 64594 24836 64606
rect 24780 64542 24782 64594
rect 24834 64542 24836 64594
rect 23212 63922 23604 63924
rect 23212 63870 23438 63922
rect 23490 63870 23604 63922
rect 23212 63868 23604 63870
rect 23436 63858 23492 63868
rect 22988 63758 22990 63810
rect 23042 63758 23044 63810
rect 22988 63746 23044 63758
rect 21084 63298 21140 63308
rect 22316 63364 22372 63374
rect 22316 63270 22372 63308
rect 21308 63140 21364 63150
rect 20972 63138 21364 63140
rect 20972 63086 21310 63138
rect 21362 63086 21364 63138
rect 20972 63084 21364 63086
rect 21308 63074 21364 63084
rect 22092 62916 22148 62926
rect 20860 62412 21140 62468
rect 18172 62356 18228 62366
rect 17388 61068 18004 61124
rect 16268 60900 16324 60910
rect 16156 59892 16212 59902
rect 16156 59798 16212 59836
rect 16268 59892 16324 60844
rect 17500 60900 17556 60910
rect 17500 60806 17556 60844
rect 17948 60898 18004 61068
rect 17948 60846 17950 60898
rect 18002 60846 18004 60898
rect 17948 60834 18004 60846
rect 18060 60900 18116 60910
rect 18172 60900 18228 62300
rect 18060 60898 18228 60900
rect 18060 60846 18062 60898
rect 18114 60846 18228 60898
rect 18060 60844 18228 60846
rect 18060 60834 18116 60844
rect 17388 60786 17444 60798
rect 17388 60734 17390 60786
rect 17442 60734 17444 60786
rect 17164 60116 17220 60126
rect 17388 60116 17444 60734
rect 17724 60786 17780 60798
rect 17724 60734 17726 60786
rect 17778 60734 17780 60786
rect 17612 60228 17668 60238
rect 17612 60134 17668 60172
rect 17164 60114 17444 60116
rect 17164 60062 17166 60114
rect 17218 60062 17444 60114
rect 17164 60060 17444 60062
rect 16492 60004 16548 60014
rect 16940 60004 16996 60014
rect 16492 60002 16996 60004
rect 16492 59950 16494 60002
rect 16546 59950 16942 60002
rect 16994 59950 16996 60002
rect 16492 59948 16996 59950
rect 16492 59938 16548 59948
rect 16940 59938 16996 59948
rect 16268 59890 16436 59892
rect 16268 59838 16270 59890
rect 16322 59838 16436 59890
rect 16268 59836 16436 59838
rect 16268 59826 16324 59836
rect 15708 59442 16100 59444
rect 15708 59390 15710 59442
rect 15762 59390 16100 59442
rect 15708 59388 16100 59390
rect 16380 59444 16436 59836
rect 16716 59780 16772 59790
rect 16380 59388 16660 59444
rect 15708 59378 15764 59388
rect 15932 59218 15988 59230
rect 15932 59166 15934 59218
rect 15986 59166 15988 59218
rect 15932 58996 15988 59166
rect 16492 59218 16548 59230
rect 16492 59166 16494 59218
rect 16546 59166 16548 59218
rect 15596 58940 16436 58996
rect 14924 57698 14980 57708
rect 15036 58156 15316 58212
rect 15372 58212 15428 58222
rect 14140 56926 14142 56978
rect 14194 56926 14196 56978
rect 14140 56914 14196 56926
rect 15036 56978 15092 58156
rect 15372 58118 15428 58156
rect 15036 56926 15038 56978
rect 15090 56926 15092 56978
rect 15036 56914 15092 56926
rect 13804 56702 13806 56754
rect 13858 56702 13860 56754
rect 13804 56690 13860 56702
rect 13916 56754 13972 56766
rect 13916 56702 13918 56754
rect 13970 56702 13972 56754
rect 13692 56254 13694 56306
rect 13746 56254 13748 56306
rect 13692 56242 13748 56254
rect 13916 56644 13972 56702
rect 14252 56756 14308 56766
rect 14252 56662 14308 56700
rect 15148 56756 15204 56766
rect 15148 56662 15204 56700
rect 13132 56196 13188 56206
rect 13356 56196 13412 56206
rect 13132 56194 13356 56196
rect 13132 56142 13134 56194
rect 13186 56142 13356 56194
rect 13132 56140 13356 56142
rect 13132 56130 13188 56140
rect 13356 56102 13412 56140
rect 13468 56196 13524 56206
rect 13468 56194 13636 56196
rect 13468 56142 13470 56194
rect 13522 56142 13636 56194
rect 13468 56140 13636 56142
rect 13468 56130 13524 56140
rect 12012 53116 12628 53172
rect 12012 53058 12068 53116
rect 12012 53006 12014 53058
rect 12066 53006 12068 53058
rect 12012 52994 12068 53006
rect 12572 53058 12628 53116
rect 12572 53006 12574 53058
rect 12626 53006 12628 53058
rect 12572 52994 12628 53006
rect 12796 53228 13076 53284
rect 13132 55972 13188 55982
rect 12348 52946 12404 52958
rect 12348 52894 12350 52946
rect 12402 52894 12404 52946
rect 12348 52836 12404 52894
rect 12348 52770 12404 52780
rect 12684 52946 12740 52958
rect 12684 52894 12686 52946
rect 12738 52894 12740 52946
rect 12348 52276 12404 52286
rect 12684 52276 12740 52894
rect 12348 52274 12740 52276
rect 12348 52222 12350 52274
rect 12402 52222 12740 52274
rect 12348 52220 12740 52222
rect 12348 52210 12404 52220
rect 12236 51938 12292 51950
rect 12236 51886 12238 51938
rect 12290 51886 12292 51938
rect 12236 50708 12292 51886
rect 12460 51940 12516 51950
rect 12460 51938 12740 51940
rect 12460 51886 12462 51938
rect 12514 51886 12740 51938
rect 12460 51884 12740 51886
rect 12460 51874 12516 51884
rect 12236 50642 12292 50652
rect 12684 49812 12740 51884
rect 12684 49718 12740 49756
rect 12348 49700 12404 49710
rect 12348 49606 12404 49644
rect 12572 48244 12628 48254
rect 12460 48130 12516 48142
rect 12460 48078 12462 48130
rect 12514 48078 12516 48130
rect 12236 47460 12292 47470
rect 12236 47366 12292 47404
rect 12460 46788 12516 48078
rect 12572 47346 12628 48188
rect 12572 47294 12574 47346
rect 12626 47294 12628 47346
rect 12572 47282 12628 47294
rect 12796 47012 12852 53228
rect 12908 53060 12964 53070
rect 12908 52162 12964 53004
rect 13132 52948 13188 55916
rect 13580 55468 13636 56140
rect 13916 56194 13972 56588
rect 14028 56642 14084 56654
rect 14028 56590 14030 56642
rect 14082 56590 14084 56642
rect 14028 56420 14084 56590
rect 14700 56644 14756 56654
rect 14700 56550 14756 56588
rect 14924 56642 14980 56654
rect 14924 56590 14926 56642
rect 14978 56590 14980 56642
rect 14924 56420 14980 56590
rect 14028 56364 14980 56420
rect 13916 56142 13918 56194
rect 13970 56142 13972 56194
rect 13916 56130 13972 56142
rect 14028 56196 14084 56206
rect 14028 56102 14084 56140
rect 13468 55412 13636 55468
rect 13468 55300 13524 55412
rect 13468 55234 13524 55244
rect 13580 55076 13636 55086
rect 13580 54982 13636 55020
rect 13356 54180 13412 54190
rect 13020 52892 13188 52948
rect 13244 54124 13356 54180
rect 13020 52276 13076 52892
rect 13132 52724 13188 52734
rect 13244 52724 13300 54124
rect 13356 54114 13412 54124
rect 14140 54180 14196 56364
rect 14252 56082 14308 56094
rect 14252 56030 14254 56082
rect 14306 56030 14308 56082
rect 14252 55972 14308 56030
rect 14588 56084 14644 56094
rect 14588 55990 14644 56028
rect 15148 56082 15204 56094
rect 15148 56030 15150 56082
rect 15202 56030 15204 56082
rect 14252 55906 14308 55916
rect 15148 55468 15204 56030
rect 15260 55972 15316 55982
rect 15260 55878 15316 55916
rect 14700 55412 15204 55468
rect 14476 55300 14532 55310
rect 14476 55206 14532 55244
rect 14588 55074 14644 55086
rect 14588 55022 14590 55074
rect 14642 55022 14644 55074
rect 14588 54852 14644 55022
rect 14252 54796 14644 54852
rect 14252 54514 14308 54796
rect 14700 54740 14756 55412
rect 14588 54684 14756 54740
rect 14588 54626 14644 54684
rect 14588 54574 14590 54626
rect 14642 54574 14644 54626
rect 14588 54562 14644 54574
rect 14252 54462 14254 54514
rect 14306 54462 14308 54514
rect 14252 54450 14308 54462
rect 14476 54516 14532 54526
rect 14812 54516 14868 54526
rect 15148 54516 15204 54526
rect 14476 54422 14532 54460
rect 14700 54514 15204 54516
rect 14700 54462 14814 54514
rect 14866 54462 15150 54514
rect 15202 54462 15204 54514
rect 14700 54460 15204 54462
rect 14140 54114 14196 54124
rect 14588 53172 14644 53182
rect 14700 53172 14756 54460
rect 14812 54450 14868 54460
rect 15148 54450 15204 54460
rect 15484 54516 15540 54526
rect 15484 54422 15540 54460
rect 14588 53170 14756 53172
rect 14588 53118 14590 53170
rect 14642 53118 14756 53170
rect 14588 53116 14756 53118
rect 14588 53106 14644 53116
rect 14812 53060 14868 53070
rect 14812 52966 14868 53004
rect 14924 52946 14980 52958
rect 14924 52894 14926 52946
rect 14978 52894 14980 52946
rect 13692 52836 13748 52846
rect 13132 52722 13300 52724
rect 13132 52670 13134 52722
rect 13186 52670 13300 52722
rect 13132 52668 13300 52670
rect 13580 52834 13748 52836
rect 13580 52782 13694 52834
rect 13746 52782 13748 52834
rect 13580 52780 13748 52782
rect 13132 52658 13188 52668
rect 13020 52220 13300 52276
rect 12908 52110 12910 52162
rect 12962 52110 12964 52162
rect 12908 52052 12964 52110
rect 12908 51996 13188 52052
rect 12908 51828 12964 51838
rect 12908 51602 12964 51772
rect 12908 51550 12910 51602
rect 12962 51550 12964 51602
rect 12908 51538 12964 51550
rect 13132 51602 13188 51996
rect 13132 51550 13134 51602
rect 13186 51550 13188 51602
rect 13132 51538 13188 51550
rect 13244 50428 13300 52220
rect 13580 52164 13636 52780
rect 13692 52770 13748 52780
rect 14924 52388 14980 52894
rect 14700 52332 14980 52388
rect 13468 52162 13636 52164
rect 13468 52110 13582 52162
rect 13634 52110 13636 52162
rect 13468 52108 13636 52110
rect 13468 51828 13524 52108
rect 13580 52098 13636 52108
rect 13916 52162 13972 52174
rect 13916 52110 13918 52162
rect 13970 52110 13972 52162
rect 13356 51604 13412 51614
rect 13356 51510 13412 51548
rect 13468 51490 13524 51772
rect 13468 51438 13470 51490
rect 13522 51438 13524 51490
rect 13468 51426 13524 51438
rect 13916 51604 13972 52110
rect 13916 50428 13972 51548
rect 14476 52164 14532 52174
rect 14364 51492 14420 51502
rect 14364 50818 14420 51436
rect 14476 51380 14532 52108
rect 14588 51380 14644 51390
rect 14476 51378 14644 51380
rect 14476 51326 14590 51378
rect 14642 51326 14644 51378
rect 14476 51324 14644 51326
rect 14700 51380 14756 52332
rect 14924 52276 14980 52332
rect 14924 52210 14980 52220
rect 14812 52162 14868 52174
rect 14812 52110 14814 52162
rect 14866 52110 14868 52162
rect 14812 51604 14868 52110
rect 15036 52162 15092 52174
rect 15036 52110 15038 52162
rect 15090 52110 15092 52162
rect 15036 51716 15092 52110
rect 15260 52164 15316 52174
rect 15260 52070 15316 52108
rect 15036 51660 15316 51716
rect 14812 51548 15092 51604
rect 15036 51492 15092 51548
rect 15036 51398 15092 51436
rect 14700 51324 14868 51380
rect 14588 51314 14644 51324
rect 14812 51156 14868 51324
rect 15260 51378 15316 51660
rect 15260 51326 15262 51378
rect 15314 51326 15316 51378
rect 15148 51266 15204 51278
rect 15148 51214 15150 51266
rect 15202 51214 15204 51266
rect 15148 51156 15204 51214
rect 14812 51100 15204 51156
rect 14364 50766 14366 50818
rect 14418 50766 14420 50818
rect 14364 50754 14420 50766
rect 13132 50372 13300 50428
rect 12908 47348 12964 47358
rect 12908 47346 13076 47348
rect 12908 47294 12910 47346
rect 12962 47294 13076 47346
rect 12908 47292 13076 47294
rect 12908 47282 12964 47292
rect 12796 46956 12964 47012
rect 12572 46788 12628 46798
rect 12460 46786 12628 46788
rect 12460 46734 12574 46786
rect 12626 46734 12628 46786
rect 12460 46732 12628 46734
rect 12572 46722 12628 46732
rect 12796 46786 12852 46798
rect 12796 46734 12798 46786
rect 12850 46734 12852 46786
rect 11900 46674 12068 46676
rect 11900 46622 11902 46674
rect 11954 46622 12068 46674
rect 11900 46620 12068 46622
rect 11900 46610 11956 46620
rect 11900 46116 11956 46126
rect 11900 41860 11956 46060
rect 12012 45780 12068 46620
rect 12684 46564 12740 46574
rect 12124 46562 12740 46564
rect 12124 46510 12686 46562
rect 12738 46510 12740 46562
rect 12124 46508 12740 46510
rect 12124 46002 12180 46508
rect 12684 46498 12740 46508
rect 12796 46116 12852 46734
rect 12796 46050 12852 46060
rect 12124 45950 12126 46002
rect 12178 45950 12180 46002
rect 12124 45938 12180 45950
rect 12796 45890 12852 45902
rect 12796 45838 12798 45890
rect 12850 45838 12852 45890
rect 12012 45724 12516 45780
rect 12460 45332 12516 45724
rect 12796 45444 12852 45838
rect 12796 45378 12852 45388
rect 12460 45238 12516 45276
rect 12908 44548 12964 46956
rect 13020 46676 13076 47292
rect 13132 46900 13188 50372
rect 13692 50370 13748 50382
rect 13692 50318 13694 50370
rect 13746 50318 13748 50370
rect 13244 49812 13300 49822
rect 13244 49718 13300 49756
rect 13692 49700 13748 50318
rect 13692 49634 13748 49644
rect 13804 50372 13972 50428
rect 14028 50482 14084 50494
rect 14028 50430 14030 50482
rect 14082 50430 14084 50482
rect 13580 48354 13636 48366
rect 13580 48302 13582 48354
rect 13634 48302 13636 48354
rect 13356 48244 13412 48254
rect 13356 47908 13412 48188
rect 13356 47842 13412 47852
rect 13580 47572 13636 48302
rect 13692 48132 13748 48142
rect 13692 48038 13748 48076
rect 13468 47516 13636 47572
rect 13692 47908 13748 47918
rect 13356 47460 13412 47470
rect 13356 47366 13412 47404
rect 13132 46834 13188 46844
rect 13468 47012 13524 47516
rect 13692 47458 13748 47852
rect 13692 47406 13694 47458
rect 13746 47406 13748 47458
rect 13692 47394 13748 47406
rect 13580 47348 13636 47358
rect 13580 47254 13636 47292
rect 13132 46676 13188 46686
rect 13020 46620 13132 46676
rect 13132 46610 13188 46620
rect 13468 46674 13524 46956
rect 13468 46622 13470 46674
rect 13522 46622 13524 46674
rect 13468 46610 13524 46622
rect 13580 46004 13636 46014
rect 13580 45666 13636 45948
rect 13580 45614 13582 45666
rect 13634 45614 13636 45666
rect 13580 45444 13636 45614
rect 13580 45378 13636 45388
rect 12684 44492 12964 44548
rect 13804 44548 13860 50372
rect 13916 49700 13972 49710
rect 14028 49700 14084 50430
rect 14252 50372 14308 50382
rect 14252 50370 14420 50372
rect 14252 50318 14254 50370
rect 14306 50318 14420 50370
rect 14252 50316 14420 50318
rect 14252 50306 14308 50316
rect 13972 49644 14084 49700
rect 14364 49812 14420 50316
rect 13916 49606 13972 49644
rect 14028 47460 14084 47470
rect 14028 47366 14084 47404
rect 13916 46674 13972 46686
rect 13916 46622 13918 46674
rect 13970 46622 13972 46674
rect 13916 45220 13972 46622
rect 14028 46116 14084 46126
rect 14028 46002 14084 46060
rect 14028 45950 14030 46002
rect 14082 45950 14084 46002
rect 14028 45938 14084 45950
rect 14028 45220 14084 45230
rect 13916 45164 14028 45220
rect 14028 45154 14084 45164
rect 13804 44492 14084 44548
rect 12572 42754 12628 42766
rect 12572 42702 12574 42754
rect 12626 42702 12628 42754
rect 12348 42532 12404 42542
rect 12348 42438 12404 42476
rect 12572 42308 12628 42702
rect 12236 42252 12628 42308
rect 11900 41794 11956 41804
rect 12124 42196 12180 42206
rect 12124 41636 12180 42140
rect 11788 38222 11790 38274
rect 11842 38222 11844 38274
rect 11788 38210 11844 38222
rect 11900 41580 12180 41636
rect 12236 42084 12292 42252
rect 11004 37986 11060 37996
rect 11452 38052 11508 38062
rect 11900 38052 11956 41580
rect 12236 40626 12292 42028
rect 12684 41300 12740 44492
rect 13468 44436 13524 44446
rect 13468 44210 13524 44380
rect 13468 44158 13470 44210
rect 13522 44158 13524 44210
rect 13468 44146 13524 44158
rect 13692 44322 13748 44334
rect 13692 44270 13694 44322
rect 13746 44270 13748 44322
rect 13692 43652 13748 44270
rect 13468 43596 13748 43652
rect 13916 43650 13972 43662
rect 13916 43598 13918 43650
rect 13970 43598 13972 43650
rect 13468 43540 13524 43596
rect 13804 43540 13860 43550
rect 12908 42532 12964 42542
rect 12796 41972 12852 41982
rect 12908 41972 12964 42476
rect 13468 42196 13524 43484
rect 13692 43538 13860 43540
rect 13692 43486 13806 43538
rect 13858 43486 13860 43538
rect 13692 43484 13860 43486
rect 13468 42130 13524 42140
rect 13580 43316 13636 43326
rect 13580 42082 13636 43260
rect 13580 42030 13582 42082
rect 13634 42030 13636 42082
rect 13580 42018 13636 42030
rect 12796 41970 12964 41972
rect 12796 41918 12798 41970
rect 12850 41918 12964 41970
rect 12796 41916 12964 41918
rect 12796 41906 12852 41916
rect 12460 41244 12740 41300
rect 12348 40964 12404 40974
rect 12348 40870 12404 40908
rect 12460 40740 12516 41244
rect 12684 41076 12740 41086
rect 12684 40982 12740 41020
rect 12236 40574 12238 40626
rect 12290 40574 12292 40626
rect 12236 40562 12292 40574
rect 12348 40684 12516 40740
rect 12572 40740 12628 40750
rect 12348 40404 12404 40684
rect 12572 40628 12628 40684
rect 12460 40572 12628 40628
rect 12460 40514 12516 40572
rect 12460 40462 12462 40514
rect 12514 40462 12516 40514
rect 12460 40450 12516 40462
rect 12796 40516 12852 40526
rect 11452 38050 11732 38052
rect 11452 37998 11454 38050
rect 11506 37998 11732 38050
rect 11452 37996 11732 37998
rect 11452 37986 11508 37996
rect 10220 37266 10612 37268
rect 10220 37214 10222 37266
rect 10274 37214 10612 37266
rect 10220 37212 10612 37214
rect 10668 37660 10836 37716
rect 11228 37938 11284 37950
rect 11228 37886 11230 37938
rect 11282 37886 11284 37938
rect 10220 37156 10276 37212
rect 9996 37100 10276 37156
rect 9996 36036 10052 37100
rect 9996 35970 10052 35980
rect 10556 35924 10612 35934
rect 10332 35810 10388 35822
rect 10332 35758 10334 35810
rect 10386 35758 10388 35810
rect 9884 34862 9886 34914
rect 9938 34862 9940 34914
rect 9660 34290 9716 34300
rect 9884 34244 9940 34862
rect 9548 33966 9550 34018
rect 9602 33966 9604 34018
rect 9548 33954 9604 33966
rect 9772 34188 9940 34244
rect 10108 35698 10164 35710
rect 10108 35646 10110 35698
rect 10162 35646 10164 35698
rect 9548 33572 9604 33582
rect 9212 32116 9268 32126
rect 9100 32060 9212 32116
rect 9212 32050 9268 32060
rect 8652 31892 8708 31902
rect 8764 31892 8932 31948
rect 7420 28366 7422 28418
rect 7474 28366 7476 28418
rect 7420 28354 7476 28366
rect 7644 30770 8036 30772
rect 7644 30718 7758 30770
rect 7810 30718 8036 30770
rect 7644 30716 8036 30718
rect 8092 31778 8148 31790
rect 8092 31726 8094 31778
rect 8146 31726 8148 31778
rect 7644 28196 7700 30716
rect 7756 30706 7812 30716
rect 7756 29988 7812 29998
rect 7812 29932 7924 29988
rect 7756 29894 7812 29932
rect 7308 28140 7700 28196
rect 7756 29426 7812 29438
rect 7756 29374 7758 29426
rect 7810 29374 7812 29426
rect 7308 27412 7364 28140
rect 7756 27972 7812 29374
rect 7868 28530 7924 29932
rect 8092 29764 8148 31726
rect 8092 29698 8148 29708
rect 8204 30210 8260 30222
rect 8204 30158 8206 30210
rect 8258 30158 8260 30210
rect 7868 28478 7870 28530
rect 7922 28478 7924 28530
rect 7868 28466 7924 28478
rect 7308 27346 7364 27356
rect 7420 27916 7812 27972
rect 7420 27076 7476 27916
rect 7980 27860 8036 27870
rect 7532 27804 7980 27860
rect 7532 27746 7588 27804
rect 7980 27766 8036 27804
rect 7532 27694 7534 27746
rect 7586 27694 7588 27746
rect 7532 27682 7588 27694
rect 8204 27636 8260 30158
rect 7868 27580 8260 27636
rect 8428 30212 8484 31892
rect 8652 31798 8708 31836
rect 7868 27300 7924 27580
rect 8428 27300 8484 30156
rect 8876 31778 8932 31892
rect 8876 31726 8878 31778
rect 8930 31726 8932 31778
rect 8876 29988 8932 31726
rect 9548 30996 9604 33516
rect 9772 31892 9828 34188
rect 9884 33908 9940 33918
rect 10108 33908 10164 35646
rect 9940 33852 10164 33908
rect 10220 35364 10276 35374
rect 10220 34130 10276 35308
rect 10332 35026 10388 35758
rect 10332 34974 10334 35026
rect 10386 34974 10388 35026
rect 10332 34962 10388 34974
rect 10444 35140 10500 35150
rect 10444 34242 10500 35084
rect 10556 34916 10612 35868
rect 10668 35138 10724 37660
rect 11228 37380 11284 37886
rect 11340 37380 11396 37390
rect 11228 37324 11340 37380
rect 11340 37286 11396 37324
rect 11004 37268 11060 37278
rect 11004 36708 11060 37212
rect 11116 37044 11172 37054
rect 11116 37042 11284 37044
rect 11116 36990 11118 37042
rect 11170 36990 11284 37042
rect 11116 36988 11284 36990
rect 11116 36978 11172 36988
rect 11004 36652 11172 36708
rect 11116 36370 11172 36652
rect 11228 36484 11284 36988
rect 11452 36484 11508 36494
rect 11228 36482 11508 36484
rect 11228 36430 11454 36482
rect 11506 36430 11508 36482
rect 11228 36428 11508 36430
rect 11116 36318 11118 36370
rect 11170 36318 11172 36370
rect 10780 36260 10836 36270
rect 10780 36166 10836 36204
rect 11004 36258 11060 36270
rect 11004 36206 11006 36258
rect 11058 36206 11060 36258
rect 11004 36148 11060 36206
rect 11004 35588 11060 36092
rect 11004 35522 11060 35532
rect 10668 35086 10670 35138
rect 10722 35086 10724 35138
rect 10668 35074 10724 35086
rect 10556 34914 10724 34916
rect 10556 34862 10558 34914
rect 10610 34862 10724 34914
rect 10556 34860 10724 34862
rect 10556 34850 10612 34860
rect 10444 34190 10446 34242
rect 10498 34190 10500 34242
rect 10444 34178 10500 34190
rect 10220 34078 10222 34130
rect 10274 34078 10276 34130
rect 9884 33814 9940 33852
rect 10220 33572 10276 34078
rect 10220 33506 10276 33516
rect 10668 33348 10724 34860
rect 10780 34804 10836 34814
rect 10780 34242 10836 34748
rect 10780 34190 10782 34242
rect 10834 34190 10836 34242
rect 10780 33460 10836 34190
rect 11116 34020 11172 36318
rect 11340 35698 11396 36428
rect 11452 36418 11508 36428
rect 11340 35646 11342 35698
rect 11394 35646 11396 35698
rect 11340 35476 11396 35646
rect 11564 36372 11620 36382
rect 11564 35700 11620 36316
rect 11676 35922 11732 37996
rect 11788 37996 11956 38052
rect 12012 40348 12404 40404
rect 12572 40404 12628 40414
rect 12796 40404 12852 40460
rect 12572 40402 12852 40404
rect 12572 40350 12574 40402
rect 12626 40350 12852 40402
rect 12572 40348 12852 40350
rect 12012 38052 12068 40348
rect 12572 40338 12628 40348
rect 12796 39844 12852 39854
rect 12796 39730 12852 39788
rect 12796 39678 12798 39730
rect 12850 39678 12852 39730
rect 12796 39666 12852 39678
rect 12348 39618 12404 39630
rect 12348 39566 12350 39618
rect 12402 39566 12404 39618
rect 12124 39060 12180 39070
rect 12124 38946 12180 39004
rect 12124 38894 12126 38946
rect 12178 38894 12180 38946
rect 12124 38882 12180 38894
rect 12348 38946 12404 39566
rect 12796 39506 12852 39518
rect 12796 39454 12798 39506
rect 12850 39454 12852 39506
rect 12796 39060 12852 39454
rect 12908 39060 12964 41916
rect 13580 40740 13636 40750
rect 13580 40626 13636 40684
rect 13580 40574 13582 40626
rect 13634 40574 13636 40626
rect 13580 40562 13636 40574
rect 13356 40516 13412 40526
rect 13356 40422 13412 40460
rect 13692 40290 13748 43484
rect 13804 43474 13860 43484
rect 13804 42532 13860 42542
rect 13916 42532 13972 43598
rect 13860 42476 13972 42532
rect 13804 42438 13860 42476
rect 13916 41076 13972 41086
rect 13804 40404 13860 40414
rect 13804 40310 13860 40348
rect 13692 40238 13694 40290
rect 13746 40238 13748 40290
rect 13692 40226 13748 40238
rect 13916 40292 13972 41020
rect 13916 40226 13972 40236
rect 14028 40068 14084 44492
rect 14140 43092 14196 43102
rect 14140 42642 14196 43036
rect 14140 42590 14142 42642
rect 14194 42590 14196 42642
rect 14140 42578 14196 42590
rect 14140 41860 14196 41870
rect 14364 41860 14420 49756
rect 14812 49812 14868 49822
rect 14812 49810 15092 49812
rect 14812 49758 14814 49810
rect 14866 49758 15092 49810
rect 14812 49756 15092 49758
rect 14812 49746 14868 49756
rect 15036 49026 15092 49756
rect 15036 48974 15038 49026
rect 15090 48974 15092 49026
rect 14812 48242 14868 48254
rect 14812 48190 14814 48242
rect 14866 48190 14868 48242
rect 14812 48132 14868 48190
rect 15036 48132 15092 48974
rect 15260 48354 15316 51326
rect 15596 50428 15652 58940
rect 16156 58772 16212 58782
rect 16212 58716 16324 58772
rect 16156 58706 16212 58716
rect 15820 58324 15876 58334
rect 16156 58324 16212 58334
rect 15820 58322 16212 58324
rect 15820 58270 15822 58322
rect 15874 58270 16158 58322
rect 16210 58270 16212 58322
rect 15820 58268 16212 58270
rect 15820 58258 15876 58268
rect 16156 58212 16212 58268
rect 16156 58146 16212 58156
rect 16044 57092 16100 57102
rect 16044 56194 16100 57036
rect 16156 56980 16212 56990
rect 16268 56980 16324 58716
rect 16380 58658 16436 58940
rect 16380 58606 16382 58658
rect 16434 58606 16436 58658
rect 16380 58594 16436 58606
rect 16492 58212 16548 59166
rect 16604 58660 16660 59388
rect 16716 59442 16772 59724
rect 16716 59390 16718 59442
rect 16770 59390 16772 59442
rect 16716 59378 16772 59390
rect 17164 59444 17220 60060
rect 17164 59378 17220 59388
rect 17612 59332 17668 59342
rect 17612 59238 17668 59276
rect 17724 59218 17780 60734
rect 18060 60562 18116 60574
rect 18060 60510 18062 60562
rect 18114 60510 18116 60562
rect 18060 59892 18116 60510
rect 18060 59332 18116 59836
rect 18172 59780 18228 60844
rect 18732 60004 18788 62412
rect 18956 62374 19012 62412
rect 19180 62354 19236 62366
rect 19180 62302 19182 62354
rect 19234 62302 19236 62354
rect 19180 62132 19236 62302
rect 19516 62356 19572 62366
rect 19852 62356 19908 62366
rect 19572 62354 19908 62356
rect 19572 62302 19854 62354
rect 19906 62302 19908 62354
rect 19572 62300 19908 62302
rect 19516 62262 19572 62300
rect 19852 62290 19908 62300
rect 20076 62354 20132 62366
rect 20076 62302 20078 62354
rect 20130 62302 20132 62354
rect 20076 62132 20132 62302
rect 20412 62354 20468 62366
rect 20412 62302 20414 62354
rect 20466 62302 20468 62354
rect 20412 62244 20468 62302
rect 20412 62178 20468 62188
rect 20860 62244 20916 62254
rect 20860 62150 20916 62188
rect 19180 62076 20132 62132
rect 19180 61572 19236 62076
rect 20300 61796 20356 61806
rect 20300 61794 21028 61796
rect 20300 61742 20302 61794
rect 20354 61742 21028 61794
rect 20300 61740 21028 61742
rect 20300 61730 20356 61740
rect 18844 61516 19236 61572
rect 18844 60674 18900 61516
rect 19964 61460 20020 61470
rect 18844 60622 18846 60674
rect 18898 60622 18900 60674
rect 18844 60452 18900 60622
rect 18844 60386 18900 60396
rect 18956 61458 20020 61460
rect 18956 61406 19966 61458
rect 20018 61406 20020 61458
rect 18956 61404 20020 61406
rect 18956 60226 19012 61404
rect 19964 61394 20020 61404
rect 20412 61458 20468 61470
rect 20412 61406 20414 61458
rect 20466 61406 20468 61458
rect 20188 61348 20244 61358
rect 20412 61348 20468 61406
rect 20188 61346 20468 61348
rect 20188 61294 20190 61346
rect 20242 61294 20468 61346
rect 20188 61292 20468 61294
rect 20636 61458 20692 61470
rect 20636 61406 20638 61458
rect 20690 61406 20692 61458
rect 20636 61348 20692 61406
rect 20748 61348 20804 61358
rect 20636 61346 20804 61348
rect 20636 61294 20750 61346
rect 20802 61294 20804 61346
rect 20636 61292 20804 61294
rect 20188 61282 20244 61292
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 18956 60174 18958 60226
rect 19010 60174 19012 60226
rect 18956 60162 19012 60174
rect 20188 60452 20244 60462
rect 18844 60004 18900 60014
rect 18732 60002 18900 60004
rect 18732 59950 18846 60002
rect 18898 59950 18900 60002
rect 18732 59948 18900 59950
rect 18844 59938 18900 59948
rect 19852 60002 19908 60014
rect 19852 59950 19854 60002
rect 19906 59950 19908 60002
rect 18172 59714 18228 59724
rect 19852 59780 19908 59950
rect 20188 60002 20244 60396
rect 20188 59950 20190 60002
rect 20242 59950 20244 60002
rect 20188 59938 20244 59950
rect 19852 59714 19908 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 18060 59266 18116 59276
rect 17724 59166 17726 59218
rect 17778 59166 17780 59218
rect 17724 59154 17780 59166
rect 18060 59108 18116 59118
rect 18060 59014 18116 59052
rect 20300 58996 20356 61292
rect 20748 61282 20804 61292
rect 20972 60898 21028 61740
rect 20972 60846 20974 60898
rect 21026 60846 21028 60898
rect 20972 60834 21028 60846
rect 21084 60676 21140 62412
rect 20300 58930 20356 58940
rect 20524 60620 21140 60676
rect 21756 61570 21812 61582
rect 21756 61518 21758 61570
rect 21810 61518 21812 61570
rect 21756 60786 21812 61518
rect 21756 60734 21758 60786
rect 21810 60734 21812 60786
rect 21756 60676 21812 60734
rect 16716 58660 16772 58670
rect 16604 58658 16772 58660
rect 16604 58606 16718 58658
rect 16770 58606 16772 58658
rect 16604 58604 16772 58606
rect 16716 58594 16772 58604
rect 16492 58146 16548 58156
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19740 57876 19796 57886
rect 16604 57764 16660 57774
rect 19628 57764 19684 57774
rect 16156 56978 16548 56980
rect 16156 56926 16158 56978
rect 16210 56926 16548 56978
rect 16156 56924 16548 56926
rect 16156 56914 16212 56924
rect 16492 56866 16548 56924
rect 16492 56814 16494 56866
rect 16546 56814 16548 56866
rect 16492 56802 16548 56814
rect 16044 56142 16046 56194
rect 16098 56142 16100 56194
rect 16044 56130 16100 56142
rect 16492 52500 16548 52510
rect 15708 52388 15764 52398
rect 16156 52388 16212 52398
rect 15708 52386 16212 52388
rect 15708 52334 15710 52386
rect 15762 52334 16158 52386
rect 16210 52334 16212 52386
rect 15708 52332 16212 52334
rect 15708 52322 15764 52332
rect 16156 52322 16212 52332
rect 16492 52386 16548 52444
rect 16492 52334 16494 52386
rect 16546 52334 16548 52386
rect 16492 52322 16548 52334
rect 15932 52164 15988 52174
rect 15932 52070 15988 52108
rect 16604 50428 16660 57708
rect 19516 57762 19684 57764
rect 19516 57710 19630 57762
rect 19682 57710 19684 57762
rect 19516 57708 19684 57710
rect 19404 57652 19460 57662
rect 19404 57558 19460 57596
rect 19068 57540 19124 57550
rect 17276 56756 17332 56766
rect 17276 56754 17892 56756
rect 17276 56702 17278 56754
rect 17330 56702 17892 56754
rect 17276 56700 17892 56702
rect 17276 56690 17332 56700
rect 17836 55970 17892 56700
rect 17836 55918 17838 55970
rect 17890 55918 17892 55970
rect 17836 55906 17892 55918
rect 17948 56194 18004 56206
rect 17948 56142 17950 56194
rect 18002 56142 18004 56194
rect 17948 55468 18004 56142
rect 19068 56194 19124 57484
rect 19516 57092 19572 57708
rect 19628 57698 19684 57708
rect 19740 57762 19796 57820
rect 20300 57876 20356 57886
rect 20356 57820 20468 57876
rect 20300 57810 20356 57820
rect 19740 57710 19742 57762
rect 19794 57710 19796 57762
rect 19740 57698 19796 57710
rect 20076 57650 20132 57662
rect 20076 57598 20078 57650
rect 20130 57598 20132 57650
rect 19516 57036 20020 57092
rect 19404 56980 19460 56990
rect 19516 56980 19572 57036
rect 19404 56978 19572 56980
rect 19404 56926 19406 56978
rect 19458 56926 19572 56978
rect 19404 56924 19572 56926
rect 19404 56914 19460 56924
rect 19852 56868 19908 56878
rect 19852 56756 19908 56812
rect 19068 56142 19070 56194
rect 19122 56142 19124 56194
rect 19068 56130 19124 56142
rect 19628 56754 19908 56756
rect 19628 56702 19854 56754
rect 19906 56702 19908 56754
rect 19628 56700 19908 56702
rect 18172 55972 18228 55982
rect 18732 55972 18788 55982
rect 18172 55970 18788 55972
rect 18172 55918 18174 55970
rect 18226 55918 18734 55970
rect 18786 55918 18788 55970
rect 18172 55916 18788 55918
rect 18172 55906 18228 55916
rect 18732 55906 18788 55916
rect 17948 55412 18116 55468
rect 16940 55076 16996 55086
rect 16716 54404 16772 54414
rect 16716 54310 16772 54348
rect 15260 48302 15262 48354
rect 15314 48302 15316 48354
rect 15260 48290 15316 48302
rect 15372 50372 15652 50428
rect 16492 50372 16660 50428
rect 15148 48132 15204 48142
rect 15036 48130 15204 48132
rect 15036 48078 15150 48130
rect 15202 48078 15204 48130
rect 15036 48076 15204 48078
rect 14812 48066 14868 48076
rect 15148 48066 15204 48076
rect 15260 47572 15316 47582
rect 15148 47516 15260 47572
rect 14588 47236 14644 47246
rect 14588 47234 14756 47236
rect 14588 47182 14590 47234
rect 14642 47182 14756 47234
rect 14588 47180 14756 47182
rect 14588 47170 14644 47180
rect 14700 47124 14756 47180
rect 14476 46676 14532 46686
rect 14532 46620 14644 46676
rect 14476 46582 14532 46620
rect 14476 45330 14532 45342
rect 14476 45278 14478 45330
rect 14530 45278 14532 45330
rect 14476 45220 14532 45278
rect 14476 45154 14532 45164
rect 14588 45106 14644 46620
rect 14588 45054 14590 45106
rect 14642 45054 14644 45106
rect 14588 42868 14644 45054
rect 14700 43762 14756 47068
rect 14812 46674 14868 46686
rect 14812 46622 14814 46674
rect 14866 46622 14868 46674
rect 14812 45892 14868 46622
rect 14812 45836 14980 45892
rect 14812 45668 14868 45678
rect 14812 45574 14868 45612
rect 14812 45220 14868 45230
rect 14924 45220 14980 45836
rect 14868 45164 14980 45220
rect 15036 45890 15092 45902
rect 15036 45838 15038 45890
rect 15090 45838 15092 45890
rect 14812 45154 14868 45164
rect 15036 45108 15092 45838
rect 15036 45042 15092 45052
rect 15148 44322 15204 47516
rect 15260 47506 15316 47516
rect 15372 45668 15428 50372
rect 16268 49252 16324 49262
rect 16268 49138 16324 49196
rect 16268 49086 16270 49138
rect 16322 49086 16324 49138
rect 16268 49074 16324 49086
rect 15596 49028 15652 49038
rect 15596 49026 16212 49028
rect 15596 48974 15598 49026
rect 15650 48974 16212 49026
rect 15596 48972 16212 48974
rect 15596 48962 15652 48972
rect 15708 48354 15764 48366
rect 15708 48302 15710 48354
rect 15762 48302 15764 48354
rect 15484 47348 15540 47358
rect 15708 47348 15764 48302
rect 15932 48242 15988 48254
rect 15932 48190 15934 48242
rect 15986 48190 15988 48242
rect 15484 47346 15764 47348
rect 15484 47294 15486 47346
rect 15538 47294 15764 47346
rect 15484 47292 15764 47294
rect 15820 47458 15876 47470
rect 15820 47406 15822 47458
rect 15874 47406 15876 47458
rect 15484 47282 15540 47292
rect 15820 47124 15876 47406
rect 15932 47348 15988 48190
rect 16156 48132 16212 48972
rect 16156 48076 16324 48132
rect 16268 47570 16324 48076
rect 16268 47518 16270 47570
rect 16322 47518 16324 47570
rect 16268 47506 16324 47518
rect 16492 47572 16548 50372
rect 16716 49140 16772 49150
rect 16716 49026 16772 49084
rect 16716 48974 16718 49026
rect 16770 48974 16772 49026
rect 16716 48962 16772 48974
rect 16492 47506 16548 47516
rect 16604 48132 16660 48142
rect 16044 47458 16100 47470
rect 16044 47406 16046 47458
rect 16098 47406 16100 47458
rect 16044 47348 16100 47406
rect 16380 47460 16436 47470
rect 16380 47366 16436 47404
rect 16604 47458 16660 48076
rect 16604 47406 16606 47458
rect 16658 47406 16660 47458
rect 16604 47394 16660 47406
rect 15932 47292 16100 47348
rect 15820 47058 15876 47068
rect 15932 46564 15988 46574
rect 15932 46470 15988 46508
rect 16044 46340 16100 47292
rect 15708 46284 16100 46340
rect 15484 45780 15540 45790
rect 15484 45686 15540 45724
rect 15372 45602 15428 45612
rect 15596 45666 15652 45678
rect 15596 45614 15598 45666
rect 15650 45614 15652 45666
rect 15372 45220 15428 45230
rect 15596 45220 15652 45614
rect 15372 45218 15652 45220
rect 15372 45166 15374 45218
rect 15426 45166 15652 45218
rect 15372 45164 15652 45166
rect 15372 44436 15428 45164
rect 15708 44994 15764 46284
rect 15820 45892 15876 45902
rect 15820 45798 15876 45836
rect 15820 45668 15876 45678
rect 15876 45612 15988 45668
rect 15820 45602 15876 45612
rect 15708 44942 15710 44994
rect 15762 44942 15764 44994
rect 15708 44930 15764 44942
rect 15820 45108 15876 45118
rect 15372 44370 15428 44380
rect 15820 44436 15876 45052
rect 15820 44370 15876 44380
rect 15148 44270 15150 44322
rect 15202 44270 15204 44322
rect 15148 44258 15204 44270
rect 15484 44212 15540 44222
rect 15484 44210 15652 44212
rect 15484 44158 15486 44210
rect 15538 44158 15652 44210
rect 15484 44156 15652 44158
rect 15484 44146 15540 44156
rect 14700 43710 14702 43762
rect 14754 43710 14756 43762
rect 14700 43698 14756 43710
rect 15372 44098 15428 44110
rect 15372 44046 15374 44098
rect 15426 44046 15428 44098
rect 14812 43538 14868 43550
rect 14812 43486 14814 43538
rect 14866 43486 14868 43538
rect 14700 42868 14756 42878
rect 14588 42812 14700 42868
rect 14700 42802 14756 42812
rect 14700 42084 14756 42094
rect 14700 41970 14756 42028
rect 14700 41918 14702 41970
rect 14754 41918 14756 41970
rect 14700 41906 14756 41918
rect 14140 40180 14196 41804
rect 14252 41804 14420 41860
rect 14588 41860 14644 41870
rect 14252 40628 14308 41804
rect 14588 41766 14644 41804
rect 14476 41748 14532 41758
rect 14252 40562 14308 40572
rect 14364 41692 14476 41748
rect 14364 40516 14420 41692
rect 14476 41682 14532 41692
rect 14588 40964 14644 40974
rect 14364 40422 14420 40460
rect 14476 40908 14588 40964
rect 14252 40404 14308 40414
rect 14252 40310 14308 40348
rect 14364 40292 14420 40302
rect 14140 40124 14308 40180
rect 13692 40012 14084 40068
rect 13468 39394 13524 39406
rect 13468 39342 13470 39394
rect 13522 39342 13524 39394
rect 13132 39060 13188 39070
rect 12908 39058 13188 39060
rect 12908 39006 13134 39058
rect 13186 39006 13188 39058
rect 12908 39004 13188 39006
rect 12348 38894 12350 38946
rect 12402 38894 12404 38946
rect 12236 38836 12292 38846
rect 12236 38274 12292 38780
rect 12348 38612 12404 38894
rect 12684 38948 12740 38958
rect 12460 38836 12516 38846
rect 12460 38742 12516 38780
rect 12684 38834 12740 38892
rect 12684 38782 12686 38834
rect 12738 38782 12740 38834
rect 12404 38556 12628 38612
rect 12348 38546 12404 38556
rect 12236 38222 12238 38274
rect 12290 38222 12292 38274
rect 12236 38210 12292 38222
rect 12572 38274 12628 38556
rect 12572 38222 12574 38274
rect 12626 38222 12628 38274
rect 12572 38210 12628 38222
rect 12012 37996 12628 38052
rect 11788 36596 11844 37996
rect 12572 37490 12628 37996
rect 12572 37438 12574 37490
rect 12626 37438 12628 37490
rect 12572 37426 12628 37438
rect 12236 37378 12292 37390
rect 12236 37326 12238 37378
rect 12290 37326 12292 37378
rect 11900 37268 11956 37278
rect 11900 37174 11956 37212
rect 11900 36596 11956 36606
rect 11788 36594 11956 36596
rect 11788 36542 11902 36594
rect 11954 36542 11956 36594
rect 11788 36540 11956 36542
rect 11900 36530 11956 36540
rect 12236 36372 12292 37326
rect 12460 37380 12516 37390
rect 12460 37286 12516 37324
rect 12684 37268 12740 38782
rect 12796 38724 12852 39004
rect 13132 38994 13188 39004
rect 12796 38162 12852 38668
rect 13468 38724 13524 39342
rect 13468 38658 13524 38668
rect 13692 38274 13748 40012
rect 14140 39620 14196 39630
rect 13804 39618 14196 39620
rect 13804 39566 14142 39618
rect 14194 39566 14196 39618
rect 13804 39564 14196 39566
rect 13804 39506 13860 39564
rect 14140 39554 14196 39564
rect 14252 39620 14308 40124
rect 14252 39554 14308 39564
rect 13804 39454 13806 39506
rect 13858 39454 13860 39506
rect 13804 39442 13860 39454
rect 13692 38222 13694 38274
rect 13746 38222 13748 38274
rect 13692 38210 13748 38222
rect 14140 38948 14196 38958
rect 12796 38110 12798 38162
rect 12850 38110 12852 38162
rect 12796 38098 12852 38110
rect 14028 38050 14084 38062
rect 14028 37998 14030 38050
rect 14082 37998 14084 38050
rect 14028 37716 14084 37998
rect 14028 37650 14084 37660
rect 14140 37490 14196 38892
rect 14364 38668 14420 40236
rect 14476 40180 14532 40908
rect 14588 40870 14644 40908
rect 14812 40740 14868 43486
rect 15036 42756 15092 42766
rect 15036 42082 15092 42700
rect 15372 42420 15428 44046
rect 15484 43540 15540 43550
rect 15484 43446 15540 43484
rect 15596 43316 15652 44156
rect 15484 43260 15652 43316
rect 15484 42756 15540 43260
rect 15932 42978 15988 45612
rect 16156 44436 16212 44446
rect 16156 44342 16212 44380
rect 16380 43876 16436 43886
rect 16380 43650 16436 43820
rect 16380 43598 16382 43650
rect 16434 43598 16436 43650
rect 16380 43586 16436 43598
rect 16156 43428 16212 43438
rect 16156 43334 16212 43372
rect 15932 42926 15934 42978
rect 15986 42926 15988 42978
rect 15932 42914 15988 42926
rect 16156 42980 16212 42990
rect 15484 42690 15540 42700
rect 15596 42644 15652 42654
rect 15596 42642 15764 42644
rect 15596 42590 15598 42642
rect 15650 42590 15764 42642
rect 15596 42588 15764 42590
rect 15596 42578 15652 42588
rect 15372 42364 15540 42420
rect 15036 42030 15038 42082
rect 15090 42030 15092 42082
rect 15036 42018 15092 42030
rect 15148 42084 15204 42094
rect 14588 40684 14868 40740
rect 15148 41186 15204 42028
rect 15372 41970 15428 41982
rect 15372 41918 15374 41970
rect 15426 41918 15428 41970
rect 15260 41748 15316 41758
rect 15260 41654 15316 41692
rect 15372 41636 15428 41918
rect 15484 41860 15540 42364
rect 15596 42084 15652 42094
rect 15596 41990 15652 42028
rect 15596 41860 15652 41870
rect 15484 41804 15596 41860
rect 15596 41794 15652 41804
rect 15372 41570 15428 41580
rect 15148 41134 15150 41186
rect 15202 41134 15204 41186
rect 14588 40626 14644 40684
rect 14588 40574 14590 40626
rect 14642 40574 14644 40626
rect 14588 40562 14644 40574
rect 14924 40628 14980 40638
rect 15148 40628 15204 41134
rect 14980 40572 15092 40628
rect 14924 40562 14980 40572
rect 14812 40404 14868 40414
rect 14812 40310 14868 40348
rect 14476 40124 14980 40180
rect 14588 39956 14644 39966
rect 14588 39730 14644 39900
rect 14588 39678 14590 39730
rect 14642 39678 14644 39730
rect 14588 39666 14644 39678
rect 14812 39956 14868 39966
rect 14812 39730 14868 39900
rect 14812 39678 14814 39730
rect 14866 39678 14868 39730
rect 14812 39666 14868 39678
rect 14924 39618 14980 40124
rect 14924 39566 14926 39618
rect 14978 39566 14980 39618
rect 14924 39554 14980 39566
rect 15036 38668 15092 40572
rect 15148 40562 15204 40572
rect 15708 41186 15764 42588
rect 15820 42532 15876 42542
rect 15820 42438 15876 42476
rect 15708 41134 15710 41186
rect 15762 41134 15764 41186
rect 15708 40964 15764 41134
rect 15148 40404 15204 40414
rect 15148 40402 15316 40404
rect 15148 40350 15150 40402
rect 15202 40350 15316 40402
rect 15148 40348 15316 40350
rect 15148 40338 15204 40348
rect 14140 37438 14142 37490
rect 14194 37438 14196 37490
rect 14140 37426 14196 37438
rect 14252 38612 14420 38668
rect 14924 38612 15092 38668
rect 15148 39620 15204 39630
rect 14252 37268 14308 38612
rect 14812 38050 14868 38062
rect 14812 37998 14814 38050
rect 14866 37998 14868 38050
rect 14700 37940 14756 37950
rect 14476 37884 14700 37940
rect 12236 36306 12292 36316
rect 12572 37212 12740 37268
rect 14140 37212 14308 37268
rect 14364 37378 14420 37390
rect 14364 37326 14366 37378
rect 14418 37326 14420 37378
rect 12572 36036 12628 37212
rect 12796 36484 12852 36494
rect 13468 36484 13524 36494
rect 12852 36428 12964 36484
rect 12796 36390 12852 36428
rect 12684 36260 12740 36270
rect 12684 36166 12740 36204
rect 12572 35980 12740 36036
rect 11676 35870 11678 35922
rect 11730 35870 11732 35922
rect 11676 35858 11732 35870
rect 11676 35700 11732 35710
rect 11564 35698 11732 35700
rect 11564 35646 11678 35698
rect 11730 35646 11732 35698
rect 11564 35644 11732 35646
rect 11676 35634 11732 35644
rect 12012 35700 12068 35710
rect 12012 35698 12292 35700
rect 12012 35646 12014 35698
rect 12066 35646 12292 35698
rect 12012 35644 12292 35646
rect 12012 35634 12068 35644
rect 11340 35410 11396 35420
rect 12236 35140 12292 35644
rect 12348 35698 12404 35710
rect 12348 35646 12350 35698
rect 12402 35646 12404 35698
rect 12348 35364 12404 35646
rect 12572 35700 12628 35710
rect 12572 35606 12628 35644
rect 12348 35298 12404 35308
rect 12236 35084 12628 35140
rect 12572 34802 12628 35084
rect 12572 34750 12574 34802
rect 12626 34750 12628 34802
rect 12572 34738 12628 34750
rect 11452 34020 11508 34030
rect 11116 34018 11508 34020
rect 11116 33966 11454 34018
rect 11506 33966 11508 34018
rect 11116 33964 11508 33966
rect 10892 33460 10948 33470
rect 10780 33458 10948 33460
rect 10780 33406 10894 33458
rect 10946 33406 10948 33458
rect 10780 33404 10948 33406
rect 10668 33292 10836 33348
rect 10668 32786 10724 32798
rect 10668 32734 10670 32786
rect 10722 32734 10724 32786
rect 10332 32564 10388 32574
rect 10332 32470 10388 32508
rect 10556 32450 10612 32462
rect 10556 32398 10558 32450
rect 10610 32398 10612 32450
rect 9772 31826 9828 31836
rect 10444 32116 10500 32126
rect 9996 30996 10052 31006
rect 9548 30994 10052 30996
rect 9548 30942 9998 30994
rect 10050 30942 10052 30994
rect 9548 30940 10052 30942
rect 9660 30212 9716 30222
rect 9660 30210 9828 30212
rect 9660 30158 9662 30210
rect 9714 30158 9828 30210
rect 9660 30156 9828 30158
rect 9660 30146 9716 30156
rect 8876 29922 8932 29932
rect 9660 29988 9716 29998
rect 9660 29894 9716 29932
rect 9324 29876 9380 29886
rect 9100 29540 9156 29550
rect 8540 29314 8596 29326
rect 8540 29262 8542 29314
rect 8594 29262 8596 29314
rect 8540 27636 8596 29262
rect 9100 28756 9156 29484
rect 8652 28754 9156 28756
rect 8652 28702 9102 28754
rect 9154 28702 9156 28754
rect 8652 28700 9156 28702
rect 8652 28082 8708 28700
rect 9100 28690 9156 28700
rect 8652 28030 8654 28082
rect 8706 28030 8708 28082
rect 8652 28018 8708 28030
rect 8652 27636 8708 27646
rect 8540 27580 8652 27636
rect 8652 27570 8708 27580
rect 8540 27300 8596 27310
rect 8428 27298 8596 27300
rect 8428 27246 8542 27298
rect 8594 27246 8596 27298
rect 8428 27244 8596 27246
rect 7868 27206 7924 27244
rect 8540 27234 8596 27244
rect 7420 27010 7476 27020
rect 9324 27074 9380 29820
rect 9772 29540 9828 30156
rect 9772 29446 9828 29484
rect 9548 29428 9604 29438
rect 9548 29334 9604 29372
rect 9660 28644 9716 28654
rect 9324 27022 9326 27074
rect 9378 27022 9380 27074
rect 9324 27010 9380 27022
rect 9548 28196 9604 28206
rect 9548 27860 9604 28140
rect 6972 26962 7140 26964
rect 6972 26910 6974 26962
rect 7026 26910 7140 26962
rect 6972 26908 7140 26910
rect 6972 26898 7028 26908
rect 7084 26852 7140 26908
rect 7084 26786 7140 26796
rect 7868 26852 7924 26862
rect 7924 26796 8036 26852
rect 7868 26786 7924 26796
rect 7868 26178 7924 26190
rect 7868 26126 7870 26178
rect 7922 26126 7924 26178
rect 7644 25508 7700 25518
rect 7644 25414 7700 25452
rect 7868 25282 7924 26126
rect 7980 25506 8036 26796
rect 9548 26514 9604 27804
rect 9548 26462 9550 26514
rect 9602 26462 9604 26514
rect 9548 26450 9604 26462
rect 9660 27746 9716 28588
rect 9660 27694 9662 27746
rect 9714 27694 9716 27746
rect 8764 26290 8820 26302
rect 8764 26238 8766 26290
rect 8818 26238 8820 26290
rect 7980 25454 7982 25506
rect 8034 25454 8036 25506
rect 7980 25442 8036 25454
rect 8204 26180 8260 26190
rect 8204 25506 8260 26124
rect 8204 25454 8206 25506
rect 8258 25454 8260 25506
rect 8204 25442 8260 25454
rect 8652 25508 8708 25518
rect 8764 25508 8820 26238
rect 8652 25506 8820 25508
rect 8652 25454 8654 25506
rect 8706 25454 8820 25506
rect 8652 25452 8820 25454
rect 8652 25442 8708 25452
rect 7868 25230 7870 25282
rect 7922 25230 7924 25282
rect 7868 25218 7924 25230
rect 8428 25284 8484 25294
rect 8428 24946 8484 25228
rect 8764 25172 8820 25452
rect 9324 25396 9380 25406
rect 9324 25302 9380 25340
rect 8876 25172 8932 25182
rect 8764 25116 8876 25172
rect 8428 24894 8430 24946
rect 8482 24894 8484 24946
rect 8428 24882 8484 24894
rect 8876 24946 8932 25116
rect 9660 25172 9716 27694
rect 9884 27860 9940 27870
rect 9884 26180 9940 27804
rect 9996 27636 10052 30940
rect 10108 30100 10164 30110
rect 10108 30006 10164 30044
rect 10444 29650 10500 32060
rect 10444 29598 10446 29650
rect 10498 29598 10500 29650
rect 10444 29586 10500 29598
rect 10556 30100 10612 32398
rect 10668 31778 10724 32734
rect 10668 31726 10670 31778
rect 10722 31726 10724 31778
rect 10668 31714 10724 31726
rect 10556 29426 10612 30044
rect 10556 29374 10558 29426
rect 10610 29374 10612 29426
rect 10556 29362 10612 29374
rect 10780 29764 10836 33292
rect 10892 29876 10948 33404
rect 11228 33346 11284 33358
rect 11228 33294 11230 33346
rect 11282 33294 11284 33346
rect 11228 30884 11284 33294
rect 11452 33236 11508 33964
rect 12460 33460 12516 33470
rect 11452 33170 11508 33180
rect 11676 33346 11732 33358
rect 11676 33294 11678 33346
rect 11730 33294 11732 33346
rect 11564 32562 11620 32574
rect 11564 32510 11566 32562
rect 11618 32510 11620 32562
rect 11564 32452 11620 32510
rect 11564 32386 11620 32396
rect 11676 31948 11732 33294
rect 12236 33346 12292 33358
rect 12236 33294 12238 33346
rect 12290 33294 12292 33346
rect 11900 32788 11956 32798
rect 11900 32694 11956 32732
rect 12236 32452 12292 33294
rect 12236 32386 12292 32396
rect 11340 31892 11732 31948
rect 12012 32228 12068 32238
rect 11340 31778 11396 31892
rect 11340 31726 11342 31778
rect 11394 31726 11396 31778
rect 11340 31714 11396 31726
rect 11340 30884 11396 30894
rect 11228 30828 11340 30884
rect 11340 30324 11396 30828
rect 11564 30770 11620 31892
rect 11788 30996 11844 31006
rect 11564 30718 11566 30770
rect 11618 30718 11620 30770
rect 11564 30706 11620 30718
rect 11676 30994 11844 30996
rect 11676 30942 11790 30994
rect 11842 30942 11844 30994
rect 11676 30940 11844 30942
rect 10892 29810 10948 29820
rect 11228 30322 11396 30324
rect 11228 30270 11342 30322
rect 11394 30270 11396 30322
rect 11228 30268 11396 30270
rect 10780 29428 10836 29708
rect 10780 29362 10836 29372
rect 11116 29540 11172 29550
rect 11004 29314 11060 29326
rect 11004 29262 11006 29314
rect 11058 29262 11060 29314
rect 11004 28196 11060 29262
rect 11116 28754 11172 29484
rect 11116 28702 11118 28754
rect 11170 28702 11172 28754
rect 11116 28690 11172 28702
rect 11004 28130 11060 28140
rect 11004 27972 11060 27982
rect 10108 27636 10164 27646
rect 9996 27580 10108 27636
rect 10108 26962 10164 27580
rect 11004 27412 11060 27916
rect 11004 27074 11060 27356
rect 11004 27022 11006 27074
rect 11058 27022 11060 27074
rect 11004 27010 11060 27022
rect 10108 26910 10110 26962
rect 10162 26910 10164 26962
rect 10108 26898 10164 26910
rect 10668 26852 10724 26862
rect 10668 26514 10724 26796
rect 11228 26852 11284 30268
rect 11340 30258 11396 30268
rect 11564 29876 11620 29886
rect 11676 29876 11732 30940
rect 11788 30930 11844 30940
rect 11620 29820 11732 29876
rect 11564 29810 11620 29820
rect 11340 29652 11396 29662
rect 11340 29538 11396 29596
rect 11340 29486 11342 29538
rect 11394 29486 11396 29538
rect 11340 29474 11396 29486
rect 11452 29540 11508 29550
rect 11452 27970 11508 29484
rect 11452 27918 11454 27970
rect 11506 27918 11508 27970
rect 11452 27906 11508 27918
rect 12012 27636 12068 32172
rect 12460 31890 12516 33404
rect 12684 33458 12740 35980
rect 12908 35922 12964 36428
rect 13468 36390 13524 36428
rect 12908 35870 12910 35922
rect 12962 35870 12964 35922
rect 12908 35858 12964 35870
rect 13580 36258 13636 36270
rect 13804 36260 13860 36270
rect 13580 36206 13582 36258
rect 13634 36206 13636 36258
rect 13580 35924 13636 36206
rect 13580 35858 13636 35868
rect 13692 36258 13860 36260
rect 13692 36206 13806 36258
rect 13858 36206 13860 36258
rect 13692 36204 13860 36206
rect 12796 35810 12852 35822
rect 12796 35758 12798 35810
rect 12850 35758 12852 35810
rect 12796 35140 12852 35758
rect 13580 35588 13636 35598
rect 13580 35494 13636 35532
rect 12796 35074 12852 35084
rect 12684 33406 12686 33458
rect 12738 33406 12740 33458
rect 12684 33394 12740 33406
rect 12796 34914 12852 34926
rect 12796 34862 12798 34914
rect 12850 34862 12852 34914
rect 12796 33348 12852 34862
rect 12796 32788 12852 33292
rect 13020 33572 13076 33582
rect 13020 33348 13076 33516
rect 13020 33346 13300 33348
rect 13020 33294 13022 33346
rect 13074 33294 13300 33346
rect 13020 33292 13300 33294
rect 13020 33282 13076 33292
rect 12796 32722 12852 32732
rect 12460 31838 12462 31890
rect 12514 31838 12516 31890
rect 12460 31826 12516 31838
rect 12796 32562 12852 32574
rect 12796 32510 12798 32562
rect 12850 32510 12852 32562
rect 12796 31892 12852 32510
rect 12796 31826 12852 31836
rect 13132 32450 13188 32462
rect 13132 32398 13134 32450
rect 13186 32398 13188 32450
rect 12124 31778 12180 31790
rect 12124 31726 12126 31778
rect 12178 31726 12180 31778
rect 12124 29316 12180 31726
rect 12348 31778 12404 31790
rect 12348 31726 12350 31778
rect 12402 31726 12404 31778
rect 12348 31668 12404 31726
rect 13132 31668 13188 32398
rect 13244 31780 13300 33292
rect 13468 33236 13524 33246
rect 13244 31724 13412 31780
rect 12348 31612 13188 31668
rect 12908 30996 12964 31006
rect 12236 30884 12292 30894
rect 12236 30882 12404 30884
rect 12236 30830 12238 30882
rect 12290 30830 12404 30882
rect 12236 30828 12404 30830
rect 12236 30818 12292 30828
rect 12348 29652 12404 30828
rect 12348 29538 12404 29596
rect 12348 29486 12350 29538
rect 12402 29486 12404 29538
rect 12348 29474 12404 29486
rect 12124 29250 12180 29260
rect 12796 29316 12852 29326
rect 12348 29092 12404 29102
rect 12348 28532 12404 29036
rect 12236 28530 12404 28532
rect 12236 28478 12350 28530
rect 12402 28478 12404 28530
rect 12236 28476 12404 28478
rect 11676 27580 12068 27636
rect 12124 27858 12180 27870
rect 12124 27806 12126 27858
rect 12178 27806 12180 27858
rect 11564 27300 11620 27310
rect 11564 27074 11620 27244
rect 11564 27022 11566 27074
rect 11618 27022 11620 27074
rect 11564 27010 11620 27022
rect 11228 26786 11284 26796
rect 11564 26516 11620 26526
rect 11676 26516 11732 27580
rect 12124 27524 12180 27806
rect 12012 27468 12180 27524
rect 12012 27188 12068 27468
rect 10668 26462 10670 26514
rect 10722 26462 10724 26514
rect 10668 26450 10724 26462
rect 11116 26514 11732 26516
rect 11116 26462 11566 26514
rect 11618 26462 11732 26514
rect 11116 26460 11732 26462
rect 11788 26852 11844 26862
rect 11788 26514 11844 26796
rect 11788 26462 11790 26514
rect 11842 26462 11844 26514
rect 10444 26290 10500 26302
rect 10444 26238 10446 26290
rect 10498 26238 10500 26290
rect 9996 26180 10052 26190
rect 9884 26178 10052 26180
rect 9884 26126 9998 26178
rect 10050 26126 10052 26178
rect 9884 26124 10052 26126
rect 9996 26114 10052 26124
rect 10444 25284 10500 26238
rect 11116 26290 11172 26460
rect 11564 26450 11620 26460
rect 11116 26238 11118 26290
rect 11170 26238 11172 26290
rect 11116 26226 11172 26238
rect 10556 26180 10612 26190
rect 11788 26180 11844 26462
rect 10556 26086 10612 26124
rect 11564 26124 11844 26180
rect 11564 25618 11620 26124
rect 11564 25566 11566 25618
rect 11618 25566 11620 25618
rect 11564 25554 11620 25566
rect 12012 25284 12068 27132
rect 12236 27186 12292 28476
rect 12348 28466 12404 28476
rect 12796 28418 12852 29260
rect 12908 28642 12964 30940
rect 13132 29428 13188 31612
rect 13356 31556 13412 31724
rect 13468 31778 13524 33180
rect 13692 33124 13748 36204
rect 13804 36194 13860 36204
rect 13916 35698 13972 35710
rect 13916 35646 13918 35698
rect 13970 35646 13972 35698
rect 13804 35588 13860 35598
rect 13804 33346 13860 35532
rect 13916 33572 13972 35646
rect 13916 33506 13972 33516
rect 14140 33458 14196 37212
rect 14364 35588 14420 37326
rect 14476 37378 14532 37884
rect 14700 37846 14756 37884
rect 14476 37326 14478 37378
rect 14530 37326 14532 37378
rect 14476 37314 14532 37326
rect 14812 37378 14868 37998
rect 14924 37828 14980 38612
rect 15036 37828 15092 37838
rect 14924 37772 15036 37828
rect 14812 37326 14814 37378
rect 14866 37326 14868 37378
rect 14812 37314 14868 37326
rect 14924 37268 14980 37278
rect 14924 37174 14980 37212
rect 15036 35810 15092 37772
rect 15148 37044 15204 39564
rect 15260 38948 15316 40348
rect 15708 40402 15764 40908
rect 15708 40350 15710 40402
rect 15762 40350 15764 40402
rect 15708 40338 15764 40350
rect 16044 41972 16100 41982
rect 16156 41972 16212 42924
rect 16380 42868 16436 42878
rect 16380 42774 16436 42812
rect 16492 42756 16548 42766
rect 16492 42662 16548 42700
rect 16828 42642 16884 42654
rect 16828 42590 16830 42642
rect 16882 42590 16884 42642
rect 16828 42084 16884 42590
rect 16828 42018 16884 42028
rect 16044 41970 16212 41972
rect 16044 41918 16046 41970
rect 16098 41918 16212 41970
rect 16044 41916 16212 41918
rect 16716 41972 16772 41982
rect 15372 40292 15428 40302
rect 15372 40198 15428 40236
rect 15932 39620 15988 39630
rect 15932 39526 15988 39564
rect 16044 39396 16100 41916
rect 16716 41878 16772 41916
rect 16380 41860 16436 41870
rect 16380 41074 16436 41804
rect 16380 41022 16382 41074
rect 16434 41022 16436 41074
rect 16380 41010 16436 41022
rect 16492 41748 16548 41758
rect 16492 39956 16548 41692
rect 16716 40514 16772 40526
rect 16716 40462 16718 40514
rect 16770 40462 16772 40514
rect 16604 40180 16660 40190
rect 16604 40086 16660 40124
rect 16492 39900 16660 39956
rect 15932 39340 16100 39396
rect 16492 39506 16548 39518
rect 16492 39454 16494 39506
rect 16546 39454 16548 39506
rect 15260 38882 15316 38892
rect 15820 39060 15876 39070
rect 15708 38834 15764 38846
rect 15708 38782 15710 38834
rect 15762 38782 15764 38834
rect 15372 38612 15428 38622
rect 15372 38518 15428 38556
rect 15372 38388 15428 38398
rect 15372 37266 15428 38332
rect 15708 38052 15764 38782
rect 15820 38722 15876 39004
rect 15820 38670 15822 38722
rect 15874 38670 15876 38722
rect 15820 38658 15876 38670
rect 15708 37986 15764 37996
rect 15932 37604 15988 39340
rect 15932 37538 15988 37548
rect 16044 38834 16100 38846
rect 16044 38782 16046 38834
rect 16098 38782 16100 38834
rect 16044 37828 16100 38782
rect 16492 38388 16548 39454
rect 16492 38322 16548 38332
rect 16492 38164 16548 38174
rect 16156 37828 16212 37838
rect 16044 37826 16212 37828
rect 16044 37774 16158 37826
rect 16210 37774 16212 37826
rect 16044 37772 16212 37774
rect 15372 37214 15374 37266
rect 15426 37214 15428 37266
rect 15372 37202 15428 37214
rect 15932 37268 15988 37278
rect 16044 37268 16100 37772
rect 16156 37762 16212 37772
rect 15932 37266 16100 37268
rect 15932 37214 15934 37266
rect 15986 37214 16100 37266
rect 15932 37212 16100 37214
rect 16492 37266 16548 38108
rect 16492 37214 16494 37266
rect 16546 37214 16548 37266
rect 15148 36950 15204 36988
rect 15820 36594 15876 36606
rect 15820 36542 15822 36594
rect 15874 36542 15876 36594
rect 15036 35758 15038 35810
rect 15090 35758 15092 35810
rect 15036 35746 15092 35758
rect 15708 36482 15764 36494
rect 15708 36430 15710 36482
rect 15762 36430 15764 36482
rect 15708 35700 15764 36430
rect 15708 35634 15764 35644
rect 15820 35698 15876 36542
rect 15820 35646 15822 35698
rect 15874 35646 15876 35698
rect 14364 35522 14420 35532
rect 14140 33406 14142 33458
rect 14194 33406 14196 33458
rect 14140 33394 14196 33406
rect 14252 35140 14308 35150
rect 13804 33294 13806 33346
rect 13858 33294 13860 33346
rect 13804 33282 13860 33294
rect 14252 33234 14308 35084
rect 15372 34916 15428 34926
rect 15372 34914 15540 34916
rect 15372 34862 15374 34914
rect 15426 34862 15540 34914
rect 15372 34860 15540 34862
rect 15372 34850 15428 34860
rect 15148 34692 15204 34702
rect 15148 34354 15204 34636
rect 15148 34302 15150 34354
rect 15202 34302 15204 34354
rect 15148 34290 15204 34302
rect 15484 34020 15540 34860
rect 15820 34692 15876 35646
rect 15820 34626 15876 34636
rect 15484 33954 15540 33964
rect 15148 33572 15204 33582
rect 14588 33460 14644 33470
rect 14588 33366 14644 33404
rect 14812 33348 14868 33358
rect 14812 33254 14868 33292
rect 14252 33182 14254 33234
rect 14306 33182 14308 33234
rect 14252 33124 14308 33182
rect 13692 33068 13860 33124
rect 14252 33068 14532 33124
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31714 13524 31726
rect 13580 32562 13636 32574
rect 13580 32510 13582 32562
rect 13634 32510 13636 32562
rect 13580 31780 13636 32510
rect 13580 31714 13636 31724
rect 13692 32340 13748 32350
rect 13692 31778 13748 32284
rect 13692 31726 13694 31778
rect 13746 31726 13748 31778
rect 13692 31714 13748 31726
rect 13804 31778 13860 33068
rect 13804 31726 13806 31778
rect 13858 31726 13860 31778
rect 13804 31714 13860 31726
rect 13916 32676 13972 32686
rect 13356 31500 13524 31556
rect 13468 29764 13524 31500
rect 13916 31444 13972 32620
rect 13804 31388 13972 31444
rect 14028 32452 14084 32462
rect 13132 29362 13188 29372
rect 13244 29708 13524 29764
rect 13580 31332 13636 31342
rect 13580 30210 13636 31276
rect 13580 30158 13582 30210
rect 13634 30158 13636 30210
rect 12908 28590 12910 28642
rect 12962 28590 12964 28642
rect 12908 28578 12964 28590
rect 12796 28366 12798 28418
rect 12850 28366 12852 28418
rect 12796 28354 12852 28366
rect 13244 28082 13300 29708
rect 13468 29540 13524 29550
rect 13468 29426 13524 29484
rect 13468 29374 13470 29426
rect 13522 29374 13524 29426
rect 13468 29362 13524 29374
rect 13468 29204 13524 29214
rect 13468 29110 13524 29148
rect 13580 29092 13636 30158
rect 13580 29026 13636 29036
rect 13804 30210 13860 31388
rect 14028 31218 14084 32396
rect 14476 31948 14532 33068
rect 15148 32786 15204 33516
rect 15148 32734 15150 32786
rect 15202 32734 15204 32786
rect 15148 32722 15204 32734
rect 15820 33460 15876 33470
rect 15820 33346 15876 33404
rect 15820 33294 15822 33346
rect 15874 33294 15876 33346
rect 14588 32676 14644 32686
rect 14924 32676 14980 32686
rect 14644 32674 14980 32676
rect 14644 32622 14926 32674
rect 14978 32622 14980 32674
rect 14644 32620 14980 32622
rect 14588 32582 14644 32620
rect 14924 32610 14980 32620
rect 15372 32562 15428 32574
rect 15372 32510 15374 32562
rect 15426 32510 15428 32562
rect 14812 32340 14868 32350
rect 14812 32246 14868 32284
rect 15372 32116 15428 32510
rect 15372 32050 15428 32060
rect 14252 31892 14308 31902
rect 14476 31892 14644 31948
rect 14252 31798 14308 31836
rect 14028 31166 14030 31218
rect 14082 31166 14084 31218
rect 14028 31154 14084 31166
rect 14140 31780 14196 31790
rect 13916 30996 13972 31006
rect 13916 30902 13972 30940
rect 13804 30158 13806 30210
rect 13858 30158 13860 30210
rect 13468 28756 13524 28766
rect 13804 28756 13860 30158
rect 14140 30210 14196 31724
rect 14476 31332 14532 31342
rect 14476 31106 14532 31276
rect 14476 31054 14478 31106
rect 14530 31054 14532 31106
rect 14476 31042 14532 31054
rect 14140 30158 14142 30210
rect 14194 30158 14196 30210
rect 13244 28030 13246 28082
rect 13298 28030 13300 28082
rect 13244 28018 13300 28030
rect 13356 28754 13524 28756
rect 13356 28702 13470 28754
rect 13522 28702 13524 28754
rect 13356 28700 13524 28702
rect 13132 27858 13188 27870
rect 13132 27806 13134 27858
rect 13186 27806 13188 27858
rect 12348 27746 12404 27758
rect 12348 27694 12350 27746
rect 12402 27694 12404 27746
rect 12348 27300 12404 27694
rect 12348 27234 12404 27244
rect 13132 27300 13188 27806
rect 13356 27748 13412 28700
rect 13468 28690 13524 28700
rect 13580 28700 13860 28756
rect 14028 28868 14084 28878
rect 13356 27682 13412 27692
rect 13468 27858 13524 27870
rect 13468 27806 13470 27858
rect 13522 27806 13524 27858
rect 13132 27234 13188 27244
rect 12236 27134 12238 27186
rect 12290 27134 12292 27186
rect 12236 27122 12292 27134
rect 12348 27076 12404 27086
rect 12236 26964 12292 26974
rect 12124 25508 12180 25518
rect 12236 25508 12292 26908
rect 12348 26402 12404 27020
rect 13468 26962 13524 27806
rect 13580 27076 13636 28700
rect 14028 28644 14084 28812
rect 14028 28578 14084 28588
rect 13580 27010 13636 27020
rect 13692 28532 13748 28542
rect 13468 26910 13470 26962
rect 13522 26910 13524 26962
rect 12348 26350 12350 26402
rect 12402 26350 12404 26402
rect 12348 26338 12404 26350
rect 13244 26852 13300 26862
rect 13244 26290 13300 26796
rect 13468 26404 13524 26910
rect 13692 26964 13748 28476
rect 13916 28530 13972 28542
rect 13916 28478 13918 28530
rect 13970 28478 13972 28530
rect 13916 28308 13972 28478
rect 14028 28420 14084 28430
rect 14028 28326 14084 28364
rect 13916 28242 13972 28252
rect 14140 28084 14196 30158
rect 14252 30212 14308 30222
rect 14252 29426 14308 30156
rect 14252 29374 14254 29426
rect 14306 29374 14308 29426
rect 14252 29362 14308 29374
rect 14588 28644 14644 31892
rect 15484 31780 15540 31790
rect 15820 31780 15876 33294
rect 15932 32676 15988 37212
rect 16492 37156 16548 37214
rect 16604 38162 16660 39900
rect 16716 39060 16772 40462
rect 16940 40292 16996 55020
rect 18060 55076 18116 55412
rect 18396 55076 18452 55086
rect 18060 55074 18452 55076
rect 18060 55022 18398 55074
rect 18450 55022 18452 55074
rect 18060 55020 18452 55022
rect 17836 53844 17892 53854
rect 17836 53730 17892 53788
rect 17836 53678 17838 53730
rect 17890 53678 17892 53730
rect 17836 53666 17892 53678
rect 17948 53618 18004 53630
rect 17948 53566 17950 53618
rect 18002 53566 18004 53618
rect 17948 53508 18004 53566
rect 17948 53442 18004 53452
rect 17500 52948 17556 52958
rect 17500 52854 17556 52892
rect 17500 50932 17556 50942
rect 17388 48916 17444 48926
rect 17388 48822 17444 48860
rect 17052 45892 17108 45902
rect 17052 45798 17108 45836
rect 17500 45780 17556 50876
rect 17612 47460 17668 47470
rect 17668 47404 17780 47460
rect 17612 47366 17668 47404
rect 17724 46676 17780 47404
rect 17948 47124 18004 47134
rect 17724 46674 17892 46676
rect 17724 46622 17726 46674
rect 17778 46622 17892 46674
rect 17724 46620 17892 46622
rect 17724 46610 17780 46620
rect 17836 45890 17892 46620
rect 17836 45838 17838 45890
rect 17890 45838 17892 45890
rect 17836 45826 17892 45838
rect 17948 46562 18004 47068
rect 17948 46510 17950 46562
rect 18002 46510 18004 46562
rect 17948 46002 18004 46510
rect 17948 45950 17950 46002
rect 18002 45950 18004 46002
rect 17500 45724 17780 45780
rect 17500 45218 17556 45230
rect 17500 45166 17502 45218
rect 17554 45166 17556 45218
rect 17052 44212 17108 44222
rect 17052 44210 17220 44212
rect 17052 44158 17054 44210
rect 17106 44158 17220 44210
rect 17052 44156 17220 44158
rect 17052 44146 17108 44156
rect 17164 43428 17220 44156
rect 17500 43652 17556 45166
rect 17612 44996 17668 45006
rect 17724 44996 17780 45724
rect 17612 44994 17780 44996
rect 17612 44942 17614 44994
rect 17666 44942 17780 44994
rect 17612 44940 17780 44942
rect 17612 44930 17668 44940
rect 17836 43876 17892 43886
rect 17948 43876 18004 45950
rect 18060 45332 18116 55020
rect 18396 55010 18452 55020
rect 18284 54516 18340 54526
rect 18284 54422 18340 54460
rect 19068 54516 19124 54526
rect 18732 53844 18788 53854
rect 18732 53750 18788 53788
rect 18396 53730 18452 53742
rect 18396 53678 18398 53730
rect 18450 53678 18452 53730
rect 18172 53506 18228 53518
rect 18172 53454 18174 53506
rect 18226 53454 18228 53506
rect 18172 53058 18228 53454
rect 18396 53508 18452 53678
rect 19068 53618 19124 54460
rect 19628 54516 19684 56700
rect 19852 56690 19908 56700
rect 19964 56644 20020 57036
rect 20076 56980 20132 57598
rect 20300 57652 20356 57662
rect 20300 57558 20356 57596
rect 20188 56980 20244 56990
rect 20076 56978 20244 56980
rect 20076 56926 20190 56978
rect 20242 56926 20244 56978
rect 20076 56924 20244 56926
rect 20188 56914 20244 56924
rect 20300 56868 20356 56878
rect 20412 56868 20468 57820
rect 20524 57874 20580 60620
rect 21756 59668 21812 60620
rect 21980 59778 22036 59790
rect 21980 59726 21982 59778
rect 22034 59726 22036 59778
rect 21980 59668 22036 59726
rect 21756 59612 22036 59668
rect 21084 58996 21140 59006
rect 20524 57822 20526 57874
rect 20578 57822 20580 57874
rect 20524 57810 20580 57822
rect 20748 58324 20804 58334
rect 20748 57652 20804 58268
rect 20748 57558 20804 57596
rect 20748 56868 20804 56878
rect 20300 56866 20692 56868
rect 20300 56814 20302 56866
rect 20354 56814 20692 56866
rect 20300 56812 20692 56814
rect 20300 56802 20356 56812
rect 20076 56644 20132 56682
rect 19964 56642 20244 56644
rect 19964 56590 20078 56642
rect 20130 56590 20244 56642
rect 19964 56588 20244 56590
rect 20076 56578 20132 56588
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20188 56196 20244 56588
rect 20300 56196 20356 56206
rect 20188 56194 20356 56196
rect 20188 56142 20302 56194
rect 20354 56142 20356 56194
rect 20188 56140 20356 56142
rect 20300 56130 20356 56140
rect 20636 55972 20692 56812
rect 20748 56774 20804 56812
rect 20748 55972 20804 55982
rect 20636 55970 20804 55972
rect 20636 55918 20750 55970
rect 20802 55918 20804 55970
rect 20636 55916 20804 55918
rect 20748 55906 20804 55916
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19628 54450 19684 54460
rect 20524 53844 20580 53854
rect 19852 53732 19908 53742
rect 19852 53638 19908 53676
rect 19964 53732 20020 53742
rect 19964 53730 20468 53732
rect 19964 53678 19966 53730
rect 20018 53678 20468 53730
rect 19964 53676 20468 53678
rect 19964 53666 20020 53676
rect 19068 53566 19070 53618
rect 19122 53566 19124 53618
rect 19068 53554 19124 53566
rect 19404 53620 19460 53630
rect 18620 53508 18676 53518
rect 18396 53506 18676 53508
rect 18396 53454 18622 53506
rect 18674 53454 18676 53506
rect 18396 53452 18676 53454
rect 18172 53006 18174 53058
rect 18226 53006 18228 53058
rect 18172 52994 18228 53006
rect 18508 52274 18564 53452
rect 18620 53442 18676 53452
rect 18844 53508 18900 53518
rect 18844 53414 18900 53452
rect 18508 52222 18510 52274
rect 18562 52222 18564 52274
rect 18508 52210 18564 52222
rect 19404 52274 19460 53564
rect 19628 53508 19684 53518
rect 19628 52612 19684 53452
rect 20076 53508 20132 53546
rect 20300 53508 20356 53518
rect 20076 53442 20132 53452
rect 20188 53506 20356 53508
rect 20188 53454 20302 53506
rect 20354 53454 20356 53506
rect 20188 53452 20356 53454
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19628 52546 19684 52556
rect 19404 52222 19406 52274
rect 19458 52222 19460 52274
rect 19404 52210 19460 52222
rect 20188 52274 20244 53452
rect 20300 53442 20356 53452
rect 20188 52222 20190 52274
rect 20242 52222 20244 52274
rect 20188 52210 20244 52222
rect 20300 52836 20356 52846
rect 19180 52164 19236 52174
rect 19180 52070 19236 52108
rect 20300 52164 20356 52780
rect 20412 52386 20468 53676
rect 20524 53506 20580 53788
rect 20636 53620 20692 53630
rect 20636 53526 20692 53564
rect 20524 53454 20526 53506
rect 20578 53454 20580 53506
rect 20524 52836 20580 53454
rect 20636 53284 20692 53294
rect 20636 52948 20692 53228
rect 20636 52854 20692 52892
rect 20524 52770 20580 52780
rect 20412 52334 20414 52386
rect 20466 52334 20468 52386
rect 20412 52322 20468 52334
rect 20524 52612 20580 52622
rect 20300 52098 20356 52108
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19628 50482 19684 50494
rect 19628 50430 19630 50482
rect 19682 50430 19684 50482
rect 19628 50428 19684 50430
rect 20524 50428 20580 52556
rect 20748 52388 20804 52398
rect 20748 52294 20804 52332
rect 19516 50372 19684 50428
rect 19740 50372 19796 50382
rect 20412 50372 20580 50428
rect 19292 49924 19348 49934
rect 19292 49830 19348 49868
rect 19180 49810 19236 49822
rect 19180 49758 19182 49810
rect 19234 49758 19236 49810
rect 19180 49700 19236 49758
rect 19180 49634 19236 49644
rect 19404 49812 19460 49822
rect 19292 49588 19348 49598
rect 19404 49588 19460 49756
rect 19292 49586 19460 49588
rect 19292 49534 19294 49586
rect 19346 49534 19460 49586
rect 19292 49532 19460 49534
rect 19292 49522 19348 49532
rect 19068 49140 19124 49150
rect 19068 48468 19124 49084
rect 19516 49138 19572 50372
rect 19740 50370 20244 50372
rect 19740 50318 19742 50370
rect 19794 50318 20244 50370
rect 19740 50316 20244 50318
rect 19740 50306 19796 50316
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20188 49924 20244 50316
rect 20300 49924 20356 49934
rect 20188 49868 20300 49924
rect 20300 49810 20356 49868
rect 20412 49922 20468 50372
rect 20412 49870 20414 49922
rect 20466 49870 20468 49922
rect 20412 49858 20468 49870
rect 20300 49758 20302 49810
rect 20354 49758 20356 49810
rect 19740 49700 19796 49710
rect 19516 49086 19518 49138
rect 19570 49086 19572 49138
rect 19516 49074 19572 49086
rect 19628 49644 19740 49700
rect 19068 48466 19348 48468
rect 19068 48414 19070 48466
rect 19122 48414 19348 48466
rect 19068 48412 19348 48414
rect 19068 48402 19124 48412
rect 19068 47570 19124 47582
rect 19068 47518 19070 47570
rect 19122 47518 19124 47570
rect 18172 47460 18228 47470
rect 18172 47366 18228 47404
rect 19068 47460 19124 47518
rect 19068 47394 19124 47404
rect 18284 47346 18340 47358
rect 18284 47294 18286 47346
rect 18338 47294 18340 47346
rect 18284 47236 18340 47294
rect 18284 47170 18340 47180
rect 18620 47234 18676 47246
rect 18620 47182 18622 47234
rect 18674 47182 18676 47234
rect 18620 47124 18676 47182
rect 18620 47058 18676 47068
rect 18172 46116 18228 46126
rect 18172 46022 18228 46060
rect 19292 46004 19348 48412
rect 19628 48130 19684 49644
rect 19740 49634 19796 49644
rect 20076 48914 20132 48926
rect 20076 48862 20078 48914
rect 20130 48862 20132 48914
rect 20076 48804 20132 48862
rect 20188 48916 20244 48926
rect 20188 48822 20244 48860
rect 20076 48738 20132 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20300 48468 20356 49758
rect 20524 49700 20580 49710
rect 20524 49606 20580 49644
rect 20412 48914 20468 48926
rect 20412 48862 20414 48914
rect 20466 48862 20468 48914
rect 20412 48692 20468 48862
rect 20636 48916 20692 48926
rect 20636 48822 20692 48860
rect 20412 48626 20468 48636
rect 20524 48804 20580 48814
rect 19964 48412 20356 48468
rect 19964 48242 20020 48412
rect 20412 48356 20468 48366
rect 20524 48356 20580 48748
rect 20412 48354 20580 48356
rect 20412 48302 20414 48354
rect 20466 48302 20580 48354
rect 20412 48300 20580 48302
rect 20412 48290 20468 48300
rect 19964 48190 19966 48242
rect 20018 48190 20020 48242
rect 19964 48178 20020 48190
rect 19628 48078 19630 48130
rect 19682 48078 19684 48130
rect 19628 48066 19684 48078
rect 20972 48132 21028 48142
rect 20972 48038 21028 48076
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19404 46676 19460 46686
rect 19404 46582 19460 46620
rect 19740 46452 19796 46462
rect 19740 46358 19796 46396
rect 18060 45276 18228 45332
rect 17892 43820 18004 43876
rect 18060 45106 18116 45118
rect 18060 45054 18062 45106
rect 18114 45054 18116 45106
rect 17836 43810 17892 43820
rect 18060 43764 18116 45054
rect 18060 43698 18116 43708
rect 17164 41074 17220 43372
rect 17276 43596 17556 43652
rect 17276 41748 17332 43596
rect 17500 43538 17556 43596
rect 17500 43486 17502 43538
rect 17554 43486 17556 43538
rect 17500 43474 17556 43486
rect 17724 43650 17780 43662
rect 17724 43598 17726 43650
rect 17778 43598 17780 43650
rect 17276 41682 17332 41692
rect 17388 43426 17444 43438
rect 17388 43374 17390 43426
rect 17442 43374 17444 43426
rect 17164 41022 17166 41074
rect 17218 41022 17220 41074
rect 17164 41010 17220 41022
rect 17388 40516 17444 43374
rect 17724 42196 17780 43598
rect 18172 43540 18228 45276
rect 18620 45106 18676 45118
rect 18620 45054 18622 45106
rect 18674 45054 18676 45106
rect 17388 40450 17444 40460
rect 17500 42140 17780 42196
rect 18060 43484 18228 43540
rect 18396 43650 18452 43662
rect 18396 43598 18398 43650
rect 18450 43598 18452 43650
rect 16940 40226 16996 40236
rect 17276 40404 17332 40414
rect 16716 38994 16772 39004
rect 16604 38110 16606 38162
rect 16658 38110 16660 38162
rect 16604 37268 16660 38110
rect 17052 38050 17108 38062
rect 17052 37998 17054 38050
rect 17106 37998 17108 38050
rect 17052 37940 17108 37998
rect 16828 37716 16884 37726
rect 16604 37202 16660 37212
rect 16716 37492 16772 37502
rect 16268 37100 16548 37156
rect 16716 37154 16772 37436
rect 16828 37378 16884 37660
rect 16828 37326 16830 37378
rect 16882 37326 16884 37378
rect 16828 37314 16884 37326
rect 16716 37102 16718 37154
rect 16770 37102 16772 37154
rect 16268 36594 16324 37100
rect 16716 37090 16772 37102
rect 17052 37044 17108 37884
rect 16828 36988 17108 37044
rect 16828 36932 16884 36988
rect 16268 36542 16270 36594
rect 16322 36542 16324 36594
rect 16268 36530 16324 36542
rect 16716 36876 16884 36932
rect 16044 35588 16100 35598
rect 16044 32900 16100 35532
rect 16268 34802 16324 34814
rect 16268 34750 16270 34802
rect 16322 34750 16324 34802
rect 16268 34692 16324 34750
rect 16268 34626 16324 34636
rect 16716 34690 16772 36876
rect 17276 36594 17332 40348
rect 17500 40402 17556 42140
rect 18060 41524 18116 43484
rect 18396 42980 18452 43598
rect 18620 43652 18676 45054
rect 18732 44996 18788 45006
rect 18732 44322 18788 44940
rect 19292 44436 19348 45948
rect 20188 46228 20244 46238
rect 20188 46002 20244 46172
rect 21084 46228 21140 58940
rect 21308 56868 21364 56878
rect 21756 56868 21812 59612
rect 22092 59556 22148 62860
rect 22428 61460 22484 61470
rect 22428 61458 22596 61460
rect 22428 61406 22430 61458
rect 22482 61406 22596 61458
rect 22428 61404 22596 61406
rect 22428 61394 22484 61404
rect 22540 60228 22596 61404
rect 22652 61348 22708 61358
rect 22652 60788 22708 61292
rect 22652 60694 22708 60732
rect 23212 60676 23268 60686
rect 23212 60582 23268 60620
rect 23548 60676 23604 63868
rect 23660 63858 23716 63868
rect 24780 63252 24836 64542
rect 25452 64484 25508 65326
rect 27356 65378 27412 67172
rect 29148 66162 29204 67172
rect 29148 66110 29150 66162
rect 29202 66110 29204 66162
rect 29148 66098 29204 66110
rect 31164 66162 31220 67172
rect 31164 66110 31166 66162
rect 31218 66110 31220 66162
rect 31164 66098 31220 66110
rect 33180 66162 33236 67172
rect 33180 66110 33182 66162
rect 33234 66110 33236 66162
rect 33180 66098 33236 66110
rect 35084 66164 35140 67172
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 36988 66386 37044 69200
rect 39004 66500 39060 69200
rect 39004 66434 39060 66444
rect 40796 66500 40852 66510
rect 40796 66406 40852 66444
rect 36988 66334 36990 66386
rect 37042 66334 37044 66386
rect 36988 66322 37044 66334
rect 39228 66276 39284 66286
rect 39788 66276 39844 66286
rect 39228 66274 39396 66276
rect 39228 66222 39230 66274
rect 39282 66222 39396 66274
rect 39228 66220 39396 66222
rect 39228 66210 39284 66220
rect 35196 66164 35252 66174
rect 35084 66162 35252 66164
rect 35084 66110 35198 66162
rect 35250 66110 35252 66162
rect 35084 66108 35252 66110
rect 35196 66098 35252 66108
rect 34860 65602 34916 65614
rect 34860 65550 34862 65602
rect 34914 65550 34916 65602
rect 27356 65326 27358 65378
rect 27410 65326 27412 65378
rect 27356 65314 27412 65326
rect 29708 65490 29764 65502
rect 29708 65438 29710 65490
rect 29762 65438 29764 65490
rect 29708 65380 29764 65438
rect 33852 65492 33908 65502
rect 30268 65380 30324 65390
rect 29708 65378 30324 65380
rect 29708 65326 30270 65378
rect 30322 65326 30324 65378
rect 29708 65324 30324 65326
rect 30268 64932 30324 65324
rect 30268 64866 30324 64876
rect 25452 64418 25508 64428
rect 26908 64818 26964 64830
rect 33516 64820 33572 64830
rect 26908 64766 26910 64818
rect 26962 64766 26964 64818
rect 26684 64260 26740 64270
rect 26908 64260 26964 64766
rect 32508 64818 33572 64820
rect 32508 64766 33518 64818
rect 33570 64766 33572 64818
rect 32508 64764 33572 64766
rect 27804 64708 27860 64718
rect 26740 64204 26964 64260
rect 27244 64482 27300 64494
rect 27244 64430 27246 64482
rect 27298 64430 27300 64482
rect 26684 63922 26740 64204
rect 26684 63870 26686 63922
rect 26738 63870 26740 63922
rect 26684 63858 26740 63870
rect 26348 63810 26404 63822
rect 27132 63812 27188 63822
rect 26348 63758 26350 63810
rect 26402 63758 26404 63810
rect 26348 63700 26404 63758
rect 24780 63186 24836 63196
rect 26236 63252 26292 63262
rect 26236 63158 26292 63196
rect 26124 63026 26180 63038
rect 26124 62974 26126 63026
rect 26178 62974 26180 63026
rect 26124 62916 26180 62974
rect 26124 62850 26180 62860
rect 25900 62132 25956 62142
rect 24556 61682 24612 61694
rect 24556 61630 24558 61682
rect 24610 61630 24612 61682
rect 24556 61460 24612 61630
rect 24892 61460 24948 61470
rect 24556 61458 24948 61460
rect 24556 61406 24894 61458
rect 24946 61406 24948 61458
rect 24556 61404 24948 61406
rect 23548 60610 23604 60620
rect 22652 60228 22708 60238
rect 22540 60226 22708 60228
rect 22540 60174 22654 60226
rect 22706 60174 22708 60226
rect 22540 60172 22708 60174
rect 22652 60162 22708 60172
rect 23996 60002 24052 60014
rect 23996 59950 23998 60002
rect 24050 59950 24052 60002
rect 22988 59892 23044 59902
rect 23324 59892 23380 59902
rect 22988 59890 23380 59892
rect 22988 59838 22990 59890
rect 23042 59838 23326 59890
rect 23378 59838 23380 59890
rect 22988 59836 23380 59838
rect 22988 59826 23044 59836
rect 23324 59826 23380 59836
rect 23996 59892 24052 59950
rect 22764 59780 22820 59790
rect 22764 59778 22932 59780
rect 22764 59726 22766 59778
rect 22818 59726 22932 59778
rect 22764 59724 22932 59726
rect 22764 59714 22820 59724
rect 21308 56866 21812 56868
rect 21308 56814 21310 56866
rect 21362 56814 21812 56866
rect 21308 56812 21812 56814
rect 21980 59500 22148 59556
rect 21308 55524 21364 56812
rect 21196 53844 21252 53854
rect 21196 53060 21252 53788
rect 21308 53284 21364 55468
rect 21364 53228 21588 53284
rect 21308 53218 21364 53228
rect 21420 53060 21476 53070
rect 21196 53058 21476 53060
rect 21196 53006 21422 53058
rect 21474 53006 21476 53058
rect 21196 53004 21476 53006
rect 21420 52994 21476 53004
rect 21532 52274 21588 53228
rect 21532 52222 21534 52274
rect 21586 52222 21588 52274
rect 21532 52210 21588 52222
rect 21980 50036 22036 59500
rect 22876 57762 22932 59724
rect 22876 57710 22878 57762
rect 22930 57710 22932 57762
rect 22764 57652 22820 57662
rect 22092 57650 22820 57652
rect 22092 57598 22766 57650
rect 22818 57598 22820 57650
rect 22092 57596 22820 57598
rect 22092 56978 22148 57596
rect 22764 57586 22820 57596
rect 22092 56926 22094 56978
rect 22146 56926 22148 56978
rect 22092 56914 22148 56926
rect 22652 57426 22708 57438
rect 22652 57374 22654 57426
rect 22706 57374 22708 57426
rect 22652 56306 22708 57374
rect 22652 56254 22654 56306
rect 22706 56254 22708 56306
rect 22652 56242 22708 56254
rect 22876 55468 22932 57710
rect 23996 57762 24052 59836
rect 24892 59890 24948 61404
rect 25004 61348 25060 61358
rect 25564 61348 25620 61358
rect 25900 61348 25956 62076
rect 26348 61460 26404 63644
rect 27020 63810 27188 63812
rect 27020 63758 27134 63810
rect 27186 63758 27188 63810
rect 27020 63756 27188 63758
rect 26684 63140 26740 63150
rect 26684 63046 26740 63084
rect 26460 63028 26516 63038
rect 26460 62934 26516 62972
rect 27020 62916 27076 63756
rect 27132 63746 27188 63756
rect 27244 63700 27300 64430
rect 27356 64482 27412 64494
rect 27356 64430 27358 64482
rect 27410 64430 27412 64482
rect 27356 64036 27412 64430
rect 27468 64482 27524 64494
rect 27468 64430 27470 64482
rect 27522 64430 27524 64482
rect 27468 64260 27524 64430
rect 27468 64194 27524 64204
rect 27804 64146 27860 64652
rect 27916 64706 27972 64718
rect 27916 64654 27918 64706
rect 27970 64654 27972 64706
rect 27916 64484 27972 64654
rect 29036 64706 29092 64718
rect 29036 64654 29038 64706
rect 29090 64654 29092 64706
rect 28700 64484 28756 64494
rect 29036 64484 29092 64654
rect 27916 64428 28420 64484
rect 27804 64094 27806 64146
rect 27858 64094 27860 64146
rect 27804 64082 27860 64094
rect 28140 64260 28196 64270
rect 27468 64036 27524 64046
rect 27356 64034 27524 64036
rect 27356 63982 27470 64034
rect 27522 63982 27524 64034
rect 27356 63980 27524 63982
rect 27468 63970 27524 63980
rect 27580 64034 27636 64046
rect 27580 63982 27582 64034
rect 27634 63982 27636 64034
rect 27580 63812 27636 63982
rect 28028 63924 28084 63934
rect 27916 63922 28084 63924
rect 27916 63870 28030 63922
rect 28082 63870 28084 63922
rect 27916 63868 28084 63870
rect 27580 63756 27860 63812
rect 27244 63634 27300 63644
rect 27132 63140 27188 63150
rect 27132 63046 27188 63084
rect 27580 63138 27636 63150
rect 27580 63086 27582 63138
rect 27634 63086 27636 63138
rect 27020 62822 27076 62860
rect 27244 63028 27300 63038
rect 27244 62914 27300 62972
rect 27244 62862 27246 62914
rect 27298 62862 27300 62914
rect 27244 62356 27300 62862
rect 27580 62916 27636 63086
rect 27804 63138 27860 63756
rect 27804 63086 27806 63138
rect 27858 63086 27860 63138
rect 27804 63074 27860 63086
rect 27580 62850 27636 62860
rect 27244 62290 27300 62300
rect 27692 62244 27748 62254
rect 27916 62244 27972 63868
rect 28028 63858 28084 63868
rect 28140 63700 28196 64204
rect 28028 63644 28196 63700
rect 28252 63700 28308 63710
rect 28028 63026 28084 63644
rect 28140 63140 28196 63150
rect 28252 63140 28308 63644
rect 28140 63138 28308 63140
rect 28140 63086 28142 63138
rect 28194 63086 28308 63138
rect 28140 63084 28308 63086
rect 28140 63074 28196 63084
rect 28028 62974 28030 63026
rect 28082 62974 28084 63026
rect 28028 62962 28084 62974
rect 28364 62356 28420 64428
rect 28588 64482 29092 64484
rect 28588 64430 28702 64482
rect 28754 64430 29092 64482
rect 28588 64428 29092 64430
rect 29148 64708 29204 64718
rect 28364 62290 28420 62300
rect 28476 62916 28532 62926
rect 28588 62916 28644 64428
rect 28700 64418 28756 64428
rect 28812 63812 28868 63822
rect 28812 63810 29092 63812
rect 28812 63758 28814 63810
rect 28866 63758 29092 63810
rect 28812 63756 29092 63758
rect 28812 63746 28868 63756
rect 28532 62914 28644 62916
rect 28532 62862 28590 62914
rect 28642 62862 28644 62914
rect 28532 62860 28644 62862
rect 27692 62242 27972 62244
rect 27692 62190 27694 62242
rect 27746 62190 27972 62242
rect 27692 62188 27972 62190
rect 27692 62132 27748 62188
rect 27692 62066 27748 62076
rect 25004 61346 25508 61348
rect 25004 61294 25006 61346
rect 25058 61294 25508 61346
rect 25004 61292 25508 61294
rect 25004 61282 25060 61292
rect 24892 59838 24894 59890
rect 24946 59838 24948 59890
rect 24892 59826 24948 59838
rect 25116 61124 25172 61134
rect 24668 59556 24724 59566
rect 24668 57876 24724 59500
rect 25116 59108 25172 61068
rect 25452 61012 25508 61292
rect 25564 61254 25620 61292
rect 25788 61346 25956 61348
rect 25788 61294 25902 61346
rect 25954 61294 25956 61346
rect 25788 61292 25956 61294
rect 25452 60918 25508 60956
rect 25452 60788 25508 60798
rect 25228 60564 25284 60574
rect 25452 60564 25508 60732
rect 25676 60676 25732 60686
rect 25788 60676 25844 61292
rect 25900 61282 25956 61292
rect 26124 61404 26404 61460
rect 26012 61012 26068 61022
rect 26012 60918 26068 60956
rect 25900 60788 25956 60798
rect 25900 60694 25956 60732
rect 25732 60620 25844 60676
rect 25676 60610 25732 60620
rect 25228 60562 25508 60564
rect 25228 60510 25230 60562
rect 25282 60510 25508 60562
rect 25228 60508 25508 60510
rect 25228 60498 25284 60508
rect 25452 60114 25508 60508
rect 25564 60562 25620 60574
rect 25564 60510 25566 60562
rect 25618 60510 25620 60562
rect 25564 60228 25620 60510
rect 25564 60172 25956 60228
rect 25452 60062 25454 60114
rect 25506 60062 25508 60114
rect 25452 60050 25508 60062
rect 25900 60002 25956 60172
rect 25900 59950 25902 60002
rect 25954 59950 25956 60002
rect 25900 59938 25956 59950
rect 25116 59042 25172 59052
rect 26012 59778 26068 59790
rect 26012 59726 26014 59778
rect 26066 59726 26068 59778
rect 25788 58660 25844 58670
rect 24668 57810 24724 57820
rect 25340 58658 25844 58660
rect 25340 58606 25790 58658
rect 25842 58606 25844 58658
rect 25340 58604 25844 58606
rect 25340 58322 25396 58604
rect 25788 58594 25844 58604
rect 25676 58436 25732 58446
rect 25676 58342 25732 58380
rect 25340 58270 25342 58322
rect 25394 58270 25396 58322
rect 25340 57874 25396 58270
rect 26012 58324 26068 59726
rect 26124 58658 26180 61404
rect 28140 61236 28196 61246
rect 27244 60898 27300 60910
rect 27244 60846 27246 60898
rect 27298 60846 27300 60898
rect 26236 60786 26292 60798
rect 26236 60734 26238 60786
rect 26290 60734 26292 60786
rect 26236 60004 26292 60734
rect 27132 60788 27188 60798
rect 26460 60004 26516 60014
rect 26236 60002 26516 60004
rect 26236 59950 26462 60002
rect 26514 59950 26516 60002
rect 26236 59948 26516 59950
rect 26460 59938 26516 59948
rect 26572 59892 26628 59902
rect 26572 59798 26628 59836
rect 27020 59444 27076 59454
rect 27132 59444 27188 60732
rect 27244 60564 27300 60846
rect 27804 60900 27860 60910
rect 27804 60806 27860 60844
rect 27244 60498 27300 60508
rect 27468 60786 27524 60798
rect 27468 60734 27470 60786
rect 27522 60734 27524 60786
rect 27468 60004 27524 60734
rect 27692 60786 27748 60798
rect 27692 60734 27694 60786
rect 27746 60734 27748 60786
rect 27692 60676 27748 60734
rect 27916 60788 27972 60798
rect 27916 60694 27972 60732
rect 27692 60610 27748 60620
rect 28028 60564 28084 60574
rect 27916 60508 28028 60564
rect 27804 60116 27860 60126
rect 27916 60116 27972 60508
rect 28028 60498 28084 60508
rect 27804 60114 27972 60116
rect 27804 60062 27806 60114
rect 27858 60062 27972 60114
rect 27804 60060 27972 60062
rect 27804 60050 27860 60060
rect 27468 59938 27524 59948
rect 28028 60002 28084 60014
rect 28028 59950 28030 60002
rect 28082 59950 28084 60002
rect 27020 59442 27188 59444
rect 27020 59390 27022 59442
rect 27074 59390 27188 59442
rect 27020 59388 27188 59390
rect 27468 59778 27524 59790
rect 27468 59726 27470 59778
rect 27522 59726 27524 59778
rect 27020 59378 27076 59388
rect 27356 59220 27412 59230
rect 27468 59220 27524 59726
rect 27356 59218 27524 59220
rect 27356 59166 27358 59218
rect 27410 59166 27524 59218
rect 27356 59164 27524 59166
rect 27356 59154 27412 59164
rect 26124 58606 26126 58658
rect 26178 58606 26180 58658
rect 26124 58594 26180 58606
rect 27468 59108 27524 59164
rect 27804 59108 27860 59118
rect 28028 59108 28084 59950
rect 27468 59106 28084 59108
rect 27468 59054 27806 59106
rect 27858 59054 28084 59106
rect 27468 59052 28084 59054
rect 27356 58548 27412 58558
rect 27020 58546 27412 58548
rect 27020 58494 27358 58546
rect 27410 58494 27412 58546
rect 27020 58492 27412 58494
rect 26684 58436 26740 58446
rect 26684 58342 26740 58380
rect 26012 58258 26068 58268
rect 25340 57822 25342 57874
rect 25394 57822 25396 57874
rect 25340 57810 25396 57822
rect 25452 58210 25508 58222
rect 25452 58158 25454 58210
rect 25506 58158 25508 58210
rect 23996 57710 23998 57762
rect 24050 57710 24052 57762
rect 23996 57698 24052 57710
rect 23660 57650 23716 57662
rect 23660 57598 23662 57650
rect 23714 57598 23716 57650
rect 22988 56196 23044 56206
rect 22988 56082 23044 56140
rect 23660 56196 23716 57598
rect 24668 57650 24724 57662
rect 24668 57598 24670 57650
rect 24722 57598 24724 57650
rect 23660 56130 23716 56140
rect 23772 57538 23828 57550
rect 23772 57486 23774 57538
rect 23826 57486 23828 57538
rect 22988 56030 22990 56082
rect 23042 56030 23044 56082
rect 22988 56018 23044 56030
rect 22428 55412 22932 55468
rect 23660 55860 23716 55870
rect 23548 55412 23604 55422
rect 23660 55412 23716 55804
rect 22316 53844 22372 53854
rect 22316 53750 22372 53788
rect 22428 53506 22484 55412
rect 23548 55410 23716 55412
rect 23548 55358 23550 55410
rect 23602 55358 23716 55410
rect 23548 55356 23716 55358
rect 23772 55410 23828 57486
rect 24668 57090 24724 57598
rect 25452 57204 25508 58158
rect 26124 58210 26180 58222
rect 26124 58158 26126 58210
rect 26178 58158 26180 58210
rect 24668 57038 24670 57090
rect 24722 57038 24724 57090
rect 24668 57026 24724 57038
rect 25116 57148 25508 57204
rect 25676 57652 25732 57662
rect 26124 57652 26180 58158
rect 25676 57650 26180 57652
rect 25676 57598 25678 57650
rect 25730 57598 26180 57650
rect 25676 57596 26180 57598
rect 26236 58212 26292 58222
rect 24220 56978 24276 56990
rect 24220 56926 24222 56978
rect 24274 56926 24276 56978
rect 24220 56644 24276 56926
rect 24780 56756 24836 56766
rect 25116 56756 25172 57148
rect 25676 57092 25732 57596
rect 25676 57026 25732 57036
rect 25452 56868 25508 56878
rect 26124 56868 26180 56878
rect 25452 56866 26180 56868
rect 25452 56814 25454 56866
rect 25506 56814 26126 56866
rect 26178 56814 26180 56866
rect 25452 56812 26180 56814
rect 25452 56802 25508 56812
rect 24780 56754 25172 56756
rect 24780 56702 24782 56754
rect 24834 56702 25118 56754
rect 25170 56702 25172 56754
rect 24780 56700 25172 56702
rect 24668 56644 24724 56654
rect 24220 56642 24724 56644
rect 24220 56590 24670 56642
rect 24722 56590 24724 56642
rect 24220 56588 24724 56590
rect 23772 55358 23774 55410
rect 23826 55358 23828 55410
rect 23548 55346 23604 55356
rect 23772 55346 23828 55358
rect 23884 56196 23940 56206
rect 24220 56196 24276 56588
rect 24668 56578 24724 56588
rect 24780 56420 24836 56700
rect 25116 56690 25172 56700
rect 23884 56194 24276 56196
rect 23884 56142 23886 56194
rect 23938 56142 24276 56194
rect 23884 56140 24276 56142
rect 24444 56364 24836 56420
rect 23884 55298 23940 56140
rect 23884 55246 23886 55298
rect 23938 55246 23940 55298
rect 23884 55234 23940 55246
rect 24108 55972 24164 55982
rect 23324 54068 23380 54078
rect 23324 53954 23380 54012
rect 23324 53902 23326 53954
rect 23378 53902 23380 53954
rect 23324 53890 23380 53902
rect 24108 53842 24164 55916
rect 24444 55970 24500 56364
rect 24444 55918 24446 55970
rect 24498 55918 24500 55970
rect 24444 55860 24500 55918
rect 24444 55794 24500 55804
rect 25340 55970 25396 55982
rect 25340 55918 25342 55970
rect 25394 55918 25396 55970
rect 25228 55524 25284 55534
rect 25340 55468 25396 55918
rect 25228 55412 25396 55468
rect 24108 53790 24110 53842
rect 24162 53790 24164 53842
rect 24108 53778 24164 53790
rect 24780 54068 24836 54078
rect 23884 53732 23940 53742
rect 24780 53732 24836 54012
rect 23884 53730 24052 53732
rect 23884 53678 23886 53730
rect 23938 53678 24052 53730
rect 23884 53676 24052 53678
rect 23884 53666 23940 53676
rect 22652 53620 22708 53630
rect 22428 53454 22430 53506
rect 22482 53454 22484 53506
rect 22428 51492 22484 53454
rect 22540 53618 22708 53620
rect 22540 53566 22654 53618
rect 22706 53566 22708 53618
rect 22540 53564 22708 53566
rect 22540 51938 22596 53564
rect 22652 53554 22708 53564
rect 23100 53620 23156 53630
rect 23100 53526 23156 53564
rect 23548 53620 23604 53630
rect 23212 53508 23268 53518
rect 23212 53414 23268 53452
rect 23100 52948 23156 52958
rect 23100 52388 23156 52892
rect 23548 52834 23604 53564
rect 23884 53508 23940 53518
rect 23884 53058 23940 53452
rect 23996 53170 24052 53676
rect 24556 53730 24836 53732
rect 24556 53678 24782 53730
rect 24834 53678 24836 53730
rect 24556 53676 24836 53678
rect 23996 53118 23998 53170
rect 24050 53118 24052 53170
rect 23996 53106 24052 53118
rect 24332 53620 24388 53630
rect 23884 53006 23886 53058
rect 23938 53006 23940 53058
rect 23884 52994 23940 53006
rect 24220 52948 24276 52958
rect 24220 52854 24276 52892
rect 23548 52782 23550 52834
rect 23602 52782 23604 52834
rect 23548 52770 23604 52782
rect 23100 52162 23156 52332
rect 23100 52110 23102 52162
rect 23154 52110 23156 52162
rect 23100 52098 23156 52110
rect 24332 52050 24388 53564
rect 24556 52274 24612 53676
rect 24780 53666 24836 53676
rect 25228 53732 25284 55412
rect 25228 53730 25396 53732
rect 25228 53678 25230 53730
rect 25282 53678 25396 53730
rect 25228 53676 25396 53678
rect 25228 53666 25284 53676
rect 24668 53172 24724 53182
rect 24668 53078 24724 53116
rect 25340 53172 25396 53676
rect 25340 53078 25396 53116
rect 24556 52222 24558 52274
rect 24610 52222 24612 52274
rect 24556 52210 24612 52222
rect 24332 51998 24334 52050
rect 24386 51998 24388 52050
rect 24332 51986 24388 51998
rect 22540 51886 22542 51938
rect 22594 51886 22596 51938
rect 22540 51874 22596 51886
rect 22428 51426 22484 51436
rect 23772 51492 23828 51502
rect 21980 49970 22036 49980
rect 21532 49924 21588 49934
rect 21532 49922 21700 49924
rect 21532 49870 21534 49922
rect 21586 49870 21700 49922
rect 21532 49868 21700 49870
rect 21532 49858 21588 49868
rect 21196 49810 21252 49822
rect 21196 49758 21198 49810
rect 21250 49758 21252 49810
rect 21196 49588 21252 49758
rect 21420 49812 21476 49822
rect 21420 49718 21476 49756
rect 21532 49588 21588 49598
rect 21196 49586 21588 49588
rect 21196 49534 21534 49586
rect 21586 49534 21588 49586
rect 21196 49532 21588 49534
rect 21532 49522 21588 49532
rect 21420 48916 21476 48926
rect 21420 48822 21476 48860
rect 21308 48804 21364 48814
rect 21308 48710 21364 48748
rect 21532 48804 21588 48814
rect 21644 48804 21700 49868
rect 23772 49812 23828 51436
rect 25452 50594 25508 50606
rect 25452 50542 25454 50594
rect 25506 50542 25508 50594
rect 25116 50484 25172 50494
rect 25452 50484 25508 50542
rect 25116 50482 25508 50484
rect 25116 50430 25118 50482
rect 25170 50430 25508 50482
rect 25116 50428 25508 50430
rect 23772 49810 23940 49812
rect 23772 49758 23774 49810
rect 23826 49758 23940 49810
rect 23772 49756 23940 49758
rect 23772 49746 23828 49756
rect 23660 49698 23716 49710
rect 23660 49646 23662 49698
rect 23714 49646 23716 49698
rect 23436 49588 23492 49598
rect 22092 49586 23492 49588
rect 22092 49534 23438 49586
rect 23490 49534 23492 49586
rect 22092 49532 23492 49534
rect 21532 48802 21700 48804
rect 21532 48750 21534 48802
rect 21586 48750 21700 48802
rect 21532 48748 21700 48750
rect 21980 49026 22036 49038
rect 21980 48974 21982 49026
rect 22034 48974 22036 49026
rect 21532 48692 21588 48748
rect 21532 47684 21588 48636
rect 21980 48132 22036 48974
rect 22092 48466 22148 49532
rect 23436 49522 23492 49532
rect 22540 49140 22596 49150
rect 22540 49046 22596 49084
rect 22988 49140 23044 49150
rect 22988 49026 23044 49084
rect 23660 49138 23716 49646
rect 23660 49086 23662 49138
rect 23714 49086 23716 49138
rect 23660 49074 23716 49086
rect 22988 48974 22990 49026
rect 23042 48974 23044 49026
rect 22988 48962 23044 48974
rect 22092 48414 22094 48466
rect 22146 48414 22148 48466
rect 22092 48402 22148 48414
rect 23660 48804 23716 48814
rect 23660 48354 23716 48748
rect 23660 48302 23662 48354
rect 23714 48302 23716 48354
rect 23660 48290 23716 48302
rect 21980 48066 22036 48076
rect 22428 48242 22484 48254
rect 22428 48190 22430 48242
rect 22482 48190 22484 48242
rect 21532 47618 21588 47628
rect 22428 47460 22484 48190
rect 23436 48132 23492 48142
rect 22652 47684 22708 47694
rect 22652 47590 22708 47628
rect 23100 47572 23156 47582
rect 23100 47478 23156 47516
rect 22876 47460 22932 47470
rect 22428 47458 22932 47460
rect 22428 47406 22878 47458
rect 22930 47406 22932 47458
rect 22428 47404 22932 47406
rect 22876 46340 22932 47404
rect 22988 46340 23044 46350
rect 22876 46284 22988 46340
rect 22988 46274 23044 46284
rect 21084 46162 21140 46172
rect 20188 45950 20190 46002
rect 20242 45950 20244 46002
rect 20188 45938 20244 45950
rect 20748 45668 20804 45678
rect 20748 45574 20804 45612
rect 21420 45668 21476 45678
rect 21420 45574 21476 45612
rect 23100 45666 23156 45678
rect 23100 45614 23102 45666
rect 23154 45614 23156 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 22316 45332 22372 45342
rect 22316 45238 22372 45276
rect 21644 45220 21700 45230
rect 21644 45106 21700 45164
rect 21644 45054 21646 45106
rect 21698 45054 21700 45106
rect 20972 44996 21028 45006
rect 20972 44902 21028 44940
rect 18732 44270 18734 44322
rect 18786 44270 18788 44322
rect 18732 44258 18788 44270
rect 19068 44434 19348 44436
rect 19068 44382 19294 44434
rect 19346 44382 19348 44434
rect 19068 44380 19348 44382
rect 18620 43586 18676 43596
rect 19068 43540 19124 44380
rect 19292 44370 19348 44380
rect 21644 44324 21700 45054
rect 21644 44258 21700 44268
rect 21756 45218 21812 45230
rect 21756 45166 21758 45218
rect 21810 45166 21812 45218
rect 21756 45108 21812 45166
rect 22204 45220 22260 45230
rect 23100 45220 23156 45614
rect 22204 45126 22260 45164
rect 22876 45164 23156 45220
rect 23324 45332 23380 45342
rect 21756 44324 21812 45052
rect 21980 45106 22036 45118
rect 21980 45054 21982 45106
rect 22034 45054 22036 45106
rect 21980 44884 22036 45054
rect 22428 45108 22484 45118
rect 22428 45014 22484 45052
rect 22876 45106 22932 45164
rect 22876 45054 22878 45106
rect 22930 45054 22932 45106
rect 22204 44884 22260 44894
rect 21980 44828 22204 44884
rect 22204 44818 22260 44828
rect 22092 44324 22148 44334
rect 21756 44322 21924 44324
rect 21756 44270 21758 44322
rect 21810 44270 21924 44322
rect 21756 44268 21924 44270
rect 21756 44258 21812 44268
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19068 43446 19124 43484
rect 20188 43764 20244 43774
rect 19740 43428 19796 43438
rect 19740 43334 19796 43372
rect 18396 42914 18452 42924
rect 20188 42978 20244 43708
rect 21196 43652 21252 43662
rect 20860 43540 20916 43550
rect 20916 43484 21028 43540
rect 20860 43474 20916 43484
rect 20188 42926 20190 42978
rect 20242 42926 20244 42978
rect 20188 42914 20244 42926
rect 20300 42980 20356 42990
rect 18172 42756 18228 42766
rect 18172 42754 18564 42756
rect 18172 42702 18174 42754
rect 18226 42702 18564 42754
rect 18172 42700 18564 42702
rect 18172 42690 18228 42700
rect 18060 41458 18116 41468
rect 18284 41970 18340 41982
rect 18284 41918 18286 41970
rect 18338 41918 18340 41970
rect 17500 40350 17502 40402
rect 17554 40350 17556 40402
rect 17500 38668 17556 40350
rect 17836 41186 17892 41198
rect 17836 41134 17838 41186
rect 17890 41134 17892 41186
rect 17724 39732 17780 39742
rect 17724 39638 17780 39676
rect 17836 39730 17892 41134
rect 17948 40514 18004 40526
rect 17948 40462 17950 40514
rect 18002 40462 18004 40514
rect 17948 40404 18004 40462
rect 17948 40338 18004 40348
rect 18284 40516 18340 41918
rect 17836 39678 17838 39730
rect 17890 39678 17892 39730
rect 17836 38946 17892 39678
rect 17836 38894 17838 38946
rect 17890 38894 17892 38946
rect 17836 38882 17892 38894
rect 17500 38612 17780 38668
rect 17612 38052 17668 38062
rect 17500 37716 17556 37726
rect 17500 37490 17556 37660
rect 17500 37438 17502 37490
rect 17554 37438 17556 37490
rect 17500 37426 17556 37438
rect 17276 36542 17278 36594
rect 17330 36542 17332 36594
rect 17276 36530 17332 36542
rect 16716 34638 16718 34690
rect 16770 34638 16772 34690
rect 16716 34626 16772 34638
rect 16828 36482 16884 36494
rect 16828 36430 16830 36482
rect 16882 36430 16884 36482
rect 16828 34244 16884 36430
rect 17612 36370 17668 37996
rect 17724 37268 17780 38612
rect 17948 38164 18004 38174
rect 17948 38070 18004 38108
rect 17724 36482 17780 37212
rect 17724 36430 17726 36482
rect 17778 36430 17780 36482
rect 17724 36418 17780 36430
rect 18284 36484 18340 40460
rect 18284 36390 18340 36428
rect 18396 41300 18452 41310
rect 18396 37716 18452 41244
rect 17612 36318 17614 36370
rect 17666 36318 17668 36370
rect 17612 36306 17668 36318
rect 17388 35700 17444 35710
rect 17052 35476 17108 35486
rect 17052 35026 17108 35420
rect 17052 34974 17054 35026
rect 17106 34974 17108 35026
rect 17052 34962 17108 34974
rect 16156 34188 16884 34244
rect 16156 34130 16212 34188
rect 16156 34078 16158 34130
rect 16210 34078 16212 34130
rect 16156 34066 16212 34078
rect 16716 34018 16772 34030
rect 16716 33966 16718 34018
rect 16770 33966 16772 34018
rect 16716 33460 16772 33966
rect 16716 33394 16772 33404
rect 16716 33236 16772 33246
rect 16716 33142 16772 33180
rect 16044 32844 16212 32900
rect 16044 32676 16100 32686
rect 15932 32674 16100 32676
rect 15932 32622 16046 32674
rect 16098 32622 16100 32674
rect 15932 32620 16100 32622
rect 16044 32610 16100 32620
rect 16156 32564 16212 32844
rect 16828 32788 16884 34188
rect 16380 32564 16436 32574
rect 16156 32562 16436 32564
rect 16156 32510 16382 32562
rect 16434 32510 16436 32562
rect 16156 32508 16436 32510
rect 15484 31778 15876 31780
rect 15484 31726 15486 31778
rect 15538 31726 15876 31778
rect 15484 31724 15876 31726
rect 15036 31556 15092 31566
rect 15036 31462 15092 31500
rect 15484 31556 15540 31724
rect 14812 29986 14868 29998
rect 14812 29934 14814 29986
rect 14866 29934 14868 29986
rect 14812 29092 14868 29934
rect 15148 29428 15204 29438
rect 15148 29334 15204 29372
rect 15484 29428 15540 31500
rect 16156 31666 16212 31678
rect 16156 31614 16158 31666
rect 16210 31614 16212 31666
rect 15708 30884 15764 30894
rect 15708 30790 15764 30828
rect 16044 30324 16100 30334
rect 16156 30324 16212 31614
rect 16044 30322 16212 30324
rect 16044 30270 16046 30322
rect 16098 30270 16212 30322
rect 16044 30268 16212 30270
rect 16044 30258 16100 30268
rect 15820 29988 15876 29998
rect 15484 29362 15540 29372
rect 15596 29426 15652 29438
rect 15596 29374 15598 29426
rect 15650 29374 15652 29426
rect 15596 29316 15652 29374
rect 15596 29250 15652 29260
rect 14812 29026 14868 29036
rect 15372 29204 15428 29214
rect 14924 28756 14980 28794
rect 14924 28690 14980 28700
rect 14812 28644 14868 28654
rect 14588 28588 14756 28644
rect 14252 28420 14308 28430
rect 14588 28420 14644 28430
rect 14252 28418 14644 28420
rect 14252 28366 14254 28418
rect 14306 28366 14590 28418
rect 14642 28366 14644 28418
rect 14252 28364 14644 28366
rect 14252 28354 14308 28364
rect 14364 28196 14420 28206
rect 14420 28140 14532 28196
rect 14364 28130 14420 28140
rect 13916 28028 14196 28084
rect 14476 28082 14532 28140
rect 14476 28030 14478 28082
rect 14530 28030 14532 28082
rect 13916 27188 13972 28028
rect 14476 28018 14532 28030
rect 13916 27094 13972 27132
rect 14364 26964 14420 26974
rect 13692 26908 14084 26964
rect 13244 26238 13246 26290
rect 13298 26238 13300 26290
rect 13244 26226 13300 26238
rect 13356 26348 13524 26404
rect 12124 25506 12292 25508
rect 12124 25454 12126 25506
rect 12178 25454 12292 25506
rect 12124 25452 12292 25454
rect 12124 25442 12180 25452
rect 12236 25284 12292 25294
rect 12012 25282 12292 25284
rect 12012 25230 12238 25282
rect 12290 25230 12292 25282
rect 12012 25228 12292 25230
rect 10444 25218 10500 25228
rect 12236 25218 12292 25228
rect 12460 25282 12516 25294
rect 12460 25230 12462 25282
rect 12514 25230 12516 25282
rect 9660 25106 9716 25116
rect 10220 25172 10276 25182
rect 8876 24894 8878 24946
rect 8930 24894 8932 24946
rect 8876 24882 8932 24894
rect 10220 24722 10276 25116
rect 12460 24836 12516 25230
rect 12796 25284 12852 25294
rect 12852 25228 12964 25284
rect 12796 25190 12852 25228
rect 12460 24770 12516 24780
rect 10220 24670 10222 24722
rect 10274 24670 10276 24722
rect 10220 24658 10276 24670
rect 10892 24612 10948 24622
rect 10892 24518 10948 24556
rect 12908 16324 12964 25228
rect 13020 24612 13076 24622
rect 13356 24612 13412 26348
rect 13916 25618 13972 25630
rect 13916 25566 13918 25618
rect 13970 25566 13972 25618
rect 13916 25396 13972 25566
rect 13916 25330 13972 25340
rect 14028 25506 14084 26908
rect 14364 26870 14420 26908
rect 14588 26516 14644 28364
rect 14700 27970 14756 28588
rect 14812 28530 14868 28588
rect 15372 28642 15428 29148
rect 15820 28756 15876 29932
rect 15820 28662 15876 28700
rect 15372 28590 15374 28642
rect 15426 28590 15428 28642
rect 15372 28578 15428 28590
rect 14812 28478 14814 28530
rect 14866 28478 14868 28530
rect 14812 28466 14868 28478
rect 14924 28530 14980 28542
rect 14924 28478 14926 28530
rect 14978 28478 14980 28530
rect 14924 28084 14980 28478
rect 15708 28420 15764 28430
rect 15036 28084 15092 28094
rect 14924 28082 15092 28084
rect 14924 28030 15038 28082
rect 15090 28030 15092 28082
rect 14924 28028 15092 28030
rect 15708 28084 15764 28364
rect 15820 28084 15876 28094
rect 15708 28082 15876 28084
rect 15708 28030 15822 28082
rect 15874 28030 15876 28082
rect 15708 28028 15876 28030
rect 15036 28018 15092 28028
rect 14700 27918 14702 27970
rect 14754 27918 14756 27970
rect 14700 27860 14756 27918
rect 15260 27972 15316 27982
rect 15260 27878 15316 27916
rect 14700 27794 14756 27804
rect 14812 27858 14868 27870
rect 14812 27806 14814 27858
rect 14866 27806 14868 27858
rect 14812 27748 14868 27806
rect 15372 27858 15428 27870
rect 15372 27806 15374 27858
rect 15426 27806 15428 27858
rect 15372 27748 15428 27806
rect 14812 27692 15428 27748
rect 15708 27748 15764 27758
rect 15148 27188 15204 27198
rect 14700 27076 14756 27086
rect 14700 26982 14756 27020
rect 15148 26962 15204 27132
rect 15148 26910 15150 26962
rect 15202 26910 15204 26962
rect 15148 26898 15204 26910
rect 15260 27074 15316 27692
rect 15260 27022 15262 27074
rect 15314 27022 15316 27074
rect 15260 26964 15316 27022
rect 15260 26898 15316 26908
rect 15708 27186 15764 27692
rect 15820 27636 15876 28028
rect 15820 27570 15876 27580
rect 15708 27134 15710 27186
rect 15762 27134 15764 27186
rect 15708 26964 15764 27134
rect 15708 26898 15764 26908
rect 15932 27076 15988 27086
rect 14924 26852 14980 26862
rect 14588 26450 14644 26460
rect 14812 26850 14980 26852
rect 14812 26798 14926 26850
rect 14978 26798 14980 26850
rect 14812 26796 14980 26798
rect 14812 26068 14868 26796
rect 14924 26786 14980 26796
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 13580 25282 13636 25294
rect 13580 25230 13582 25282
rect 13634 25230 13636 25282
rect 13580 25172 13636 25230
rect 13468 25116 13580 25172
rect 13468 24946 13524 25116
rect 13580 25106 13636 25116
rect 13468 24894 13470 24946
rect 13522 24894 13524 24946
rect 13468 24882 13524 24894
rect 13020 24610 13412 24612
rect 13020 24558 13022 24610
rect 13074 24558 13412 24610
rect 13020 24556 13412 24558
rect 13804 24724 13860 24734
rect 13020 24546 13076 24556
rect 13804 23042 13860 24668
rect 14028 24722 14084 25454
rect 14364 26012 14868 26068
rect 14924 26516 14980 26526
rect 14364 25394 14420 26012
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 14364 25330 14420 25342
rect 14700 25508 14756 25518
rect 14924 25508 14980 26460
rect 15596 26516 15652 26526
rect 15596 26422 15652 26460
rect 15932 26516 15988 27020
rect 16268 26908 16324 32508
rect 16380 32498 16436 32508
rect 16828 32562 16884 32732
rect 16828 32510 16830 32562
rect 16882 32510 16884 32562
rect 16828 32498 16884 32510
rect 17388 34130 17444 35644
rect 17948 34692 18004 34702
rect 17948 34242 18004 34636
rect 17948 34190 17950 34242
rect 18002 34190 18004 34242
rect 17948 34178 18004 34190
rect 17388 34078 17390 34130
rect 17442 34078 17444 34130
rect 17388 31892 17444 34078
rect 17612 32788 17668 32798
rect 17612 32694 17668 32732
rect 18172 32788 18228 32798
rect 18172 32562 18228 32732
rect 18172 32510 18174 32562
rect 18226 32510 18228 32562
rect 18172 32498 18228 32510
rect 17276 31836 17388 31892
rect 16380 30098 16436 30110
rect 16380 30046 16382 30098
rect 16434 30046 16436 30098
rect 16380 29092 16436 30046
rect 16492 30100 16548 30110
rect 16492 30006 16548 30044
rect 17052 30100 17108 30110
rect 17052 30006 17108 30044
rect 17276 30098 17332 31836
rect 17388 31826 17444 31836
rect 18284 31890 18340 31902
rect 18284 31838 18286 31890
rect 18338 31838 18340 31890
rect 18284 31780 18340 31838
rect 18284 31714 18340 31724
rect 17276 30046 17278 30098
rect 17330 30046 17332 30098
rect 17276 30034 17332 30046
rect 17388 30100 17444 30110
rect 17388 30098 17780 30100
rect 17388 30046 17390 30098
rect 17442 30046 17780 30098
rect 17388 30044 17780 30046
rect 17388 30034 17444 30044
rect 16604 29988 16660 29998
rect 16604 29894 16660 29932
rect 16828 29988 16884 29998
rect 16828 29986 16996 29988
rect 16828 29934 16830 29986
rect 16882 29934 16996 29986
rect 16828 29932 16996 29934
rect 16828 29922 16884 29932
rect 16380 28868 16436 29036
rect 16380 28802 16436 28812
rect 16828 29316 16884 29326
rect 16604 28644 16660 28654
rect 16828 28644 16884 29260
rect 16604 28642 16884 28644
rect 16604 28590 16606 28642
rect 16658 28590 16884 28642
rect 16604 28588 16884 28590
rect 16604 28578 16660 28588
rect 16828 26908 16884 28588
rect 16940 28418 16996 29932
rect 17388 29426 17444 29438
rect 17388 29374 17390 29426
rect 17442 29374 17444 29426
rect 17388 29316 17444 29374
rect 17388 29250 17444 29260
rect 17724 28980 17780 30044
rect 17836 29988 17892 29998
rect 17836 29894 17892 29932
rect 18172 29316 18228 29326
rect 18172 29314 18340 29316
rect 18172 29262 18174 29314
rect 18226 29262 18340 29314
rect 18172 29260 18340 29262
rect 18172 29250 18228 29260
rect 17724 28924 18116 28980
rect 17612 28868 17668 28878
rect 17612 28756 17668 28812
rect 17388 28700 17668 28756
rect 17388 28642 17444 28700
rect 17388 28590 17390 28642
rect 17442 28590 17444 28642
rect 17388 28578 17444 28590
rect 18060 28642 18116 28924
rect 18172 28868 18228 28906
rect 18172 28802 18228 28812
rect 18060 28590 18062 28642
rect 18114 28590 18116 28642
rect 17500 28532 17556 28542
rect 17500 28438 17556 28476
rect 16940 28366 16942 28418
rect 16994 28366 16996 28418
rect 16940 28196 16996 28366
rect 17052 28420 17108 28430
rect 17052 28326 17108 28364
rect 17164 28418 17220 28430
rect 17164 28366 17166 28418
rect 17218 28366 17220 28418
rect 16940 28140 17108 28196
rect 16268 26852 16772 26908
rect 16828 26852 16996 26908
rect 15932 26422 15988 26460
rect 16492 26404 16548 26414
rect 16604 26404 16660 26414
rect 16492 26402 16604 26404
rect 16492 26350 16494 26402
rect 16546 26350 16604 26402
rect 16492 26348 16604 26350
rect 16492 26338 16548 26348
rect 14700 25506 14980 25508
rect 14700 25454 14702 25506
rect 14754 25454 14980 25506
rect 14700 25452 14980 25454
rect 15036 26178 15092 26190
rect 15036 26126 15038 26178
rect 15090 26126 15092 26178
rect 14476 25282 14532 25294
rect 14476 25230 14478 25282
rect 14530 25230 14532 25282
rect 14476 25060 14532 25230
rect 14476 24994 14532 25004
rect 14700 24946 14756 25452
rect 15036 25172 15092 26126
rect 15820 25620 15876 25630
rect 15820 25618 15988 25620
rect 15820 25566 15822 25618
rect 15874 25566 15988 25618
rect 15820 25564 15988 25566
rect 15820 25554 15876 25564
rect 15036 25106 15092 25116
rect 15596 25282 15652 25294
rect 15596 25230 15598 25282
rect 15650 25230 15652 25282
rect 14700 24894 14702 24946
rect 14754 24894 14756 24946
rect 14700 24882 14756 24894
rect 15148 25060 15204 25070
rect 15148 24946 15204 25004
rect 15148 24894 15150 24946
rect 15202 24894 15204 24946
rect 15148 24882 15204 24894
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 14028 24658 14084 24670
rect 14252 24836 14308 24846
rect 14252 24722 14308 24780
rect 14476 24836 14532 24846
rect 14476 24834 14644 24836
rect 14476 24782 14478 24834
rect 14530 24782 14644 24834
rect 14476 24780 14644 24782
rect 14476 24770 14532 24780
rect 14252 24670 14254 24722
rect 14306 24670 14308 24722
rect 14252 24658 14308 24670
rect 14364 24612 14420 24622
rect 14364 24518 14420 24556
rect 14588 24612 14644 24780
rect 14588 24546 14644 24556
rect 15596 24612 15652 25230
rect 15596 24518 15652 24556
rect 15820 25172 15876 25182
rect 15820 23716 15876 25116
rect 15820 23650 15876 23660
rect 15932 23266 15988 25564
rect 16604 25508 16660 26348
rect 16604 25414 16660 25452
rect 16044 25394 16100 25406
rect 16044 25342 16046 25394
rect 16098 25342 16100 25394
rect 16044 25284 16100 25342
rect 16268 25394 16324 25406
rect 16268 25342 16270 25394
rect 16322 25342 16324 25394
rect 16044 25228 16212 25284
rect 16156 24948 16212 25228
rect 16156 24854 16212 24892
rect 16268 24946 16324 25342
rect 16268 24894 16270 24946
rect 16322 24894 16324 24946
rect 16268 24882 16324 24894
rect 16380 25282 16436 25294
rect 16380 25230 16382 25282
rect 16434 25230 16436 25282
rect 16380 24612 16436 25230
rect 16716 25172 16772 26852
rect 16828 26292 16884 26302
rect 16828 26198 16884 26236
rect 16828 25508 16884 25518
rect 16940 25508 16996 26852
rect 17052 26404 17108 28140
rect 17164 28084 17220 28366
rect 17164 28018 17220 28028
rect 17612 27636 17668 27646
rect 17388 26404 17444 26414
rect 17052 26338 17108 26348
rect 17276 26348 17388 26404
rect 16828 25506 16996 25508
rect 16828 25454 16830 25506
rect 16882 25454 16996 25506
rect 16828 25452 16996 25454
rect 16828 25396 16884 25452
rect 17276 25396 17332 26348
rect 17388 26310 17444 26348
rect 16828 25330 16884 25340
rect 16940 25340 17332 25396
rect 17388 25508 17444 25518
rect 16492 25116 16772 25172
rect 16492 24834 16548 25116
rect 16940 25060 16996 25340
rect 16492 24782 16494 24834
rect 16546 24782 16548 24834
rect 16492 24724 16548 24782
rect 16604 25004 16996 25060
rect 16604 24834 16660 25004
rect 17388 24946 17444 25452
rect 17388 24894 17390 24946
rect 17442 24894 17444 24946
rect 17388 24882 17444 24894
rect 16604 24782 16606 24834
rect 16658 24782 16660 24834
rect 16604 24770 16660 24782
rect 17612 24834 17668 27580
rect 18060 26404 18116 28590
rect 18172 28644 18228 28654
rect 18172 28530 18228 28588
rect 18172 28478 18174 28530
rect 18226 28478 18228 28530
rect 18172 28466 18228 28478
rect 18284 28420 18340 29260
rect 18284 28354 18340 28364
rect 18172 28084 18228 28094
rect 18228 28028 18340 28084
rect 18172 27990 18228 28028
rect 18172 26850 18228 26862
rect 18172 26798 18174 26850
rect 18226 26798 18228 26850
rect 18172 26514 18228 26798
rect 18172 26462 18174 26514
rect 18226 26462 18228 26514
rect 18172 26450 18228 26462
rect 18060 26310 18116 26348
rect 17724 26292 17780 26302
rect 17724 25732 17780 26236
rect 18172 26068 18228 26078
rect 17724 25666 17780 25676
rect 17836 26066 18228 26068
rect 17836 26014 18174 26066
rect 18226 26014 18228 26066
rect 17836 26012 18228 26014
rect 17612 24782 17614 24834
rect 17666 24782 17668 24834
rect 16492 24658 16548 24668
rect 16380 23940 16436 24556
rect 17612 24388 17668 24782
rect 17724 25394 17780 25406
rect 17724 25342 17726 25394
rect 17778 25342 17780 25394
rect 17724 24610 17780 25342
rect 17836 24722 17892 26012
rect 18172 26002 18228 26012
rect 18284 25060 18340 28028
rect 18396 27188 18452 37660
rect 18508 37492 18564 42700
rect 19628 42754 19684 42766
rect 19628 42702 19630 42754
rect 19682 42702 19684 42754
rect 19180 42084 19236 42094
rect 18732 41970 18788 41982
rect 18732 41918 18734 41970
rect 18786 41918 18788 41970
rect 18732 41300 18788 41918
rect 18732 41234 18788 41244
rect 18732 41074 18788 41086
rect 18732 41022 18734 41074
rect 18786 41022 18788 41074
rect 18732 39732 18788 41022
rect 19180 41076 19236 42028
rect 19516 42082 19572 42094
rect 19516 42030 19518 42082
rect 19570 42030 19572 42082
rect 19516 41412 19572 42030
rect 19516 41346 19572 41356
rect 19180 40290 19236 41020
rect 19516 41186 19572 41198
rect 19516 41134 19518 41186
rect 19570 41134 19572 41186
rect 19404 40964 19460 40974
rect 19404 40404 19460 40908
rect 19404 40338 19460 40348
rect 19180 40238 19182 40290
rect 19234 40238 19236 40290
rect 18732 39618 18788 39676
rect 18732 39566 18734 39618
rect 18786 39566 18788 39618
rect 18732 39554 18788 39566
rect 18844 40180 18900 40190
rect 18844 39058 18900 40124
rect 18844 39006 18846 39058
rect 18898 39006 18900 39058
rect 18844 38994 18900 39006
rect 19180 38668 19236 40238
rect 19516 39508 19572 41134
rect 19628 40628 19684 42702
rect 20300 42642 20356 42924
rect 20300 42590 20302 42642
rect 20354 42590 20356 42642
rect 20300 42578 20356 42590
rect 20748 42642 20804 42654
rect 20748 42590 20750 42642
rect 20802 42590 20804 42642
rect 20524 42532 20580 42542
rect 20524 42530 20692 42532
rect 20524 42478 20526 42530
rect 20578 42478 20692 42530
rect 20524 42476 20692 42478
rect 20524 42466 20580 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19964 42196 20020 42206
rect 19964 41860 20020 42140
rect 19964 41766 20020 41804
rect 20300 41972 20356 41982
rect 19964 41074 20020 41086
rect 19964 41022 19966 41074
rect 20018 41022 20020 41074
rect 19964 40964 20020 41022
rect 20188 41076 20244 41086
rect 20188 40982 20244 41020
rect 19964 40898 20020 40908
rect 20300 40962 20356 41916
rect 20300 40910 20302 40962
rect 20354 40910 20356 40962
rect 20300 40898 20356 40910
rect 20412 41970 20468 41982
rect 20412 41918 20414 41970
rect 20466 41918 20468 41970
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19740 40628 19796 40638
rect 20412 40628 20468 41918
rect 20636 41636 20692 42476
rect 20748 42196 20804 42590
rect 20748 42130 20804 42140
rect 20748 41970 20804 41982
rect 20748 41918 20750 41970
rect 20802 41918 20804 41970
rect 20748 41748 20804 41918
rect 20748 41682 20804 41692
rect 20524 41300 20580 41310
rect 20524 41186 20580 41244
rect 20524 41134 20526 41186
rect 20578 41134 20580 41186
rect 20524 41122 20580 41134
rect 19628 40626 20468 40628
rect 19628 40574 19742 40626
rect 19794 40574 20468 40626
rect 19628 40572 20468 40574
rect 19740 40562 19796 40572
rect 20300 40404 20356 40414
rect 20188 39620 20244 39630
rect 20188 39526 20244 39564
rect 19628 39508 19684 39518
rect 19516 39452 19628 39508
rect 19628 39442 19684 39452
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19628 39060 19684 39070
rect 19628 38966 19684 39004
rect 20300 38948 20356 40348
rect 20412 40292 20468 40302
rect 20412 39508 20468 40236
rect 20636 39844 20692 41580
rect 20860 41636 20916 41646
rect 20636 39778 20692 39788
rect 20748 41412 20804 41422
rect 20412 39506 20580 39508
rect 20412 39454 20414 39506
rect 20466 39454 20580 39506
rect 20412 39452 20580 39454
rect 20412 39442 20468 39452
rect 20300 38882 20356 38892
rect 20524 38946 20580 39452
rect 20524 38894 20526 38946
rect 20578 38894 20580 38946
rect 20524 38882 20580 38894
rect 18956 38612 19236 38668
rect 19740 38724 19796 38734
rect 20748 38668 20804 41356
rect 20860 40402 20916 41580
rect 20860 40350 20862 40402
rect 20914 40350 20916 40402
rect 20860 40338 20916 40350
rect 20972 40068 21028 43484
rect 21084 42532 21140 42542
rect 21084 40180 21140 42476
rect 21196 42082 21252 43596
rect 21868 43426 21924 44268
rect 22092 44230 22148 44268
rect 22316 44212 22372 44222
rect 22652 44212 22708 44222
rect 22204 44210 22708 44212
rect 22204 44158 22318 44210
rect 22370 44158 22654 44210
rect 22706 44158 22708 44210
rect 22204 44156 22708 44158
rect 22204 43650 22260 44156
rect 22316 44146 22372 44156
rect 22652 44146 22708 44156
rect 22204 43598 22206 43650
rect 22258 43598 22260 43650
rect 22204 43586 22260 43598
rect 22764 44098 22820 44110
rect 22764 44046 22766 44098
rect 22818 44046 22820 44098
rect 22764 43650 22820 44046
rect 22764 43598 22766 43650
rect 22818 43598 22820 43650
rect 22764 43586 22820 43598
rect 22876 44098 22932 45054
rect 23324 45106 23380 45276
rect 23324 45054 23326 45106
rect 23378 45054 23380 45106
rect 23324 45042 23380 45054
rect 23100 44994 23156 45006
rect 23100 44942 23102 44994
rect 23154 44942 23156 44994
rect 23100 44884 23156 44942
rect 23100 44818 23156 44828
rect 22876 44046 22878 44098
rect 22930 44046 22932 44098
rect 22876 43876 22932 44046
rect 23324 44324 23380 44334
rect 23436 44324 23492 48076
rect 23772 48130 23828 48142
rect 23772 48078 23774 48130
rect 23826 48078 23828 48130
rect 23772 48020 23828 48078
rect 23772 47954 23828 47964
rect 23660 47460 23716 47470
rect 23660 47366 23716 47404
rect 23884 47348 23940 49756
rect 25116 49140 25172 50428
rect 25116 49074 25172 49084
rect 24444 48804 24500 48814
rect 24444 48466 24500 48748
rect 24444 48414 24446 48466
rect 24498 48414 24500 48466
rect 24332 48018 24388 48030
rect 24332 47966 24334 48018
rect 24386 47966 24388 48018
rect 24332 47572 24388 47966
rect 24332 47506 24388 47516
rect 23996 47348 24052 47358
rect 23884 47346 24052 47348
rect 23884 47294 23998 47346
rect 24050 47294 24052 47346
rect 23884 47292 24052 47294
rect 23996 47282 24052 47292
rect 23660 47236 23716 47246
rect 23660 46786 23716 47180
rect 24332 47234 24388 47246
rect 24332 47182 24334 47234
rect 24386 47182 24388 47234
rect 24332 47124 24388 47182
rect 24444 47236 24500 48414
rect 24668 48020 24724 48030
rect 24668 47684 24724 47964
rect 24668 47628 24948 47684
rect 24556 47460 24612 47470
rect 24556 47366 24612 47404
rect 24892 47346 24948 47628
rect 24892 47294 24894 47346
rect 24946 47294 24948 47346
rect 24780 47236 24836 47246
rect 24444 47234 24836 47236
rect 24444 47182 24782 47234
rect 24834 47182 24836 47234
rect 24444 47180 24836 47182
rect 24780 47170 24836 47180
rect 24892 47236 24948 47294
rect 24892 47170 24948 47180
rect 25452 47234 25508 47246
rect 25452 47182 25454 47234
rect 25506 47182 25508 47234
rect 23660 46734 23662 46786
rect 23714 46734 23716 46786
rect 23660 46722 23716 46734
rect 23996 47068 24332 47124
rect 23548 46676 23604 46686
rect 23548 46582 23604 46620
rect 23660 46340 23716 46350
rect 23660 45330 23716 46284
rect 23660 45278 23662 45330
rect 23714 45278 23716 45330
rect 23660 45266 23716 45278
rect 23324 44322 23492 44324
rect 23324 44270 23326 44322
rect 23378 44270 23492 44322
rect 23324 44268 23492 44270
rect 23324 44212 23380 44268
rect 23212 43988 23268 43998
rect 23212 43876 23268 43932
rect 22876 43820 23268 43876
rect 21868 43374 21870 43426
rect 21922 43374 21924 43426
rect 21868 43362 21924 43374
rect 22092 43540 22148 43550
rect 22092 42866 22148 43484
rect 22540 43538 22596 43550
rect 22540 43486 22542 43538
rect 22594 43486 22596 43538
rect 22316 43428 22372 43438
rect 22540 43428 22596 43486
rect 22876 43428 22932 43820
rect 23212 43762 23268 43820
rect 23212 43710 23214 43762
rect 23266 43710 23268 43762
rect 23212 43698 23268 43710
rect 22540 43372 22932 43428
rect 22316 43334 22372 43372
rect 22092 42814 22094 42866
rect 22146 42814 22148 42866
rect 22092 42802 22148 42814
rect 21308 42644 21364 42654
rect 21308 42550 21364 42588
rect 21644 42644 21700 42654
rect 21644 42642 21812 42644
rect 21644 42590 21646 42642
rect 21698 42590 21812 42642
rect 21644 42588 21812 42590
rect 21644 42578 21700 42588
rect 21532 42532 21588 42542
rect 21532 42196 21588 42476
rect 21532 42140 21700 42196
rect 21196 42030 21198 42082
rect 21250 42030 21252 42082
rect 21196 42018 21252 42030
rect 21644 42082 21700 42140
rect 21644 42030 21646 42082
rect 21698 42030 21700 42082
rect 21644 42018 21700 42030
rect 21532 41972 21588 41982
rect 21420 41970 21588 41972
rect 21420 41918 21534 41970
rect 21586 41918 21588 41970
rect 21420 41916 21588 41918
rect 21308 41524 21364 41534
rect 21196 41412 21252 41422
rect 21196 40514 21252 41356
rect 21308 41298 21364 41468
rect 21308 41246 21310 41298
rect 21362 41246 21364 41298
rect 21308 41234 21364 41246
rect 21196 40462 21198 40514
rect 21250 40462 21252 40514
rect 21196 40450 21252 40462
rect 21308 40516 21364 40526
rect 21308 40422 21364 40460
rect 21308 40180 21364 40190
rect 21084 40178 21364 40180
rect 21084 40126 21310 40178
rect 21362 40126 21364 40178
rect 21084 40124 21364 40126
rect 21308 40114 21364 40124
rect 18844 38164 18900 38174
rect 18508 37426 18564 37436
rect 18620 37604 18676 37614
rect 18508 35700 18564 35710
rect 18508 35606 18564 35644
rect 18620 35586 18676 37548
rect 18844 37266 18900 38108
rect 18844 37214 18846 37266
rect 18898 37214 18900 37266
rect 18844 36482 18900 37214
rect 18844 36430 18846 36482
rect 18898 36430 18900 36482
rect 18844 35810 18900 36430
rect 18844 35758 18846 35810
rect 18898 35758 18900 35810
rect 18844 35700 18900 35758
rect 18844 35634 18900 35644
rect 18620 35534 18622 35586
rect 18674 35534 18676 35586
rect 18620 35522 18676 35534
rect 18620 33236 18676 33246
rect 18620 32786 18676 33180
rect 18620 32734 18622 32786
rect 18674 32734 18676 32786
rect 18620 32722 18676 32734
rect 18844 32676 18900 32686
rect 18844 32582 18900 32620
rect 18508 32564 18564 32574
rect 18508 32470 18564 32508
rect 18620 31892 18676 31902
rect 18620 31798 18676 31836
rect 18956 30212 19012 38612
rect 19404 38388 19460 38398
rect 19404 36484 19460 38332
rect 19292 36482 19460 36484
rect 19292 36430 19406 36482
rect 19458 36430 19460 36482
rect 19292 36428 19460 36430
rect 19292 34354 19348 36428
rect 19404 36418 19460 36428
rect 19628 38276 19684 38286
rect 19628 36370 19684 38220
rect 19740 38162 19796 38668
rect 19740 38110 19742 38162
rect 19794 38110 19796 38162
rect 19740 38098 19796 38110
rect 20300 38612 20804 38668
rect 20860 40012 21028 40068
rect 20188 38052 20244 38062
rect 20188 37958 20244 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20300 37492 20356 38612
rect 19628 36318 19630 36370
rect 19682 36318 19684 36370
rect 19628 36306 19684 36318
rect 20188 37436 20356 37492
rect 20636 37828 20692 37838
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19964 35700 20020 35710
rect 20020 35644 20132 35700
rect 19964 35634 20020 35644
rect 20076 35026 20132 35644
rect 20076 34974 20078 35026
rect 20130 34974 20132 35026
rect 20076 34962 20132 34974
rect 19516 34692 19572 34702
rect 19292 34302 19294 34354
rect 19346 34302 19348 34354
rect 19292 34290 19348 34302
rect 19404 34690 19572 34692
rect 19404 34638 19518 34690
rect 19570 34638 19572 34690
rect 19404 34636 19572 34638
rect 19180 34020 19236 34030
rect 19068 33124 19124 33134
rect 19068 32674 19124 33068
rect 19068 32622 19070 32674
rect 19122 32622 19124 32674
rect 19068 32610 19124 32622
rect 19068 30212 19124 30222
rect 18956 30210 19124 30212
rect 18956 30158 19070 30210
rect 19122 30158 19124 30210
rect 18956 30156 19124 30158
rect 18844 29092 18900 29102
rect 18620 28532 18676 28542
rect 18620 27746 18676 28476
rect 18844 28530 18900 29036
rect 18956 28644 19012 30156
rect 19068 30146 19124 30156
rect 19180 29988 19236 33964
rect 19404 33458 19460 34636
rect 19516 34626 19572 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19404 33406 19406 33458
rect 19458 33406 19460 33458
rect 19404 32788 19460 33406
rect 20188 33346 20244 37436
rect 20300 37268 20356 37278
rect 20300 37174 20356 37212
rect 20412 37156 20468 37166
rect 20300 36484 20356 36494
rect 20300 35698 20356 36428
rect 20300 35646 20302 35698
rect 20354 35646 20356 35698
rect 20300 34354 20356 35646
rect 20300 34302 20302 34354
rect 20354 34302 20356 34354
rect 20300 34290 20356 34302
rect 20412 34132 20468 37100
rect 20636 37044 20692 37772
rect 20636 36950 20692 36988
rect 20748 36260 20804 36270
rect 20748 35812 20804 36204
rect 20860 35924 20916 40012
rect 21084 39844 21140 39854
rect 20972 38834 21028 38846
rect 20972 38782 20974 38834
rect 21026 38782 21028 38834
rect 20972 37940 21028 38782
rect 21084 38668 21140 39788
rect 21196 39620 21252 39630
rect 21196 38836 21252 39564
rect 21308 39508 21364 39518
rect 21308 39414 21364 39452
rect 21308 38836 21364 38846
rect 21196 38780 21308 38836
rect 21308 38742 21364 38780
rect 21084 38612 21252 38668
rect 21196 38162 21252 38612
rect 21420 38276 21476 41916
rect 21532 41906 21588 41916
rect 21756 40628 21812 42588
rect 22652 42084 22708 42094
rect 22316 41972 22372 41982
rect 22316 41300 22372 41916
rect 22540 41858 22596 41870
rect 22540 41806 22542 41858
rect 22594 41806 22596 41858
rect 22540 41746 22596 41806
rect 22540 41694 22542 41746
rect 22594 41694 22596 41746
rect 22540 41300 22596 41694
rect 21868 41298 22484 41300
rect 21868 41246 22318 41298
rect 22370 41246 22484 41298
rect 21868 41244 22484 41246
rect 21868 41186 21924 41244
rect 22316 41234 22372 41244
rect 21868 41134 21870 41186
rect 21922 41134 21924 41186
rect 21868 41122 21924 41134
rect 21532 40572 21812 40628
rect 21532 38388 21588 40572
rect 21868 40404 21924 40414
rect 21532 38322 21588 38332
rect 21644 39506 21700 39518
rect 21644 39454 21646 39506
rect 21698 39454 21700 39506
rect 21420 38210 21476 38220
rect 21196 38110 21198 38162
rect 21250 38110 21252 38162
rect 21196 38098 21252 38110
rect 21308 38164 21364 38174
rect 21308 38050 21364 38108
rect 21308 37998 21310 38050
rect 21362 37998 21364 38050
rect 21308 37986 21364 37998
rect 20972 37156 21028 37884
rect 21532 37938 21588 37950
rect 21532 37886 21534 37938
rect 21586 37886 21588 37938
rect 21532 37604 21588 37886
rect 21644 37828 21700 39454
rect 21644 37762 21700 37772
rect 21756 38836 21812 38846
rect 21756 37604 21812 38780
rect 21868 38276 21924 40348
rect 22316 40180 22372 40190
rect 21868 38210 21924 38220
rect 22204 40178 22372 40180
rect 22204 40126 22318 40178
rect 22370 40126 22372 40178
rect 22204 40124 22372 40126
rect 22204 39618 22260 40124
rect 22316 40114 22372 40124
rect 22204 39566 22206 39618
rect 22258 39566 22260 39618
rect 22092 37940 22148 37950
rect 22092 37846 22148 37884
rect 21532 37548 21812 37604
rect 20972 37090 21028 37100
rect 21196 37268 21252 37278
rect 21196 37154 21252 37212
rect 21196 37102 21198 37154
rect 21250 37102 21252 37154
rect 21196 37090 21252 37102
rect 21420 37266 21476 37278
rect 21420 37214 21422 37266
rect 21474 37214 21476 37266
rect 21308 36260 21364 36270
rect 21308 36166 21364 36204
rect 20860 35868 21364 35924
rect 20748 35746 20804 35756
rect 21084 35700 21140 35710
rect 20860 35698 21140 35700
rect 20860 35646 21086 35698
rect 21138 35646 21140 35698
rect 20860 35644 21140 35646
rect 20860 35252 20916 35644
rect 21084 35634 21140 35644
rect 20748 35196 20916 35252
rect 20748 34132 20804 35196
rect 21308 34916 21364 35868
rect 20860 34914 21364 34916
rect 20860 34862 21310 34914
rect 21362 34862 21364 34914
rect 20860 34860 21364 34862
rect 20860 34802 20916 34860
rect 21308 34850 21364 34860
rect 20860 34750 20862 34802
rect 20914 34750 20916 34802
rect 20860 34738 20916 34750
rect 20188 33294 20190 33346
rect 20242 33294 20244 33346
rect 19964 33124 20020 33134
rect 19404 32694 19460 32732
rect 19628 33122 20020 33124
rect 19628 33070 19966 33122
rect 20018 33070 20020 33122
rect 19628 33068 20020 33070
rect 19628 32564 19684 33068
rect 19964 33058 20020 33068
rect 20076 33124 20132 33162
rect 20076 33058 20132 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32788 20244 33294
rect 19628 32004 19684 32508
rect 19964 32732 20244 32788
rect 20300 34076 20468 34132
rect 20524 34130 20804 34132
rect 20524 34078 20750 34130
rect 20802 34078 20804 34130
rect 20524 34076 20804 34078
rect 20300 32788 20356 34076
rect 20412 32788 20468 32798
rect 20300 32786 20468 32788
rect 20300 32734 20414 32786
rect 20466 32734 20468 32786
rect 20300 32732 20468 32734
rect 19964 32676 20020 32732
rect 20412 32722 20468 32732
rect 19964 32562 20020 32620
rect 19964 32510 19966 32562
rect 20018 32510 20020 32562
rect 19964 32498 20020 32510
rect 20300 32450 20356 32462
rect 20300 32398 20302 32450
rect 20354 32398 20356 32450
rect 19852 32004 19908 32014
rect 19628 31948 19852 32004
rect 19852 31890 19908 31948
rect 19852 31838 19854 31890
rect 19906 31838 19908 31890
rect 19852 31826 19908 31838
rect 19404 31780 19460 31790
rect 19404 31686 19460 31724
rect 20300 31780 20356 32398
rect 20300 31714 20356 31724
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20300 30884 20356 30894
rect 20188 30828 20300 30884
rect 19628 30212 19684 30222
rect 19628 30118 19684 30156
rect 18956 28578 19012 28588
rect 19068 29932 19236 29988
rect 18844 28478 18846 28530
rect 18898 28478 18900 28530
rect 18844 28466 18900 28478
rect 18620 27694 18622 27746
rect 18674 27694 18676 27746
rect 18620 27636 18676 27694
rect 18620 27570 18676 27580
rect 18508 27188 18564 27198
rect 18396 27186 18564 27188
rect 18396 27134 18510 27186
rect 18562 27134 18564 27186
rect 18396 27132 18564 27134
rect 18396 26850 18452 27132
rect 18508 26908 18564 27132
rect 19068 26908 19124 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19628 28868 19684 28878
rect 19628 28756 19684 28812
rect 19180 28754 19684 28756
rect 19180 28702 19630 28754
rect 19682 28702 19684 28754
rect 19180 28700 19684 28702
rect 19180 28642 19236 28700
rect 19628 28690 19684 28700
rect 19180 28590 19182 28642
rect 19234 28590 19236 28642
rect 19180 28578 19236 28590
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 27860 19684 27870
rect 19292 27636 19348 27646
rect 18508 26852 18676 26908
rect 19068 26852 19236 26908
rect 18396 26798 18398 26850
rect 18450 26798 18452 26850
rect 18396 26786 18452 26798
rect 18620 26402 18676 26852
rect 18620 26350 18622 26402
rect 18674 26350 18676 26402
rect 18620 26338 18676 26350
rect 19180 26290 19236 26852
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 19180 25620 19236 26238
rect 19180 25554 19236 25564
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 24658 17892 24670
rect 18172 24948 18228 24958
rect 18172 24722 18228 24892
rect 18172 24670 18174 24722
rect 18226 24670 18228 24722
rect 18172 24658 18228 24670
rect 17724 24558 17726 24610
rect 17778 24558 17780 24610
rect 17724 24546 17780 24558
rect 17612 24322 17668 24332
rect 16380 23874 16436 23884
rect 16604 23716 16660 23726
rect 18284 23716 18340 25004
rect 19180 24948 19236 24958
rect 19292 24948 19348 27580
rect 19236 24892 19348 24948
rect 19180 24854 19236 24892
rect 19628 24724 19684 27804
rect 20188 26908 20244 30828
rect 20300 30818 20356 30828
rect 20524 30212 20580 34076
rect 20748 34066 20804 34076
rect 21420 34132 21476 37214
rect 21532 35476 21588 37548
rect 22204 36932 22260 39566
rect 22428 38612 22484 41244
rect 22540 41234 22596 41244
rect 22428 38546 22484 38556
rect 22540 40628 22596 40638
rect 22652 40628 22708 42028
rect 22876 41858 22932 41870
rect 22876 41806 22878 41858
rect 22930 41806 22932 41858
rect 22876 41746 22932 41806
rect 22876 41694 22878 41746
rect 22930 41694 22932 41746
rect 22876 41682 22932 41694
rect 23324 41636 23380 44156
rect 23660 44098 23716 44110
rect 23660 44046 23662 44098
rect 23714 44046 23716 44098
rect 23660 43988 23716 44046
rect 23660 43922 23716 43932
rect 23660 42084 23716 42122
rect 23660 42018 23716 42028
rect 23772 42084 23828 42094
rect 23772 42082 23940 42084
rect 23772 42030 23774 42082
rect 23826 42030 23940 42082
rect 23772 42028 23940 42030
rect 23772 42018 23828 42028
rect 23660 41860 23716 41870
rect 23660 41746 23716 41804
rect 23660 41694 23662 41746
rect 23714 41694 23716 41746
rect 23660 41682 23716 41694
rect 23324 41524 23380 41580
rect 23436 41524 23492 41534
rect 23324 41468 23436 41524
rect 23436 41458 23492 41468
rect 23772 41412 23828 41422
rect 22540 40626 22708 40628
rect 22540 40574 22542 40626
rect 22594 40574 22708 40626
rect 22540 40572 22708 40574
rect 23324 41298 23380 41310
rect 23324 41246 23326 41298
rect 23378 41246 23380 41298
rect 22204 36866 22260 36876
rect 22540 36596 22596 40572
rect 22988 40404 23044 40414
rect 22652 40292 22708 40302
rect 22988 40292 23044 40348
rect 22652 40290 23044 40292
rect 22652 40238 22654 40290
rect 22706 40238 23044 40290
rect 22652 40236 23044 40238
rect 22652 40226 22708 40236
rect 22652 39732 22708 39742
rect 23324 39732 23380 41246
rect 23772 41298 23828 41356
rect 23772 41246 23774 41298
rect 23826 41246 23828 41298
rect 23772 41234 23828 41246
rect 23436 41188 23492 41198
rect 23436 40964 23492 41132
rect 23436 40908 23716 40964
rect 23436 40740 23492 40750
rect 23436 40290 23492 40684
rect 23436 40238 23438 40290
rect 23490 40238 23492 40290
rect 23436 40226 23492 40238
rect 23436 39732 23492 39742
rect 23324 39676 23436 39732
rect 23660 39732 23716 40908
rect 23772 40404 23828 40414
rect 23884 40404 23940 42028
rect 23996 41972 24052 47068
rect 24332 47058 24388 47068
rect 25452 47124 25508 47182
rect 25452 47058 25508 47068
rect 24556 46900 24612 46910
rect 24556 46806 24612 46844
rect 24444 46676 24500 46686
rect 24108 46674 24500 46676
rect 24108 46622 24446 46674
rect 24498 46622 24500 46674
rect 24108 46620 24500 46622
rect 24108 45330 24164 46620
rect 24444 46610 24500 46620
rect 25228 46676 25284 46686
rect 24108 45278 24110 45330
rect 24162 45278 24164 45330
rect 24108 45266 24164 45278
rect 25228 45218 25284 46620
rect 25228 45166 25230 45218
rect 25282 45166 25284 45218
rect 25228 45154 25284 45166
rect 24780 45108 24836 45118
rect 24668 44994 24724 45006
rect 24668 44942 24670 44994
rect 24722 44942 24724 44994
rect 24444 44882 24500 44894
rect 24444 44830 24446 44882
rect 24498 44830 24500 44882
rect 24444 44324 24500 44830
rect 24108 44212 24164 44222
rect 24108 44118 24164 44156
rect 24444 44210 24500 44268
rect 24444 44158 24446 44210
rect 24498 44158 24500 44210
rect 24444 44146 24500 44158
rect 24668 44212 24724 44942
rect 24780 44322 24836 45052
rect 24780 44270 24782 44322
rect 24834 44270 24836 44322
rect 24780 44258 24836 44270
rect 25340 45108 25396 45118
rect 24668 44146 24724 44156
rect 25340 42866 25396 45052
rect 25564 44212 25620 44222
rect 25564 44118 25620 44156
rect 25340 42814 25342 42866
rect 25394 42814 25396 42866
rect 25340 42802 25396 42814
rect 23996 41906 24052 41916
rect 24780 42754 24836 42766
rect 24780 42702 24782 42754
rect 24834 42702 24836 42754
rect 24780 41300 24836 42702
rect 25004 42642 25060 42654
rect 25004 42590 25006 42642
rect 25058 42590 25060 42642
rect 25004 41636 25060 42590
rect 25116 41970 25172 41982
rect 25116 41918 25118 41970
rect 25170 41918 25172 41970
rect 25116 41860 25172 41918
rect 25116 41794 25172 41804
rect 25676 41746 25732 56812
rect 26124 56802 26180 56812
rect 26236 55468 26292 58156
rect 26460 57650 26516 57662
rect 26460 57598 26462 57650
rect 26514 57598 26516 57650
rect 26460 57428 26516 57598
rect 27020 57652 27076 58492
rect 27356 58482 27412 58492
rect 27020 57650 27300 57652
rect 27020 57598 27022 57650
rect 27074 57598 27300 57650
rect 27020 57596 27300 57598
rect 27020 57586 27076 57596
rect 26460 57362 26516 57372
rect 27244 57090 27300 57596
rect 27244 57038 27246 57090
rect 27298 57038 27300 57090
rect 27244 57026 27300 57038
rect 26684 56868 26740 56878
rect 26684 56774 26740 56812
rect 26796 56756 26852 56766
rect 27132 56756 27188 56766
rect 26796 56754 27188 56756
rect 26796 56702 26798 56754
rect 26850 56702 27134 56754
rect 27186 56702 27188 56754
rect 26796 56700 27188 56702
rect 26796 56690 26852 56700
rect 27132 56690 27188 56700
rect 27468 56532 27524 59052
rect 27804 59042 27860 59052
rect 27804 58434 27860 58446
rect 27804 58382 27806 58434
rect 27858 58382 27860 58434
rect 27804 57876 27860 58382
rect 28140 58322 28196 61180
rect 28364 60786 28420 60798
rect 28364 60734 28366 60786
rect 28418 60734 28420 60786
rect 28364 60228 28420 60734
rect 28364 60134 28420 60172
rect 28140 58270 28142 58322
rect 28194 58270 28196 58322
rect 28140 58258 28196 58270
rect 28028 57876 28084 57886
rect 27804 57874 28084 57876
rect 27804 57822 28030 57874
rect 28082 57822 28084 57874
rect 27804 57820 28084 57822
rect 28028 57810 28084 57820
rect 27692 57764 27748 57774
rect 27692 57670 27748 57708
rect 28252 57652 28308 57662
rect 28252 57558 28308 57596
rect 25900 55412 26292 55468
rect 27132 56476 27524 56532
rect 27692 56868 27748 56878
rect 27692 56642 27748 56812
rect 27692 56590 27694 56642
rect 27746 56590 27748 56642
rect 25788 49138 25844 49150
rect 25788 49086 25790 49138
rect 25842 49086 25844 49138
rect 25788 48804 25844 49086
rect 25788 48738 25844 48748
rect 25788 47570 25844 47582
rect 25788 47518 25790 47570
rect 25842 47518 25844 47570
rect 25788 46676 25844 47518
rect 25900 47124 25956 55412
rect 27020 55076 27076 55086
rect 26684 54628 26740 54638
rect 26684 54534 26740 54572
rect 27020 54626 27076 55020
rect 27020 54574 27022 54626
rect 27074 54574 27076 54626
rect 27020 54562 27076 54574
rect 26796 54402 26852 54414
rect 26796 54350 26798 54402
rect 26850 54350 26852 54402
rect 26796 54180 26852 54350
rect 26012 54124 26852 54180
rect 26012 53842 26068 54124
rect 26012 53790 26014 53842
rect 26066 53790 26068 53842
rect 26012 53778 26068 53790
rect 26236 50484 26292 50494
rect 26236 50390 26292 50428
rect 27132 49700 27188 56476
rect 27692 55300 27748 56590
rect 28476 56308 28532 62860
rect 28588 62850 28644 62860
rect 28924 62916 28980 62926
rect 28924 62466 28980 62860
rect 29036 62578 29092 63756
rect 29036 62526 29038 62578
rect 29090 62526 29092 62578
rect 29036 62514 29092 62526
rect 28924 62414 28926 62466
rect 28978 62414 28980 62466
rect 28924 62402 28980 62414
rect 29148 62354 29204 64652
rect 29484 64708 29540 64718
rect 29484 64614 29540 64652
rect 30380 64708 30436 64718
rect 30380 64614 30436 64652
rect 30940 64596 30996 64606
rect 30940 64502 30996 64540
rect 32508 64594 32564 64764
rect 32508 64542 32510 64594
rect 32562 64542 32564 64594
rect 29596 64482 29652 64494
rect 29596 64430 29598 64482
rect 29650 64430 29652 64482
rect 29596 63364 29652 64430
rect 29148 62302 29150 62354
rect 29202 62302 29204 62354
rect 29148 62290 29204 62302
rect 29372 63308 29652 63364
rect 29708 64482 29764 64494
rect 29708 64430 29710 64482
rect 29762 64430 29764 64482
rect 29372 62354 29428 63308
rect 29484 63026 29540 63038
rect 29484 62974 29486 63026
rect 29538 62974 29540 63026
rect 29484 62916 29540 62974
rect 29708 62916 29764 64430
rect 30828 64482 30884 64494
rect 30828 64430 30830 64482
rect 30882 64430 30884 64482
rect 30828 63812 30884 64430
rect 31052 64484 31108 64494
rect 31500 64484 31556 64494
rect 32284 64484 32340 64494
rect 31052 64482 31556 64484
rect 31052 64430 31054 64482
rect 31106 64430 31502 64482
rect 31554 64430 31556 64482
rect 31052 64428 31556 64430
rect 30940 63812 30996 63822
rect 30828 63810 30996 63812
rect 30828 63758 30942 63810
rect 30994 63758 30996 63810
rect 30828 63756 30996 63758
rect 30156 63140 30212 63150
rect 30156 63046 30212 63084
rect 30380 63138 30436 63150
rect 30380 63086 30382 63138
rect 30434 63086 30436 63138
rect 29540 62860 29764 62916
rect 29484 62822 29540 62860
rect 29372 62302 29374 62354
rect 29426 62302 29428 62354
rect 29372 62290 29428 62302
rect 29484 62356 29540 62366
rect 29484 62188 29540 62300
rect 30380 62244 30436 63086
rect 30940 63140 30996 63756
rect 30940 63074 30996 63084
rect 31052 63028 31108 64428
rect 31500 64418 31556 64428
rect 32172 64482 32340 64484
rect 32172 64430 32286 64482
rect 32338 64430 32340 64482
rect 32172 64428 32340 64430
rect 31948 64034 32004 64046
rect 31948 63982 31950 64034
rect 32002 63982 32004 64034
rect 31724 63812 31780 63822
rect 31724 63718 31780 63756
rect 31948 63588 32004 63982
rect 31948 63522 32004 63532
rect 32060 63922 32116 63934
rect 32060 63870 32062 63922
rect 32114 63870 32116 63922
rect 31276 63364 31332 63374
rect 31276 63270 31332 63308
rect 31948 63364 32004 63374
rect 31276 63140 31332 63150
rect 31164 63028 31220 63038
rect 31052 63026 31220 63028
rect 31052 62974 31166 63026
rect 31218 62974 31220 63026
rect 31052 62972 31220 62974
rect 30828 62244 30884 62254
rect 31164 62244 31220 62972
rect 31276 63026 31332 63084
rect 31276 62974 31278 63026
rect 31330 62974 31332 63026
rect 31276 62962 31332 62974
rect 31948 63026 32004 63308
rect 32060 63250 32116 63870
rect 32060 63198 32062 63250
rect 32114 63198 32116 63250
rect 32060 63186 32116 63198
rect 32172 63138 32228 64428
rect 32284 64418 32340 64428
rect 32508 64260 32564 64542
rect 32284 64204 32564 64260
rect 32620 64594 32676 64606
rect 32620 64542 32622 64594
rect 32674 64542 32676 64594
rect 32284 64146 32340 64204
rect 32284 64094 32286 64146
rect 32338 64094 32340 64146
rect 32284 64082 32340 64094
rect 32284 63924 32340 63934
rect 32508 63924 32564 63934
rect 32620 63924 32676 64542
rect 32956 64596 33012 64606
rect 32956 64502 33012 64540
rect 32340 63868 32452 63924
rect 32284 63858 32340 63868
rect 32172 63086 32174 63138
rect 32226 63086 32228 63138
rect 32172 63074 32228 63086
rect 32396 63138 32452 63868
rect 32396 63086 32398 63138
rect 32450 63086 32452 63138
rect 32396 63074 32452 63086
rect 32564 63868 32676 63924
rect 33068 64482 33124 64494
rect 33068 64430 33070 64482
rect 33122 64430 33124 64482
rect 31948 62974 31950 63026
rect 32002 62974 32004 63026
rect 31948 62962 32004 62974
rect 32508 62580 32564 63868
rect 32844 63588 32900 63598
rect 32844 62916 32900 63532
rect 33068 63364 33124 64430
rect 33292 64484 33348 64494
rect 33292 64390 33348 64428
rect 33180 63924 33236 63934
rect 33180 63810 33236 63868
rect 33516 63922 33572 64764
rect 33516 63870 33518 63922
rect 33570 63870 33572 63922
rect 33516 63858 33572 63870
rect 33180 63758 33182 63810
rect 33234 63758 33236 63810
rect 33180 63746 33236 63758
rect 33068 63298 33124 63308
rect 32844 62914 33012 62916
rect 32844 62862 32846 62914
rect 32898 62862 33012 62914
rect 32844 62860 33012 62862
rect 32844 62850 32900 62860
rect 32284 62524 32564 62580
rect 31276 62244 31332 62254
rect 30380 62242 31332 62244
rect 30380 62190 30830 62242
rect 30882 62190 31278 62242
rect 31330 62190 31332 62242
rect 30380 62188 31332 62190
rect 29484 62132 29764 62188
rect 29596 61124 29652 61134
rect 29596 60898 29652 61068
rect 29596 60846 29598 60898
rect 29650 60846 29652 60898
rect 29596 60834 29652 60846
rect 28924 60788 28980 60798
rect 28980 60732 29092 60788
rect 28924 60694 28980 60732
rect 28700 60676 28756 60686
rect 28700 60582 28756 60620
rect 29036 60002 29092 60732
rect 29036 59950 29038 60002
rect 29090 59950 29092 60002
rect 29036 59938 29092 59950
rect 29260 60228 29316 60238
rect 29260 59890 29316 60172
rect 29372 60004 29428 60014
rect 29372 59910 29428 59948
rect 29260 59838 29262 59890
rect 29314 59838 29316 59890
rect 29260 59826 29316 59838
rect 29708 58100 29764 62132
rect 30044 60676 30100 60686
rect 30044 60582 30100 60620
rect 30492 60676 30548 60686
rect 30492 60582 30548 60620
rect 30828 60676 30884 62188
rect 31276 62178 31332 62188
rect 30828 60610 30884 60620
rect 31052 61348 31108 61358
rect 29932 60564 29988 60574
rect 29932 60470 29988 60508
rect 30380 59892 30436 59902
rect 30380 59778 30436 59836
rect 30380 59726 30382 59778
rect 30434 59726 30436 59778
rect 30380 59556 30436 59726
rect 30380 59490 30436 59500
rect 30716 59778 30772 59790
rect 30716 59726 30718 59778
rect 30770 59726 30772 59778
rect 30716 59108 30772 59726
rect 31052 59780 31108 61292
rect 32284 61010 32340 62524
rect 32956 62244 33012 62860
rect 33852 62188 33908 65436
rect 34860 65492 34916 65550
rect 34860 65426 34916 65436
rect 35532 65492 35588 65502
rect 35532 65398 35588 65436
rect 36652 65490 36708 65502
rect 36652 65438 36654 65490
rect 36706 65438 36708 65490
rect 34972 65380 35028 65390
rect 34972 65286 35028 65324
rect 35644 65380 35700 65390
rect 35084 65266 35140 65278
rect 35084 65214 35086 65266
rect 35138 65214 35140 65266
rect 34636 64484 34692 64494
rect 34636 63922 34692 64428
rect 35084 64036 35140 65214
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35644 64818 35700 65324
rect 35644 64766 35646 64818
rect 35698 64766 35700 64818
rect 35644 64754 35700 64766
rect 36428 64708 36484 64718
rect 36652 64708 36708 65438
rect 37436 65378 37492 65390
rect 37436 65326 37438 65378
rect 37490 65326 37492 65378
rect 37436 65268 37492 65326
rect 37436 65202 37492 65212
rect 38556 65380 38612 65390
rect 36428 64706 36652 64708
rect 36428 64654 36430 64706
rect 36482 64654 36652 64706
rect 36428 64652 36652 64654
rect 36428 64642 36484 64652
rect 36652 64642 36708 64652
rect 37100 64708 37156 64718
rect 37100 64614 37156 64652
rect 38556 64708 38612 65324
rect 38556 64614 38612 64652
rect 39228 64594 39284 64606
rect 39228 64542 39230 64594
rect 39282 64542 39284 64594
rect 39228 64148 39284 64542
rect 39228 64082 39284 64092
rect 35196 64036 35252 64046
rect 35084 64034 35252 64036
rect 35084 63982 35198 64034
rect 35250 63982 35252 64034
rect 35084 63980 35252 63982
rect 35196 63970 35252 63980
rect 34636 63870 34638 63922
rect 34690 63870 34692 63922
rect 34636 63858 34692 63870
rect 39340 63924 39396 66220
rect 39564 66274 39844 66276
rect 39564 66222 39790 66274
rect 39842 66222 39844 66274
rect 39564 66220 39844 66222
rect 39564 65378 39620 66220
rect 39788 66210 39844 66220
rect 41020 65492 41076 69200
rect 43036 67172 43092 69200
rect 43036 67116 43876 67172
rect 43820 66498 43876 67116
rect 43820 66446 43822 66498
rect 43874 66446 43876 66498
rect 43820 66434 43876 66446
rect 45052 66500 45108 69200
rect 47068 67228 47124 69200
rect 47068 67172 47572 67228
rect 45052 66434 45108 66444
rect 46172 66274 46228 66286
rect 46172 66222 46174 66274
rect 46226 66222 46228 66274
rect 43036 66164 43092 66174
rect 43036 66070 43092 66108
rect 46172 66164 46228 66222
rect 41020 65426 41076 65436
rect 42700 65492 42756 65502
rect 39564 65326 39566 65378
rect 39618 65326 39620 65378
rect 39564 65314 39620 65326
rect 40124 65378 40180 65390
rect 40124 65326 40126 65378
rect 40178 65326 40180 65378
rect 40124 65268 40180 65326
rect 41132 65380 41188 65390
rect 41132 65286 41188 65324
rect 41580 65380 41636 65390
rect 42028 65380 42084 65390
rect 41580 65378 41860 65380
rect 41580 65326 41582 65378
rect 41634 65326 41860 65378
rect 41580 65324 41860 65326
rect 41580 65314 41636 65324
rect 39452 63924 39508 63934
rect 39340 63922 39620 63924
rect 39340 63870 39454 63922
rect 39506 63870 39620 63922
rect 39340 63868 39620 63870
rect 39452 63858 39508 63868
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 37884 62804 37940 62814
rect 37436 62468 37492 62478
rect 32732 61460 32788 61470
rect 32732 61458 32900 61460
rect 32732 61406 32734 61458
rect 32786 61406 32900 61458
rect 32732 61404 32900 61406
rect 32732 61394 32788 61404
rect 32396 61348 32452 61358
rect 32620 61348 32676 61358
rect 32396 61254 32452 61292
rect 32508 61346 32676 61348
rect 32508 61294 32622 61346
rect 32674 61294 32676 61346
rect 32508 61292 32676 61294
rect 32284 60958 32286 61010
rect 32338 60958 32340 61010
rect 31948 60786 32004 60798
rect 31948 60734 31950 60786
rect 32002 60734 32004 60786
rect 31276 60676 31332 60686
rect 31052 59714 31108 59724
rect 31164 60004 31220 60014
rect 30940 59108 30996 59118
rect 31164 59108 31220 59948
rect 30716 59106 31220 59108
rect 30716 59054 30942 59106
rect 30994 59054 31220 59106
rect 30716 59052 31220 59054
rect 29820 58324 29876 58334
rect 29820 58230 29876 58268
rect 30492 58324 30548 58334
rect 29932 58210 29988 58222
rect 29932 58158 29934 58210
rect 29986 58158 29988 58210
rect 29708 58044 29876 58100
rect 29820 57090 29876 58044
rect 29820 57038 29822 57090
rect 29874 57038 29876 57090
rect 29820 57026 29876 57038
rect 29932 56978 29988 58158
rect 30044 58210 30100 58222
rect 30044 58158 30046 58210
rect 30098 58158 30100 58210
rect 30044 57762 30100 58158
rect 30044 57710 30046 57762
rect 30098 57710 30100 57762
rect 30044 57316 30100 57710
rect 30044 57250 30100 57260
rect 30156 57652 30212 57662
rect 29932 56926 29934 56978
rect 29986 56926 29988 56978
rect 29932 56914 29988 56926
rect 28364 56306 28532 56308
rect 28364 56254 28478 56306
rect 28530 56254 28532 56306
rect 28364 56252 28532 56254
rect 28364 55300 28420 56252
rect 28476 56242 28532 56252
rect 30156 56866 30212 57596
rect 30268 57652 30324 57662
rect 30492 57652 30548 58268
rect 30268 57650 30548 57652
rect 30268 57598 30270 57650
rect 30322 57598 30548 57650
rect 30268 57596 30548 57598
rect 30604 58210 30660 58222
rect 30604 58158 30606 58210
rect 30658 58158 30660 58210
rect 30268 57586 30324 57596
rect 30156 56814 30158 56866
rect 30210 56814 30212 56866
rect 30156 55524 30212 56814
rect 30156 55468 30324 55524
rect 27692 55244 28084 55300
rect 27692 55076 27748 55086
rect 27580 55074 27748 55076
rect 27580 55022 27694 55074
rect 27746 55022 27748 55074
rect 27580 55020 27748 55022
rect 27244 54514 27300 54526
rect 27244 54462 27246 54514
rect 27298 54462 27300 54514
rect 27244 54292 27300 54462
rect 27580 54516 27636 55020
rect 27692 55010 27748 55020
rect 27804 55074 27860 55086
rect 27804 55022 27806 55074
rect 27858 55022 27860 55074
rect 27580 54422 27636 54460
rect 27804 54292 27860 55022
rect 27916 55076 27972 55086
rect 27916 54982 27972 55020
rect 27244 54236 27860 54292
rect 28028 51268 28084 55244
rect 28252 55298 28420 55300
rect 28252 55246 28366 55298
rect 28418 55246 28420 55298
rect 28252 55244 28420 55246
rect 28140 54514 28196 54526
rect 28140 54462 28142 54514
rect 28194 54462 28196 54514
rect 28140 53844 28196 54462
rect 28140 53750 28196 53788
rect 28252 53620 28308 55244
rect 28364 55234 28420 55244
rect 29260 55298 29316 55310
rect 30156 55300 30212 55310
rect 29260 55246 29262 55298
rect 29314 55246 29316 55298
rect 28476 54404 28532 54414
rect 28476 54310 28532 54348
rect 28924 54402 28980 54414
rect 28924 54350 28926 54402
rect 28978 54350 28980 54402
rect 28924 53844 28980 54350
rect 29148 54404 29204 54414
rect 29260 54404 29316 55246
rect 29484 55298 30212 55300
rect 29484 55246 30158 55298
rect 30210 55246 30212 55298
rect 29484 55244 30212 55246
rect 29372 55186 29428 55198
rect 29372 55134 29374 55186
rect 29426 55134 29428 55186
rect 29372 55076 29428 55134
rect 29372 54516 29428 55020
rect 29484 54738 29540 55244
rect 30156 55234 30212 55244
rect 30156 55076 30212 55086
rect 30268 55076 30324 55468
rect 30380 55188 30436 57596
rect 30604 57316 30660 58158
rect 30604 57250 30660 57260
rect 30828 58210 30884 58222
rect 30828 58158 30830 58210
rect 30882 58158 30884 58210
rect 30828 56866 30884 58158
rect 30940 57876 30996 59052
rect 30940 57820 31220 57876
rect 30940 57652 30996 57662
rect 30940 57558 30996 57596
rect 30828 56814 30830 56866
rect 30882 56814 30884 56866
rect 30828 56802 30884 56814
rect 30940 55858 30996 55870
rect 30940 55806 30942 55858
rect 30994 55806 30996 55858
rect 30940 55298 30996 55806
rect 30940 55246 30942 55298
rect 30994 55246 30996 55298
rect 30716 55188 30772 55198
rect 30380 55186 30772 55188
rect 30380 55134 30718 55186
rect 30770 55134 30772 55186
rect 30380 55132 30772 55134
rect 30156 55074 30324 55076
rect 30156 55022 30158 55074
rect 30210 55022 30324 55074
rect 30156 55020 30324 55022
rect 30716 55076 30772 55132
rect 30828 55076 30884 55086
rect 30716 55020 30828 55076
rect 30156 55010 30212 55020
rect 30828 55010 30884 55020
rect 29484 54686 29486 54738
rect 29538 54686 29540 54738
rect 29484 54674 29540 54686
rect 30380 54740 30436 54750
rect 29372 54460 29876 54516
rect 29260 54348 29764 54404
rect 29148 54068 29204 54348
rect 29148 54012 29428 54068
rect 29372 53956 29428 54012
rect 29372 53862 29428 53900
rect 29708 53954 29764 54348
rect 29708 53902 29710 53954
rect 29762 53902 29764 53954
rect 29708 53890 29764 53902
rect 29148 53844 29204 53854
rect 28980 53842 29204 53844
rect 28980 53790 29150 53842
rect 29202 53790 29204 53842
rect 28980 53788 29204 53790
rect 28924 53750 28980 53788
rect 29148 53778 29204 53788
rect 28028 51202 28084 51212
rect 28140 53564 28308 53620
rect 27132 49644 27636 49700
rect 27356 49476 27412 49486
rect 27356 48466 27412 49420
rect 27356 48414 27358 48466
rect 27410 48414 27412 48466
rect 27356 48402 27412 48414
rect 26124 48244 26180 48254
rect 27244 48244 27300 48254
rect 27468 48244 27524 48254
rect 26124 47346 26180 48188
rect 27132 48242 27300 48244
rect 27132 48190 27246 48242
rect 27298 48190 27300 48242
rect 27132 48188 27300 48190
rect 27132 47348 27188 48188
rect 27244 48178 27300 48188
rect 27356 48188 27468 48244
rect 26124 47294 26126 47346
rect 26178 47294 26180 47346
rect 26124 47282 26180 47294
rect 26796 47292 27188 47348
rect 25900 47068 26404 47124
rect 26012 46676 26068 46686
rect 25788 46674 26068 46676
rect 25788 46622 26014 46674
rect 26066 46622 26068 46674
rect 25788 46620 26068 46622
rect 26012 46564 26068 46620
rect 26012 46498 26068 46508
rect 26236 46562 26292 46574
rect 26236 46510 26238 46562
rect 26290 46510 26292 46562
rect 26236 46116 26292 46510
rect 26236 46050 26292 46060
rect 25900 45106 25956 45118
rect 25900 45054 25902 45106
rect 25954 45054 25956 45106
rect 25900 44210 25956 45054
rect 26236 45108 26292 45118
rect 26236 45014 26292 45052
rect 25900 44158 25902 44210
rect 25954 44158 25956 44210
rect 25900 43764 25956 44158
rect 25900 43698 25956 43708
rect 26012 42756 26068 42766
rect 26012 42662 26068 42700
rect 26236 42754 26292 42766
rect 26236 42702 26238 42754
rect 26290 42702 26292 42754
rect 25900 41972 25956 41982
rect 26236 41972 26292 42702
rect 25900 41970 26292 41972
rect 25900 41918 25902 41970
rect 25954 41918 26292 41970
rect 25900 41916 26292 41918
rect 25676 41694 25678 41746
rect 25730 41694 25732 41746
rect 25676 41682 25732 41694
rect 25788 41858 25844 41870
rect 25788 41806 25790 41858
rect 25842 41806 25844 41858
rect 25004 41580 25172 41636
rect 25116 41412 25172 41580
rect 24780 41234 24836 41244
rect 24892 41298 24948 41310
rect 24892 41246 24894 41298
rect 24946 41246 24948 41298
rect 24332 41188 24388 41198
rect 24332 40626 24388 41132
rect 24892 41188 24948 41246
rect 24892 41122 24948 41132
rect 25116 41186 25172 41356
rect 25116 41134 25118 41186
rect 25170 41134 25172 41186
rect 25116 41122 25172 41134
rect 25564 41300 25620 41310
rect 25564 41186 25620 41244
rect 25564 41134 25566 41186
rect 25618 41134 25620 41186
rect 25564 41122 25620 41134
rect 24332 40574 24334 40626
rect 24386 40574 24388 40626
rect 24332 40562 24388 40574
rect 24444 40852 24500 40862
rect 24108 40516 24164 40526
rect 24164 40460 24276 40516
rect 24108 40422 24164 40460
rect 23996 40404 24052 40414
rect 23884 40348 23996 40404
rect 23772 40310 23828 40348
rect 23772 39732 23828 39742
rect 23660 39730 23828 39732
rect 23660 39678 23774 39730
rect 23826 39678 23828 39730
rect 23660 39676 23828 39678
rect 22652 39638 22708 39676
rect 23436 38834 23492 39676
rect 23436 38782 23438 38834
rect 23490 38782 23492 38834
rect 23436 38770 23492 38782
rect 23660 38948 23716 38958
rect 23660 38834 23716 38892
rect 23660 38782 23662 38834
rect 23714 38782 23716 38834
rect 23660 38770 23716 38782
rect 22652 38722 22708 38734
rect 22652 38670 22654 38722
rect 22706 38670 22708 38722
rect 22652 38668 22708 38670
rect 23772 38668 23828 39676
rect 23996 39394 24052 40348
rect 24220 39844 24276 40460
rect 24444 40290 24500 40796
rect 24444 40238 24446 40290
rect 24498 40238 24500 40290
rect 24444 40226 24500 40238
rect 24220 39788 24388 39844
rect 23996 39342 23998 39394
rect 24050 39342 24052 39394
rect 23996 39330 24052 39342
rect 24220 39396 24276 39406
rect 24108 38834 24164 38846
rect 24108 38782 24110 38834
rect 24162 38782 24164 38834
rect 22652 38612 22932 38668
rect 22652 38276 22708 38286
rect 22708 38220 22820 38276
rect 22652 38210 22708 38220
rect 22764 37938 22820 38220
rect 22876 38052 22932 38612
rect 23212 38612 23268 38622
rect 22988 38052 23044 38062
rect 22876 38050 23044 38052
rect 22876 37998 22990 38050
rect 23042 37998 23044 38050
rect 22876 37996 23044 37998
rect 22764 37886 22766 37938
rect 22818 37886 22820 37938
rect 22764 37874 22820 37886
rect 22876 37156 22932 37194
rect 22876 37090 22932 37100
rect 22876 36932 22932 36942
rect 22540 36594 22708 36596
rect 22540 36542 22542 36594
rect 22594 36542 22708 36594
rect 22540 36540 22708 36542
rect 22540 36530 22596 36540
rect 21644 36258 21700 36270
rect 21644 36206 21646 36258
rect 21698 36206 21700 36258
rect 21644 35700 21700 36206
rect 21644 35634 21700 35644
rect 22540 35700 22596 35710
rect 21644 35476 21700 35486
rect 21532 35420 21644 35476
rect 21644 35382 21700 35420
rect 22092 34804 22148 34814
rect 21420 34066 21476 34076
rect 21868 34802 22148 34804
rect 21868 34750 22094 34802
rect 22146 34750 22148 34802
rect 21868 34748 22148 34750
rect 21308 34020 21364 34030
rect 20636 33348 20692 33358
rect 21308 33348 21364 33964
rect 20636 33346 21364 33348
rect 20636 33294 20638 33346
rect 20690 33294 21364 33346
rect 20636 33292 21364 33294
rect 21420 33346 21476 33358
rect 21420 33294 21422 33346
rect 21474 33294 21476 33346
rect 20636 32228 20692 33292
rect 21420 33124 21476 33294
rect 21420 33058 21476 33068
rect 20636 32162 20692 32172
rect 21084 32450 21140 32462
rect 21084 32398 21086 32450
rect 21138 32398 21140 32450
rect 20412 29652 20468 29662
rect 20524 29652 20580 30156
rect 21084 32004 21140 32398
rect 20412 29650 20580 29652
rect 20412 29598 20414 29650
rect 20466 29598 20580 29650
rect 20412 29596 20580 29598
rect 20972 30100 21028 30110
rect 20412 29586 20468 29596
rect 20972 29428 21028 30044
rect 21084 29876 21140 31948
rect 21532 30996 21588 31006
rect 21420 30994 21588 30996
rect 21420 30942 21534 30994
rect 21586 30942 21588 30994
rect 21420 30940 21588 30942
rect 21196 30884 21252 30894
rect 21196 30790 21252 30828
rect 21420 30100 21476 30940
rect 21532 30930 21588 30940
rect 21532 30324 21588 30334
rect 21868 30324 21924 34748
rect 22092 34738 22148 34748
rect 22540 33460 22596 35644
rect 22540 33394 22596 33404
rect 22092 33236 22148 33246
rect 22092 33142 22148 33180
rect 21980 31220 22036 31230
rect 21980 31106 22036 31164
rect 22540 31220 22596 31230
rect 22540 31126 22596 31164
rect 21980 31054 21982 31106
rect 22034 31054 22036 31106
rect 21980 31042 22036 31054
rect 22092 31108 22148 31118
rect 22092 31014 22148 31052
rect 22316 30994 22372 31006
rect 22316 30942 22318 30994
rect 22370 30942 22372 30994
rect 22092 30882 22148 30894
rect 22092 30830 22094 30882
rect 22146 30830 22148 30882
rect 22092 30772 22148 30830
rect 22092 30706 22148 30716
rect 22204 30436 22260 30446
rect 21532 30322 21924 30324
rect 21532 30270 21534 30322
rect 21586 30270 21924 30322
rect 21532 30268 21924 30270
rect 21980 30380 22204 30436
rect 21532 30258 21588 30268
rect 21532 30100 21588 30110
rect 21756 30100 21812 30110
rect 21420 30044 21532 30100
rect 21588 30098 21812 30100
rect 21588 30046 21758 30098
rect 21810 30046 21812 30098
rect 21588 30044 21812 30046
rect 21532 30034 21588 30044
rect 21756 30034 21812 30044
rect 21868 30100 21924 30110
rect 21084 29820 21812 29876
rect 21532 29540 21588 29550
rect 21532 29446 21588 29484
rect 21644 29538 21700 29550
rect 21644 29486 21646 29538
rect 21698 29486 21700 29538
rect 21084 29428 21140 29438
rect 20972 29426 21140 29428
rect 20972 29374 21086 29426
rect 21138 29374 21140 29426
rect 20972 29372 21140 29374
rect 21084 29204 21140 29372
rect 21532 29316 21588 29326
rect 21084 29138 21140 29148
rect 21196 29314 21588 29316
rect 21196 29262 21534 29314
rect 21586 29262 21588 29314
rect 21196 29260 21588 29262
rect 21196 28644 21252 29260
rect 21532 29250 21588 29260
rect 21644 28980 21700 29486
rect 20300 28588 21252 28644
rect 21308 28924 21644 28980
rect 20300 27970 20356 28588
rect 21308 28532 21364 28924
rect 21644 28914 21700 28924
rect 20300 27918 20302 27970
rect 20354 27918 20356 27970
rect 20300 27906 20356 27918
rect 20748 28476 21364 28532
rect 20748 28418 20804 28476
rect 20748 28366 20750 28418
rect 20802 28366 20804 28418
rect 20748 26908 20804 28366
rect 21756 26908 21812 29820
rect 21868 29650 21924 30044
rect 21980 30098 22036 30380
rect 22204 30370 22260 30380
rect 22316 30210 22372 30942
rect 22316 30158 22318 30210
rect 22370 30158 22372 30210
rect 21980 30046 21982 30098
rect 22034 30046 22036 30098
rect 21980 30034 22036 30046
rect 22092 30098 22148 30110
rect 22092 30046 22094 30098
rect 22146 30046 22148 30098
rect 22092 29988 22148 30046
rect 22316 30100 22372 30158
rect 22316 30034 22372 30044
rect 22204 29988 22260 29998
rect 22092 29932 22204 29988
rect 22204 29922 22260 29932
rect 22652 29764 22708 36540
rect 22764 36484 22820 36494
rect 22764 36390 22820 36428
rect 22876 35586 22932 36876
rect 22988 35700 23044 37996
rect 23100 37940 23156 37950
rect 23100 36706 23156 37884
rect 23100 36654 23102 36706
rect 23154 36654 23156 36706
rect 23100 36642 23156 36654
rect 22988 35634 23044 35644
rect 22876 35534 22878 35586
rect 22930 35534 22932 35586
rect 22876 35522 22932 35534
rect 22764 33572 22820 33582
rect 22764 31218 22820 33516
rect 22764 31166 22766 31218
rect 22818 31166 22820 31218
rect 22764 31154 22820 31166
rect 22876 30996 22932 31006
rect 22876 30902 22932 30940
rect 23100 30994 23156 31006
rect 23100 30942 23102 30994
rect 23154 30942 23156 30994
rect 23100 30436 23156 30942
rect 23212 30996 23268 38556
rect 23548 38612 23828 38668
rect 23884 38724 23940 38762
rect 23884 38658 23940 38668
rect 23996 38612 24052 38622
rect 23324 36484 23380 36494
rect 23324 35922 23380 36428
rect 23324 35870 23326 35922
rect 23378 35870 23380 35922
rect 23324 35858 23380 35870
rect 23324 35364 23380 35374
rect 23324 31218 23380 35308
rect 23548 34018 23604 38612
rect 23996 37940 24052 38556
rect 24108 38052 24164 38782
rect 24220 38612 24276 39340
rect 24220 38518 24276 38556
rect 24108 37986 24164 37996
rect 24220 38050 24276 38062
rect 24220 37998 24222 38050
rect 24274 37998 24276 38050
rect 23996 37846 24052 37884
rect 24220 37940 24276 37998
rect 24220 37874 24276 37884
rect 24332 37716 24388 39788
rect 25004 39732 25060 39742
rect 25788 39732 25844 41806
rect 25900 41186 25956 41916
rect 25900 41134 25902 41186
rect 25954 41134 25956 41186
rect 25900 41122 25956 41134
rect 26012 41188 26068 41198
rect 26012 39842 26068 41132
rect 26012 39790 26014 39842
rect 26066 39790 26068 39842
rect 26012 39778 26068 39790
rect 25004 39506 25060 39676
rect 25676 39676 25844 39732
rect 26124 39732 26180 39742
rect 25004 39454 25006 39506
rect 25058 39454 25060 39506
rect 25004 39442 25060 39454
rect 25564 39620 25620 39630
rect 24780 39172 24836 39182
rect 23996 37660 24388 37716
rect 24444 38948 24500 38958
rect 23660 37378 23716 37390
rect 23660 37326 23662 37378
rect 23714 37326 23716 37378
rect 23660 36932 23716 37326
rect 23996 37268 24052 37660
rect 23996 37212 24164 37268
rect 23660 36482 23716 36876
rect 23660 36430 23662 36482
rect 23714 36430 23716 36482
rect 23660 36418 23716 36430
rect 23884 37156 23940 37166
rect 23884 34132 23940 37100
rect 24108 36594 24164 37212
rect 24108 36542 24110 36594
rect 24162 36542 24164 36594
rect 24108 36530 24164 36542
rect 23996 36482 24052 36494
rect 23996 36430 23998 36482
rect 24050 36430 24052 36482
rect 23996 35698 24052 36430
rect 24332 36482 24388 36494
rect 24332 36430 24334 36482
rect 24386 36430 24388 36482
rect 24332 36372 24388 36430
rect 24220 35924 24276 35934
rect 24220 35830 24276 35868
rect 23996 35646 23998 35698
rect 24050 35646 24052 35698
rect 23996 35028 24052 35646
rect 24220 35028 24276 35038
rect 23996 35026 24276 35028
rect 23996 34974 24222 35026
rect 24274 34974 24276 35026
rect 23996 34972 24276 34974
rect 24220 34962 24276 34972
rect 23884 34130 24276 34132
rect 23884 34078 23886 34130
rect 23938 34078 24276 34130
rect 23884 34076 24276 34078
rect 23884 34066 23940 34076
rect 23548 33966 23550 34018
rect 23602 33966 23604 34018
rect 23548 33572 23604 33966
rect 23548 33506 23604 33516
rect 24220 33458 24276 34076
rect 24220 33406 24222 33458
rect 24274 33406 24276 33458
rect 24220 33394 24276 33406
rect 24332 33236 24388 36316
rect 24108 33180 24388 33236
rect 24444 36484 24500 38892
rect 24556 38836 24612 38846
rect 24556 38274 24612 38780
rect 24556 38222 24558 38274
rect 24610 38222 24612 38274
rect 24556 38210 24612 38222
rect 24556 37940 24612 37950
rect 24780 37940 24836 39116
rect 25564 38722 25620 39564
rect 25676 38836 25732 39676
rect 26124 39638 26180 39676
rect 26236 39618 26292 39630
rect 26236 39566 26238 39618
rect 26290 39566 26292 39618
rect 26236 38948 26292 39566
rect 26236 38882 26292 38892
rect 25676 38742 25732 38780
rect 26012 38836 26068 38846
rect 25564 38670 25566 38722
rect 25618 38670 25620 38722
rect 25564 38668 25620 38670
rect 25564 38612 25732 38668
rect 24612 37884 24836 37940
rect 24892 38164 24948 38174
rect 24556 37490 24612 37884
rect 24556 37438 24558 37490
rect 24610 37438 24612 37490
rect 24556 37426 24612 37438
rect 24556 37268 24612 37278
rect 24556 36706 24612 37212
rect 24892 37268 24948 38108
rect 25340 38052 25396 38062
rect 25340 37492 25396 37996
rect 25340 37398 25396 37436
rect 24892 37202 24948 37212
rect 25228 37156 25284 37166
rect 25228 37062 25284 37100
rect 24556 36654 24558 36706
rect 24610 36654 24612 36706
rect 24556 36642 24612 36654
rect 24668 36484 24724 36494
rect 24444 36482 24724 36484
rect 24444 36430 24670 36482
rect 24722 36430 24724 36482
rect 24444 36428 24724 36430
rect 23324 31166 23326 31218
rect 23378 31166 23380 31218
rect 23324 31154 23380 31166
rect 23884 33124 23940 33134
rect 23884 31778 23940 33068
rect 24108 32786 24164 33180
rect 24444 32788 24500 36428
rect 24668 36418 24724 36428
rect 25340 35924 25396 35934
rect 25340 35698 25396 35868
rect 25340 35646 25342 35698
rect 25394 35646 25396 35698
rect 25340 35634 25396 35646
rect 25452 35588 25508 35598
rect 25452 34018 25508 35532
rect 25676 35586 25732 38612
rect 26012 38274 26068 38780
rect 26012 38222 26014 38274
rect 26066 38222 26068 38274
rect 26012 38210 26068 38222
rect 26124 38612 26180 38622
rect 26124 38050 26180 38556
rect 26124 37998 26126 38050
rect 26178 37998 26180 38050
rect 26124 37986 26180 37998
rect 26012 37828 26068 37838
rect 26012 37378 26068 37772
rect 26012 37326 26014 37378
rect 26066 37326 26068 37378
rect 26012 35924 26068 37326
rect 26124 37380 26180 37390
rect 26124 37286 26180 37324
rect 26012 35858 26068 35868
rect 25676 35534 25678 35586
rect 25730 35534 25732 35586
rect 25676 35364 25732 35534
rect 25676 35298 25732 35308
rect 25452 33966 25454 34018
rect 25506 33966 25508 34018
rect 25452 33954 25508 33966
rect 25116 33460 25172 33470
rect 24668 33124 24724 33134
rect 24668 33030 24724 33068
rect 25116 33124 25172 33404
rect 25788 33236 25844 33246
rect 25788 33142 25844 33180
rect 25452 33124 25508 33134
rect 25116 33122 25508 33124
rect 25116 33070 25118 33122
rect 25170 33070 25454 33122
rect 25506 33070 25508 33122
rect 25116 33068 25508 33070
rect 24108 32734 24110 32786
rect 24162 32734 24164 32786
rect 24108 31892 24164 32734
rect 24108 31826 24164 31836
rect 24220 32786 24500 32788
rect 24220 32734 24446 32786
rect 24498 32734 24500 32786
rect 24220 32732 24500 32734
rect 23884 31726 23886 31778
rect 23938 31726 23940 31778
rect 23436 30996 23492 31006
rect 23212 30940 23380 30996
rect 23100 30370 23156 30380
rect 22876 29988 22932 29998
rect 22932 29932 23044 29988
rect 22876 29894 22932 29932
rect 21868 29598 21870 29650
rect 21922 29598 21924 29650
rect 21868 29586 21924 29598
rect 22316 29708 22708 29764
rect 22316 29650 22372 29708
rect 22316 29598 22318 29650
rect 22370 29598 22372 29650
rect 22092 29540 22148 29550
rect 22092 29446 22148 29484
rect 22316 27748 22372 29598
rect 22428 29540 22484 29550
rect 22428 29446 22484 29484
rect 22876 29538 22932 29550
rect 22876 29486 22878 29538
rect 22930 29486 22932 29538
rect 22876 29204 22932 29486
rect 22876 29138 22932 29148
rect 22876 27860 22932 27870
rect 22428 27748 22484 27758
rect 22316 27746 22484 27748
rect 22316 27694 22430 27746
rect 22482 27694 22484 27746
rect 22316 27692 22484 27694
rect 22428 27682 22484 27692
rect 20188 26852 20356 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19964 25620 20020 25630
rect 19964 25526 20020 25564
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19740 24724 19796 24734
rect 19628 24722 19796 24724
rect 19628 24670 19742 24722
rect 19794 24670 19796 24722
rect 19628 24668 19796 24670
rect 19740 24658 19796 24668
rect 18620 24610 18676 24622
rect 18620 24558 18622 24610
rect 18674 24558 18676 24610
rect 18620 24388 18676 24558
rect 18620 24322 18676 24332
rect 16660 23660 16772 23716
rect 16604 23622 16660 23660
rect 15932 23214 15934 23266
rect 15986 23214 15988 23266
rect 15932 23202 15988 23214
rect 13804 22990 13806 23042
rect 13858 22990 13860 23042
rect 13804 22978 13860 22990
rect 16716 23154 16772 23660
rect 18284 23650 18340 23660
rect 18844 24052 18900 24062
rect 16716 23102 16718 23154
rect 16770 23102 16772 23154
rect 16716 23044 16772 23102
rect 16716 22978 16772 22988
rect 17500 23044 17556 23054
rect 15260 20802 15316 20814
rect 15260 20750 15262 20802
rect 15314 20750 15316 20802
rect 14812 20578 14868 20590
rect 14812 20526 14814 20578
rect 14866 20526 14868 20578
rect 14812 20244 14868 20526
rect 14364 20132 14868 20188
rect 15260 20244 15316 20750
rect 15932 20692 15988 20702
rect 15932 20598 15988 20636
rect 15260 20178 15316 20188
rect 14364 19234 14420 20132
rect 17500 20020 17556 22988
rect 18620 21812 18676 21822
rect 18620 21718 18676 21756
rect 18284 21698 18340 21710
rect 18284 21646 18286 21698
rect 18338 21646 18340 21698
rect 18060 20916 18116 20926
rect 18060 20914 18228 20916
rect 18060 20862 18062 20914
rect 18114 20862 18228 20914
rect 18060 20860 18228 20862
rect 18060 20850 18116 20860
rect 18172 20132 18228 20860
rect 18172 20066 18228 20076
rect 18284 20802 18340 21646
rect 18844 21028 18900 23996
rect 19404 24052 19460 24062
rect 19404 23958 19460 23996
rect 18956 23940 19012 23950
rect 18956 23380 19012 23884
rect 19852 23938 19908 23950
rect 19852 23886 19854 23938
rect 19906 23886 19908 23938
rect 19852 23716 19908 23886
rect 19852 23650 19908 23660
rect 20300 23938 20356 26852
rect 20412 26852 20804 26908
rect 21644 26852 21812 26908
rect 22876 26964 22932 27804
rect 22876 26898 22932 26908
rect 20412 24052 20468 26852
rect 21420 25394 21476 25406
rect 21420 25342 21422 25394
rect 21474 25342 21476 25394
rect 21420 25172 21476 25342
rect 21420 25106 21476 25116
rect 21532 25282 21588 25294
rect 21532 25230 21534 25282
rect 21586 25230 21588 25282
rect 21532 24948 21588 25230
rect 20524 24892 21588 24948
rect 20524 24834 20580 24892
rect 20524 24782 20526 24834
rect 20578 24782 20580 24834
rect 20524 24770 20580 24782
rect 20412 23986 20468 23996
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18956 23314 19012 23324
rect 19628 23380 19684 23390
rect 19628 23286 19684 23324
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19292 21812 19348 21822
rect 19292 21718 19348 21756
rect 19964 21812 20020 21822
rect 19964 21718 20020 21756
rect 18956 21700 19012 21710
rect 19012 21644 19236 21700
rect 18956 21606 19012 21644
rect 18844 20972 19124 21028
rect 18284 20750 18286 20802
rect 18338 20750 18340 20802
rect 18060 20020 18116 20030
rect 17500 19964 18060 20020
rect 14364 19182 14366 19234
rect 14418 19182 14420 19234
rect 14364 19170 14420 19182
rect 17164 19346 17220 19358
rect 17164 19294 17166 19346
rect 17218 19294 17220 19346
rect 15036 19122 15092 19134
rect 15036 19070 15038 19122
rect 15090 19070 15092 19122
rect 15036 18452 15092 19070
rect 17164 19012 17220 19294
rect 17724 19346 17780 19964
rect 18060 19926 18116 19964
rect 18284 19908 18340 20750
rect 18732 20916 18788 20926
rect 18732 20802 18788 20860
rect 18732 20750 18734 20802
rect 18786 20750 18788 20802
rect 18732 20738 18788 20750
rect 18844 20802 18900 20814
rect 18844 20750 18846 20802
rect 18898 20750 18900 20802
rect 18508 20692 18564 20702
rect 18508 20598 18564 20636
rect 17724 19294 17726 19346
rect 17778 19294 17780 19346
rect 17724 19282 17780 19294
rect 18172 19852 18340 19908
rect 18396 20580 18452 20590
rect 18396 20130 18452 20524
rect 18844 20356 18900 20750
rect 18508 20300 18900 20356
rect 18508 20242 18564 20300
rect 18508 20190 18510 20242
rect 18562 20190 18564 20242
rect 18508 20178 18564 20190
rect 18396 20078 18398 20130
rect 18450 20078 18452 20130
rect 18172 19124 18228 19852
rect 18284 19236 18340 19246
rect 18396 19236 18452 20078
rect 18620 20132 18676 20142
rect 18620 20020 18676 20076
rect 18620 20018 18900 20020
rect 18620 19966 18622 20018
rect 18674 19966 18900 20018
rect 18620 19964 18900 19966
rect 18620 19954 18676 19964
rect 18284 19234 18452 19236
rect 18284 19182 18286 19234
rect 18338 19182 18452 19234
rect 18284 19180 18452 19182
rect 18284 19170 18340 19180
rect 17948 19068 18228 19124
rect 17164 18946 17220 18956
rect 17836 19012 17892 19022
rect 15036 18386 15092 18396
rect 17388 18340 17444 18350
rect 17388 17666 17444 18284
rect 17388 17614 17390 17666
rect 17442 17614 17444 17666
rect 14700 17444 14756 17454
rect 14700 16994 14756 17388
rect 17388 17332 17444 17614
rect 17724 17554 17780 17566
rect 17724 17502 17726 17554
rect 17778 17502 17780 17554
rect 17500 17444 17556 17454
rect 17500 17350 17556 17388
rect 17388 17266 17444 17276
rect 17724 17220 17780 17502
rect 17836 17444 17892 18956
rect 17948 18450 18004 19068
rect 18396 19010 18452 19022
rect 18396 18958 18398 19010
rect 18450 18958 18452 19010
rect 18396 18788 18452 18958
rect 18508 19012 18564 19022
rect 18508 18918 18564 18956
rect 18396 18732 18564 18788
rect 18508 18562 18564 18732
rect 18508 18510 18510 18562
rect 18562 18510 18564 18562
rect 18508 18498 18564 18510
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18340 18004 18398
rect 18060 18452 18116 18462
rect 18060 18358 18116 18396
rect 18284 18452 18340 18462
rect 18284 18358 18340 18396
rect 17948 18274 18004 18284
rect 17948 17668 18004 17678
rect 18396 17668 18452 17678
rect 17948 17666 18452 17668
rect 17948 17614 17950 17666
rect 18002 17614 18398 17666
rect 18450 17614 18452 17666
rect 17948 17612 18452 17614
rect 17948 17602 18004 17612
rect 18396 17602 18452 17612
rect 18284 17444 18340 17482
rect 17836 17388 18228 17444
rect 17724 17154 17780 17164
rect 16828 17108 16884 17118
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 16716 16996 16772 17006
rect 12908 16258 12964 16268
rect 14028 16882 14084 16894
rect 14028 16830 14030 16882
rect 14082 16830 14084 16882
rect 14028 16212 14084 16830
rect 14028 13746 14084 16156
rect 15932 16772 15988 16782
rect 15932 16212 15988 16716
rect 15932 16098 15988 16156
rect 16716 16210 16772 16940
rect 16828 16770 16884 17052
rect 18060 17108 18116 17118
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 17612 16884 17668 16894
rect 16716 16158 16718 16210
rect 16770 16158 16772 16210
rect 16716 16146 16772 16158
rect 15932 16046 15934 16098
rect 15986 16046 15988 16098
rect 15932 16034 15988 16046
rect 17612 15148 17668 16828
rect 17500 15092 17668 15148
rect 14700 13972 14756 13982
rect 14700 13858 14756 13916
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 17500 13970 17556 15092
rect 17500 13918 17502 13970
rect 17554 13918 17556 13970
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13682 14084 13694
rect 16828 13636 16884 13646
rect 16828 13542 16884 13580
rect 17500 13524 17556 13918
rect 17500 13458 17556 13468
rect 17836 13188 17892 13198
rect 17836 13094 17892 13132
rect 17948 12964 18004 12974
rect 17948 12870 18004 12908
rect 17836 12740 17892 12750
rect 5852 11666 5908 11676
rect 14476 11732 14532 11742
rect 14476 11394 14532 11676
rect 17724 11732 17780 11742
rect 17276 11508 17332 11518
rect 17724 11508 17780 11676
rect 17276 11414 17332 11452
rect 17500 11506 17780 11508
rect 17500 11454 17726 11506
rect 17778 11454 17780 11506
rect 17500 11452 17780 11454
rect 14476 11342 14478 11394
rect 14530 11342 14532 11394
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 14476 9826 14532 11342
rect 15148 11284 15204 11294
rect 15148 11282 15764 11284
rect 15148 11230 15150 11282
rect 15202 11230 15764 11282
rect 15148 11228 15764 11230
rect 15148 11218 15204 11228
rect 15708 10834 15764 11228
rect 15708 10782 15710 10834
rect 15762 10782 15764 10834
rect 15708 10770 15764 10782
rect 15820 11172 15876 11182
rect 15820 10722 15876 11116
rect 15820 10670 15822 10722
rect 15874 10670 15876 10722
rect 15820 10658 15876 10670
rect 14476 9774 14478 9826
rect 14530 9774 14532 9826
rect 14476 9762 14532 9774
rect 17276 9938 17332 9950
rect 17276 9886 17278 9938
rect 17330 9886 17332 9938
rect 17276 9828 17332 9886
rect 17276 9762 17332 9772
rect 15148 9716 15204 9726
rect 15148 9714 15764 9716
rect 15148 9662 15150 9714
rect 15202 9662 15764 9714
rect 15148 9660 15764 9662
rect 15148 9650 15204 9660
rect 15708 9266 15764 9660
rect 15708 9214 15710 9266
rect 15762 9214 15764 9266
rect 15708 9202 15764 9214
rect 15820 9604 15876 9614
rect 15820 9154 15876 9548
rect 15820 9102 15822 9154
rect 15874 9102 15876 9154
rect 15820 9090 15876 9102
rect 17500 9266 17556 11452
rect 17724 11442 17780 11452
rect 17724 10052 17780 10062
rect 17836 10052 17892 12684
rect 18060 10722 18116 17052
rect 18172 15148 18228 17388
rect 18284 17378 18340 17388
rect 18508 17442 18564 17454
rect 18508 17390 18510 17442
rect 18562 17390 18564 17442
rect 18396 17332 18452 17342
rect 18284 17220 18340 17230
rect 18284 17106 18340 17164
rect 18284 17054 18286 17106
rect 18338 17054 18340 17106
rect 18284 17042 18340 17054
rect 18396 16882 18452 17276
rect 18508 17108 18564 17390
rect 18508 17042 18564 17052
rect 18732 17108 18788 17118
rect 18732 17014 18788 17052
rect 18732 16884 18788 16894
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 18396 16818 18452 16830
rect 18508 16882 18788 16884
rect 18508 16830 18734 16882
rect 18786 16830 18788 16882
rect 18508 16828 18788 16830
rect 18508 15988 18564 16828
rect 18732 16818 18788 16828
rect 18844 16548 18900 19964
rect 18956 20018 19012 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18956 19234 19012 19966
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 18956 17668 19012 19182
rect 19068 19348 19124 20972
rect 19068 18452 19124 19292
rect 19068 18358 19124 18396
rect 18956 17574 19012 17612
rect 19180 17666 19236 21644
rect 19628 21698 19684 21710
rect 19628 21646 19630 21698
rect 19682 21646 19684 21698
rect 19404 20916 19460 20926
rect 19404 20822 19460 20860
rect 19628 20580 19684 21646
rect 20076 21700 20132 21710
rect 20076 20802 20132 21644
rect 20300 20916 20356 23886
rect 20748 23716 20804 23726
rect 20748 23268 20804 23660
rect 20748 23202 20804 23212
rect 20300 20850 20356 20860
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 20524 20804 20580 20814
rect 20524 20710 20580 20748
rect 20748 20692 20804 20702
rect 20748 20598 20804 20636
rect 19628 20514 19684 20524
rect 20300 20578 20356 20590
rect 20300 20526 20302 20578
rect 20354 20526 20356 20578
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20132 20244 20142
rect 20300 20132 20356 20526
rect 20188 20130 20356 20132
rect 20188 20078 20190 20130
rect 20242 20078 20356 20130
rect 20188 20076 20356 20078
rect 20188 20066 20244 20076
rect 19404 20020 19460 20030
rect 19404 19926 19460 19964
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 19180 17444 19236 17614
rect 19852 18116 19908 18126
rect 19852 17666 19908 18060
rect 21532 17780 21588 17790
rect 21644 17780 21700 26852
rect 22876 26628 22932 26638
rect 22764 26290 22820 26302
rect 22764 26238 22766 26290
rect 22818 26238 22820 26290
rect 22316 26180 22372 26190
rect 22316 26086 22372 26124
rect 22764 26180 22820 26238
rect 22764 26114 22820 26124
rect 21756 25394 21812 25406
rect 21756 25342 21758 25394
rect 21810 25342 21812 25394
rect 21756 25284 21812 25342
rect 21980 25396 22036 25406
rect 21980 25394 22372 25396
rect 21980 25342 21982 25394
rect 22034 25342 22372 25394
rect 21980 25340 22372 25342
rect 21980 25330 22036 25340
rect 21756 25218 21812 25228
rect 22204 25172 22260 25182
rect 22204 23940 22260 25116
rect 22316 24050 22372 25340
rect 22316 23998 22318 24050
rect 22370 23998 22372 24050
rect 22316 23986 22372 23998
rect 22540 25284 22596 25294
rect 21980 23714 22036 23726
rect 21980 23662 21982 23714
rect 22034 23662 22036 23714
rect 21980 23380 22036 23662
rect 21980 23314 22036 23324
rect 22204 23156 22260 23884
rect 22428 23714 22484 23726
rect 22428 23662 22430 23714
rect 22482 23662 22484 23714
rect 22428 23604 22484 23662
rect 22428 23538 22484 23548
rect 22540 23268 22596 25228
rect 22652 24612 22708 24622
rect 22652 24518 22708 24556
rect 22876 23938 22932 26572
rect 22988 24388 23044 29932
rect 23212 29652 23268 29662
rect 23212 29558 23268 29596
rect 23324 26908 23380 30940
rect 23436 29540 23492 30940
rect 23884 30212 23940 31726
rect 24108 31220 24164 31230
rect 24220 31220 24276 32732
rect 24444 32722 24500 32732
rect 24668 31668 24724 31678
rect 24668 31666 25060 31668
rect 24668 31614 24670 31666
rect 24722 31614 25060 31666
rect 24668 31612 25060 31614
rect 24668 31602 24724 31612
rect 24108 31218 24276 31220
rect 24108 31166 24110 31218
rect 24162 31166 24276 31218
rect 24108 31164 24276 31166
rect 24108 31154 24164 31164
rect 23996 30996 24052 31006
rect 23996 30902 24052 30940
rect 24332 30996 24388 31006
rect 24332 30994 24612 30996
rect 24332 30942 24334 30994
rect 24386 30942 24612 30994
rect 24332 30940 24612 30942
rect 24332 30930 24388 30940
rect 23996 30212 24052 30222
rect 23884 30156 23996 30212
rect 23996 30146 24052 30156
rect 24220 30100 24276 30110
rect 24220 29652 24276 30044
rect 24556 30098 24612 30940
rect 25004 30322 25060 31612
rect 25004 30270 25006 30322
rect 25058 30270 25060 30322
rect 25004 30258 25060 30270
rect 24556 30046 24558 30098
rect 24610 30046 24612 30098
rect 24556 30034 24612 30046
rect 24780 30098 24836 30110
rect 24780 30046 24782 30098
rect 24834 30046 24836 30098
rect 24444 29988 24500 29998
rect 24444 29894 24500 29932
rect 24332 29652 24388 29662
rect 24220 29650 24388 29652
rect 24220 29598 24334 29650
rect 24386 29598 24388 29650
rect 24220 29596 24388 29598
rect 24332 29586 24388 29596
rect 23660 29540 23716 29550
rect 23436 29484 23660 29540
rect 23660 29446 23716 29484
rect 23996 29426 24052 29438
rect 23996 29374 23998 29426
rect 24050 29374 24052 29426
rect 23996 29316 24052 29374
rect 24556 29426 24612 29438
rect 24556 29374 24558 29426
rect 24610 29374 24612 29426
rect 24556 29316 24612 29374
rect 24780 29428 24836 30046
rect 24780 29362 24836 29372
rect 23996 29260 24612 29316
rect 24556 27298 24612 29260
rect 24556 27246 24558 27298
rect 24610 27246 24612 27298
rect 24556 27234 24612 27246
rect 23996 26964 24052 26974
rect 23324 26852 23492 26908
rect 23212 26178 23268 26190
rect 23212 26126 23214 26178
rect 23266 26126 23268 26178
rect 23212 25844 23268 26126
rect 23212 25778 23268 25788
rect 23324 26180 23380 26190
rect 23324 25618 23380 26124
rect 23324 25566 23326 25618
rect 23378 25566 23380 25618
rect 23324 25554 23380 25566
rect 23436 24948 23492 26852
rect 23772 26290 23828 26302
rect 23772 26238 23774 26290
rect 23826 26238 23828 26290
rect 23772 26180 23828 26238
rect 23772 26114 23828 26124
rect 23324 24892 23492 24948
rect 22988 24322 23044 24332
rect 23100 24610 23156 24622
rect 23100 24558 23102 24610
rect 23154 24558 23156 24610
rect 22876 23886 22878 23938
rect 22930 23886 22932 23938
rect 22876 23380 22932 23886
rect 23100 23604 23156 24558
rect 23100 23538 23156 23548
rect 22428 23212 22596 23268
rect 22764 23324 22876 23380
rect 22316 23156 22372 23166
rect 22204 23154 22372 23156
rect 22204 23102 22318 23154
rect 22370 23102 22372 23154
rect 22204 23100 22372 23102
rect 22316 23090 22372 23100
rect 22428 22932 22484 23212
rect 22652 23154 22708 23166
rect 22652 23102 22654 23154
rect 22706 23102 22708 23154
rect 22316 22876 22484 22932
rect 22540 23042 22596 23054
rect 22540 22990 22542 23042
rect 22594 22990 22596 23042
rect 21756 21588 21812 21598
rect 21756 21494 21812 21532
rect 21868 20692 21924 20702
rect 21868 20598 21924 20636
rect 21756 20580 21812 20590
rect 21756 18674 21812 20524
rect 21980 20578 22036 20590
rect 21980 20526 21982 20578
rect 22034 20526 22036 20578
rect 21980 19908 22036 20526
rect 22316 20468 22372 22876
rect 22428 21700 22484 21710
rect 22540 21700 22596 22990
rect 22428 21698 22596 21700
rect 22428 21646 22430 21698
rect 22482 21646 22596 21698
rect 22428 21644 22596 21646
rect 22652 22820 22708 23102
rect 22428 21634 22484 21644
rect 22428 20802 22484 20814
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 22428 20580 22484 20750
rect 22652 20804 22708 22764
rect 22652 20738 22708 20748
rect 22764 20914 22820 23324
rect 22876 23314 22932 23324
rect 22988 23156 23044 23166
rect 22988 23062 23044 23100
rect 22764 20862 22766 20914
rect 22818 20862 22820 20914
rect 22764 20580 22820 20862
rect 22428 20524 22820 20580
rect 22316 20412 22484 20468
rect 22316 19908 22372 19918
rect 22036 19906 22372 19908
rect 22036 19854 22318 19906
rect 22370 19854 22372 19906
rect 22036 19852 22372 19854
rect 21980 19842 22036 19852
rect 22316 19842 22372 19852
rect 22428 19684 22484 20412
rect 21756 18622 21758 18674
rect 21810 18622 21812 18674
rect 21756 18610 21812 18622
rect 22316 19628 22484 19684
rect 22876 19908 22932 19918
rect 21980 18452 22036 18462
rect 21980 18450 22260 18452
rect 21980 18398 21982 18450
rect 22034 18398 22260 18450
rect 21980 18396 22260 18398
rect 21980 18386 22036 18396
rect 21868 18338 21924 18350
rect 21868 18286 21870 18338
rect 21922 18286 21924 18338
rect 21644 17724 21812 17780
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17602 19908 17614
rect 21196 17666 21252 17678
rect 21196 17614 21198 17666
rect 21250 17614 21252 17666
rect 19180 17378 19236 17388
rect 19292 17442 19348 17454
rect 19292 17390 19294 17442
rect 19346 17390 19348 17442
rect 19068 16996 19124 17006
rect 19292 16996 19348 17390
rect 19068 16994 19348 16996
rect 19068 16942 19070 16994
rect 19122 16942 19348 16994
rect 19068 16940 19348 16942
rect 19404 17442 19460 17454
rect 19404 17390 19406 17442
rect 19458 17390 19460 17442
rect 19068 16930 19124 16940
rect 18508 15922 18564 15932
rect 18620 16492 18900 16548
rect 18172 15092 18340 15148
rect 18284 14642 18340 15092
rect 18284 14590 18286 14642
rect 18338 14590 18340 14642
rect 18284 14578 18340 14590
rect 18508 14532 18564 14542
rect 18284 13746 18340 13758
rect 18284 13694 18286 13746
rect 18338 13694 18340 13746
rect 18284 13412 18340 13694
rect 18284 13188 18340 13356
rect 18284 13122 18340 13132
rect 18396 12962 18452 12974
rect 18396 12910 18398 12962
rect 18450 12910 18452 12962
rect 18284 12178 18340 12190
rect 18284 12126 18286 12178
rect 18338 12126 18340 12178
rect 18284 12068 18340 12126
rect 18284 12002 18340 12012
rect 18284 11508 18340 11518
rect 18396 11508 18452 12910
rect 18508 12740 18564 14476
rect 18620 12962 18676 16492
rect 19404 16324 19460 17390
rect 21196 17444 21252 17614
rect 21532 17666 21588 17724
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 21532 17602 21588 17614
rect 21196 17378 21252 17388
rect 21420 17442 21476 17454
rect 21420 17390 21422 17442
rect 21474 17390 21476 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 21420 17108 21476 17390
rect 20636 17052 21476 17108
rect 20636 16994 20692 17052
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16930 20692 16942
rect 18844 16268 19460 16324
rect 19628 16884 19684 16894
rect 19852 16884 19908 16894
rect 19684 16882 19908 16884
rect 19684 16830 19854 16882
rect 19906 16830 19908 16882
rect 19684 16828 19908 16830
rect 18844 16210 18900 16268
rect 18844 16158 18846 16210
rect 18898 16158 18900 16210
rect 18844 15148 18900 16158
rect 19628 16212 19684 16828
rect 19852 16818 19908 16828
rect 19740 16212 19796 16222
rect 19628 16210 19796 16212
rect 19628 16158 19742 16210
rect 19794 16158 19796 16210
rect 19628 16156 19796 16158
rect 19740 16146 19796 16156
rect 21756 16212 21812 17724
rect 21868 17666 21924 18286
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21868 17602 21924 17614
rect 22204 16884 22260 18396
rect 22316 17780 22372 19628
rect 22316 17686 22372 17724
rect 22428 18450 22484 18462
rect 22428 18398 22430 18450
rect 22482 18398 22484 18450
rect 22428 17668 22484 18398
rect 22428 17556 22484 17612
rect 22764 17556 22820 17566
rect 22428 17554 22820 17556
rect 22428 17502 22766 17554
rect 22818 17502 22820 17554
rect 22428 17500 22820 17502
rect 22764 17490 22820 17500
rect 22204 16828 22820 16884
rect 22428 16212 22484 16222
rect 21812 16156 21924 16212
rect 21756 16146 21812 16156
rect 19292 15988 19348 15998
rect 19292 15894 19348 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 21868 15538 21924 16156
rect 22428 16118 22484 16156
rect 21868 15486 21870 15538
rect 21922 15486 21924 15538
rect 21868 15474 21924 15486
rect 18732 15092 18900 15148
rect 22428 15202 22484 15214
rect 22428 15150 22430 15202
rect 22482 15150 22484 15202
rect 22428 15148 22484 15150
rect 22652 15148 22708 16828
rect 22764 16770 22820 16828
rect 22764 16718 22766 16770
rect 22818 16718 22820 16770
rect 22764 16706 22820 16718
rect 22764 16212 22820 16222
rect 22764 16098 22820 16156
rect 22764 16046 22766 16098
rect 22818 16046 22820 16098
rect 22764 16034 22820 16046
rect 22876 16100 22932 19852
rect 23212 19236 23268 19246
rect 23212 18676 23268 19180
rect 22988 18620 23268 18676
rect 22988 18450 23044 18620
rect 22988 18398 22990 18450
rect 23042 18398 23044 18450
rect 22988 18386 23044 18398
rect 23100 18452 23156 18462
rect 23100 17666 23156 18396
rect 23212 18450 23268 18620
rect 23212 18398 23214 18450
rect 23266 18398 23268 18450
rect 23212 18386 23268 18398
rect 23100 17614 23102 17666
rect 23154 17614 23156 17666
rect 23100 17602 23156 17614
rect 23324 17444 23380 24892
rect 23436 24722 23492 24734
rect 23436 24670 23438 24722
rect 23490 24670 23492 24722
rect 23436 24612 23492 24670
rect 23436 24546 23492 24556
rect 23996 24610 24052 26908
rect 24668 26962 24724 26974
rect 24668 26910 24670 26962
rect 24722 26910 24724 26962
rect 24556 26852 24612 26862
rect 24556 26758 24612 26796
rect 24108 26180 24164 26190
rect 24108 26086 24164 26124
rect 24332 26180 24388 26190
rect 24332 26178 24500 26180
rect 24332 26126 24334 26178
rect 24386 26126 24500 26178
rect 24332 26124 24500 26126
rect 24332 26114 24388 26124
rect 24108 25732 24164 25742
rect 24108 25638 24164 25676
rect 24220 25508 24276 25518
rect 24220 25414 24276 25452
rect 24108 25396 24164 25406
rect 24108 25302 24164 25340
rect 23996 24558 23998 24610
rect 24050 24558 24052 24610
rect 23436 23380 23492 23390
rect 23996 23380 24052 24558
rect 24444 25284 24500 26124
rect 24556 25844 24612 25854
rect 24556 25506 24612 25788
rect 24668 25620 24724 26910
rect 25116 26908 25172 33068
rect 25452 33058 25508 33068
rect 25452 30882 25508 30894
rect 25452 30830 25454 30882
rect 25506 30830 25508 30882
rect 25452 29988 25508 30830
rect 25788 30212 25844 30222
rect 25900 30212 25956 30222
rect 25788 30210 25900 30212
rect 25788 30158 25790 30210
rect 25842 30158 25900 30210
rect 25788 30156 25900 30158
rect 25788 30146 25844 30156
rect 25228 29538 25284 29550
rect 25228 29486 25230 29538
rect 25282 29486 25284 29538
rect 25228 29428 25284 29486
rect 25228 29362 25284 29372
rect 25452 28644 25508 29932
rect 25564 29652 25620 29662
rect 25564 29204 25620 29596
rect 25564 29138 25620 29148
rect 25452 28578 25508 28588
rect 25788 27858 25844 27870
rect 25788 27806 25790 27858
rect 25842 27806 25844 27858
rect 25788 27748 25844 27806
rect 25900 27748 25956 30156
rect 26348 29092 26404 47068
rect 26460 47012 26516 47022
rect 26460 46116 26516 46956
rect 26796 46562 26852 47292
rect 27244 47236 27300 47246
rect 27244 46898 27300 47180
rect 27244 46846 27246 46898
rect 27298 46846 27300 46898
rect 27244 46834 27300 46846
rect 26796 46510 26798 46562
rect 26850 46510 26852 46562
rect 26796 46498 26852 46510
rect 26460 46050 26516 46060
rect 27356 46114 27412 48188
rect 27468 48150 27524 48188
rect 27468 47458 27524 47470
rect 27468 47406 27470 47458
rect 27522 47406 27524 47458
rect 27468 47012 27524 47406
rect 27468 46946 27524 46956
rect 27356 46062 27358 46114
rect 27410 46062 27412 46114
rect 27356 46050 27412 46062
rect 27468 46674 27524 46686
rect 27468 46622 27470 46674
rect 27522 46622 27524 46674
rect 27244 45892 27300 45902
rect 27468 45892 27524 46622
rect 27244 45890 27524 45892
rect 27244 45838 27246 45890
rect 27298 45838 27524 45890
rect 27244 45836 27524 45838
rect 27132 42756 27188 42766
rect 27132 42662 27188 42700
rect 27244 42308 27300 45836
rect 27468 42756 27524 42766
rect 27132 42252 27300 42308
rect 27356 42754 27524 42756
rect 27356 42702 27470 42754
rect 27522 42702 27524 42754
rect 27356 42700 27524 42702
rect 26908 41970 26964 41982
rect 26908 41918 26910 41970
rect 26962 41918 26964 41970
rect 26908 41188 26964 41918
rect 27132 41410 27188 42252
rect 27244 42084 27300 42094
rect 27244 41990 27300 42028
rect 27132 41358 27134 41410
rect 27186 41358 27188 41410
rect 27132 41346 27188 41358
rect 26908 41122 26964 41132
rect 26460 41076 26516 41086
rect 26460 40982 26516 41020
rect 26572 41074 26628 41086
rect 26572 41022 26574 41074
rect 26626 41022 26628 41074
rect 26572 40852 26628 41022
rect 26572 40786 26628 40796
rect 26684 41074 26740 41086
rect 26684 41022 26686 41074
rect 26738 41022 26740 41074
rect 26460 39620 26516 39630
rect 26460 39526 26516 39564
rect 26684 39060 26740 41022
rect 27356 40964 27412 42700
rect 27468 42690 27524 42700
rect 27580 42308 27636 49644
rect 27692 48244 27748 48254
rect 27692 47236 27748 48188
rect 27916 48242 27972 48254
rect 27916 48190 27918 48242
rect 27970 48190 27972 48242
rect 27916 48020 27972 48190
rect 27916 47954 27972 47964
rect 28140 47908 28196 53564
rect 29036 53508 29092 53518
rect 28476 51378 28532 51390
rect 28476 51326 28478 51378
rect 28530 51326 28532 51378
rect 28252 50932 28308 50942
rect 28252 49924 28308 50876
rect 28364 50708 28420 50718
rect 28476 50708 28532 51326
rect 28364 50706 28532 50708
rect 28364 50654 28366 50706
rect 28418 50654 28532 50706
rect 28364 50652 28532 50654
rect 28588 51156 28644 51166
rect 28364 50642 28420 50652
rect 28588 50428 28644 51100
rect 28476 50372 28644 50428
rect 29036 50428 29092 53452
rect 29260 51378 29316 51390
rect 29260 51326 29262 51378
rect 29314 51326 29316 51378
rect 29260 51156 29316 51326
rect 29708 51266 29764 51278
rect 29708 51214 29710 51266
rect 29762 51214 29764 51266
rect 29316 51100 29540 51156
rect 29260 51090 29316 51100
rect 29372 50820 29428 50830
rect 29036 50372 29204 50428
rect 28476 50034 28532 50372
rect 28476 49982 28478 50034
rect 28530 49982 28532 50034
rect 28476 49970 28532 49982
rect 28812 50036 28868 50046
rect 28364 49924 28420 49934
rect 28252 49922 28420 49924
rect 28252 49870 28366 49922
rect 28418 49870 28420 49922
rect 28252 49868 28420 49870
rect 28364 49858 28420 49868
rect 28700 49812 28756 49822
rect 28700 49718 28756 49756
rect 28812 49810 28868 49980
rect 28812 49758 28814 49810
rect 28866 49758 28868 49810
rect 28812 49746 28868 49758
rect 28364 48356 28420 48366
rect 28420 48300 28644 48356
rect 28364 48262 28420 48300
rect 28252 48244 28308 48254
rect 28252 48150 28308 48188
rect 28364 48020 28420 48030
rect 28364 47926 28420 47964
rect 28140 47852 28308 47908
rect 27692 47170 27748 47180
rect 27916 45890 27972 45902
rect 27916 45838 27918 45890
rect 27970 45838 27972 45890
rect 27916 45108 27972 45838
rect 27916 45042 27972 45052
rect 27804 42868 27860 42878
rect 27692 42756 27748 42766
rect 27804 42756 27860 42812
rect 27692 42754 27860 42756
rect 27692 42702 27694 42754
rect 27746 42702 27860 42754
rect 27692 42700 27860 42702
rect 27692 42690 27748 42700
rect 27468 42252 27636 42308
rect 27468 41298 27524 42252
rect 27692 41748 27748 41758
rect 27468 41246 27470 41298
rect 27522 41246 27524 41298
rect 27468 41234 27524 41246
rect 27580 41746 27748 41748
rect 27580 41694 27694 41746
rect 27746 41694 27748 41746
rect 27580 41692 27748 41694
rect 27804 41748 27860 42700
rect 27916 42196 27972 42206
rect 27916 41970 27972 42140
rect 27916 41918 27918 41970
rect 27970 41918 27972 41970
rect 27916 41906 27972 41918
rect 28028 42194 28084 42206
rect 28028 42142 28030 42194
rect 28082 42142 28084 42194
rect 28028 41972 28084 42142
rect 28028 41906 28084 41916
rect 28140 41970 28196 41982
rect 28140 41918 28142 41970
rect 28194 41918 28196 41970
rect 27804 41692 27972 41748
rect 27580 41300 27636 41692
rect 27692 41682 27748 41692
rect 27356 40898 27412 40908
rect 27468 40962 27524 40974
rect 27468 40910 27470 40962
rect 27522 40910 27524 40962
rect 27468 40628 27524 40910
rect 27580 40740 27636 41244
rect 27804 41412 27860 41422
rect 27692 40964 27748 40974
rect 27804 40964 27860 41356
rect 27692 40962 27860 40964
rect 27692 40910 27694 40962
rect 27746 40910 27860 40962
rect 27692 40908 27860 40910
rect 27692 40898 27748 40908
rect 27804 40740 27860 40908
rect 27580 40684 27748 40740
rect 27468 40562 27524 40572
rect 27132 40402 27188 40414
rect 27132 40350 27134 40402
rect 27186 40350 27188 40402
rect 26908 39172 26964 39182
rect 27132 39172 27188 40350
rect 27580 40404 27636 40414
rect 27580 40292 27636 40348
rect 26964 39116 27188 39172
rect 27244 40290 27636 40292
rect 27244 40238 27582 40290
rect 27634 40238 27636 40290
rect 27244 40236 27636 40238
rect 26908 39106 26964 39116
rect 26684 38994 26740 39004
rect 26572 38948 26628 38958
rect 26572 38610 26628 38892
rect 27020 38834 27076 39116
rect 27020 38782 27022 38834
rect 27074 38782 27076 38834
rect 27020 38770 27076 38782
rect 27244 38834 27300 40236
rect 27580 40226 27636 40236
rect 27692 40068 27748 40684
rect 27804 40402 27860 40684
rect 27804 40350 27806 40402
rect 27858 40350 27860 40402
rect 27804 40338 27860 40350
rect 27580 40012 27748 40068
rect 27468 39396 27524 39406
rect 27468 39302 27524 39340
rect 27244 38782 27246 38834
rect 27298 38782 27300 38834
rect 26908 38724 26964 38734
rect 26908 38630 26964 38668
rect 26572 38558 26574 38610
rect 26626 38558 26628 38610
rect 26572 38546 26628 38558
rect 27020 38164 27076 38174
rect 27020 38070 27076 38108
rect 26572 38052 26628 38062
rect 26572 37266 26628 37996
rect 27132 38050 27188 38062
rect 27132 37998 27134 38050
rect 27186 37998 27188 38050
rect 26572 37214 26574 37266
rect 26626 37214 26628 37266
rect 26572 37202 26628 37214
rect 26796 37378 26852 37390
rect 26796 37326 26798 37378
rect 26850 37326 26852 37378
rect 26796 37268 26852 37326
rect 26796 37202 26852 37212
rect 27132 37380 27188 37998
rect 27132 37266 27188 37324
rect 27132 37214 27134 37266
rect 27186 37214 27188 37266
rect 27132 37202 27188 37214
rect 27244 37042 27300 38782
rect 27244 36990 27246 37042
rect 27298 36990 27300 37042
rect 27244 36978 27300 36990
rect 27356 38612 27412 38622
rect 27356 36706 27412 38556
rect 27580 38162 27636 40012
rect 27916 39730 27972 41692
rect 28140 41412 28196 41918
rect 28140 41346 28196 41356
rect 28028 41188 28084 41198
rect 28028 41186 28196 41188
rect 28028 41134 28030 41186
rect 28082 41134 28196 41186
rect 28028 41132 28196 41134
rect 28028 41122 28084 41132
rect 28140 40964 28196 41132
rect 28028 40740 28084 40750
rect 28028 40290 28084 40684
rect 28028 40238 28030 40290
rect 28082 40238 28084 40290
rect 28028 40226 28084 40238
rect 27916 39678 27918 39730
rect 27970 39678 27972 39730
rect 27916 39666 27972 39678
rect 27916 39396 27972 39406
rect 27692 39060 27748 39070
rect 27692 38966 27748 39004
rect 27916 39058 27972 39340
rect 27916 39006 27918 39058
rect 27970 39006 27972 39058
rect 27916 38994 27972 39006
rect 28028 38836 28084 38846
rect 28028 38742 28084 38780
rect 27580 38110 27582 38162
rect 27634 38110 27636 38162
rect 27580 38098 27636 38110
rect 28140 38162 28196 40908
rect 28140 38110 28142 38162
rect 28194 38110 28196 38162
rect 28140 38098 28196 38110
rect 27468 38052 27524 38062
rect 27468 37958 27524 37996
rect 27580 37940 27636 37950
rect 27580 37492 27636 37884
rect 28140 37940 28196 37950
rect 28140 37846 28196 37884
rect 27580 37266 27636 37436
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 37202 27636 37214
rect 27356 36654 27358 36706
rect 27410 36654 27412 36706
rect 27356 36642 27412 36654
rect 27020 36594 27076 36606
rect 27020 36542 27022 36594
rect 27074 36542 27076 36594
rect 26908 36482 26964 36494
rect 26908 36430 26910 36482
rect 26962 36430 26964 36482
rect 26908 36372 26964 36430
rect 27020 36484 27076 36542
rect 27076 36428 27300 36484
rect 27020 36418 27076 36428
rect 26908 36306 26964 36316
rect 27244 35922 27300 36428
rect 27804 36260 27860 36270
rect 27244 35870 27246 35922
rect 27298 35870 27300 35922
rect 27244 35858 27300 35870
rect 27580 36258 27860 36260
rect 27580 36206 27806 36258
rect 27858 36206 27860 36258
rect 27580 36204 27860 36206
rect 27356 35812 27412 35822
rect 27580 35812 27636 36204
rect 27804 36194 27860 36204
rect 28252 35924 28308 47852
rect 28476 47572 28532 47582
rect 28476 47478 28532 47516
rect 28588 46786 28644 48300
rect 28588 46734 28590 46786
rect 28642 46734 28644 46786
rect 28588 46564 28644 46734
rect 28700 46788 28756 46798
rect 28700 46694 28756 46732
rect 28924 46676 28980 46686
rect 28924 46674 29092 46676
rect 28924 46622 28926 46674
rect 28978 46622 29092 46674
rect 28924 46620 29092 46622
rect 28924 46610 28980 46620
rect 28588 46508 28756 46564
rect 28588 45666 28644 45678
rect 28588 45614 28590 45666
rect 28642 45614 28644 45666
rect 28476 45108 28532 45118
rect 28588 45108 28644 45614
rect 28700 45330 28756 46508
rect 29036 45890 29092 46620
rect 29036 45838 29038 45890
rect 29090 45838 29092 45890
rect 29036 45826 29092 45838
rect 29148 45892 29204 50372
rect 29372 50034 29428 50764
rect 29484 50594 29540 51100
rect 29708 50932 29764 51214
rect 29820 51154 29876 54460
rect 30380 54068 30436 54684
rect 30940 54628 30996 55246
rect 30828 54572 30940 54628
rect 30828 54514 30884 54572
rect 30940 54562 30996 54572
rect 30828 54462 30830 54514
rect 30882 54462 30884 54514
rect 30380 53618 30436 54012
rect 30380 53566 30382 53618
rect 30434 53566 30436 53618
rect 30380 53554 30436 53566
rect 30604 54402 30660 54414
rect 30604 54350 30606 54402
rect 30658 54350 30660 54402
rect 30044 53508 30100 53518
rect 30044 53414 30100 53452
rect 30604 53508 30660 54350
rect 30604 53442 30660 53452
rect 30716 53732 30772 53742
rect 30716 52836 30772 53676
rect 30828 52836 30884 54462
rect 30828 52780 31108 52836
rect 30716 52050 30772 52780
rect 30940 52276 30996 52286
rect 30940 52164 30996 52220
rect 30716 51998 30718 52050
rect 30770 51998 30772 52050
rect 30716 51986 30772 51998
rect 30828 52162 30996 52164
rect 30828 52110 30942 52162
rect 30994 52110 30996 52162
rect 30828 52108 30996 52110
rect 29820 51102 29822 51154
rect 29874 51102 29876 51154
rect 29820 51090 29876 51102
rect 30044 51378 30100 51390
rect 30044 51326 30046 51378
rect 30098 51326 30100 51378
rect 29708 50706 29764 50876
rect 29708 50654 29710 50706
rect 29762 50654 29764 50706
rect 29708 50642 29764 50654
rect 29820 50708 29876 50718
rect 29484 50542 29486 50594
rect 29538 50542 29540 50594
rect 29484 50530 29540 50542
rect 29596 50596 29652 50606
rect 29372 49982 29374 50034
rect 29426 49982 29428 50034
rect 29372 49970 29428 49982
rect 29484 50036 29540 50046
rect 29596 50036 29652 50540
rect 29820 50036 29876 50652
rect 29932 50036 29988 50046
rect 29484 50034 29652 50036
rect 29484 49982 29486 50034
rect 29538 49982 29652 50034
rect 29484 49980 29652 49982
rect 29708 50034 29988 50036
rect 29708 49982 29934 50034
rect 29986 49982 29988 50034
rect 29708 49980 29988 49982
rect 30044 50036 30100 51326
rect 30716 50708 30772 50718
rect 30156 50596 30212 50606
rect 30380 50596 30436 50606
rect 30212 50594 30436 50596
rect 30212 50542 30382 50594
rect 30434 50542 30436 50594
rect 30212 50540 30436 50542
rect 30156 50502 30212 50540
rect 30380 50530 30436 50540
rect 30716 50594 30772 50652
rect 30716 50542 30718 50594
rect 30770 50542 30772 50594
rect 30716 50530 30772 50542
rect 30604 50484 30660 50522
rect 30604 50418 30660 50428
rect 30828 50372 30884 52108
rect 30940 52098 30996 52108
rect 30940 50820 30996 50830
rect 30940 50594 30996 50764
rect 30940 50542 30942 50594
rect 30994 50542 30996 50594
rect 30940 50530 30996 50542
rect 30716 50316 30884 50372
rect 30156 50036 30212 50046
rect 30044 50034 30212 50036
rect 30044 49982 30158 50034
rect 30210 49982 30212 50034
rect 30044 49980 30212 49982
rect 29484 49970 29540 49980
rect 29260 49812 29316 49822
rect 29708 49812 29764 49980
rect 29932 49970 29988 49980
rect 30156 49970 30212 49980
rect 30492 50036 30548 50046
rect 29260 49810 29764 49812
rect 29260 49758 29262 49810
rect 29314 49758 29764 49810
rect 29260 49756 29764 49758
rect 29820 49812 29876 49822
rect 29260 46114 29316 49756
rect 29820 49718 29876 49756
rect 30492 49140 30548 49980
rect 30492 49074 30548 49084
rect 29372 48356 29428 48366
rect 29372 47682 29428 48300
rect 29372 47630 29374 47682
rect 29426 47630 29428 47682
rect 29372 46562 29428 47630
rect 29372 46510 29374 46562
rect 29426 46510 29428 46562
rect 29372 46498 29428 46510
rect 29484 47234 29540 47246
rect 29484 47182 29486 47234
rect 29538 47182 29540 47234
rect 29260 46062 29262 46114
rect 29314 46062 29316 46114
rect 29260 46050 29316 46062
rect 29484 46004 29540 47182
rect 29596 47236 29652 47246
rect 29596 47234 29876 47236
rect 29596 47182 29598 47234
rect 29650 47182 29876 47234
rect 29596 47180 29876 47182
rect 29596 47170 29652 47180
rect 29820 46788 29876 47180
rect 29708 46004 29764 46014
rect 29484 46002 29764 46004
rect 29484 45950 29710 46002
rect 29762 45950 29764 46002
rect 29484 45948 29764 45950
rect 29708 45938 29764 45948
rect 29820 46004 29876 46732
rect 29820 45938 29876 45948
rect 30156 46228 30212 46238
rect 29148 45836 29428 45892
rect 28700 45278 28702 45330
rect 28754 45278 28756 45330
rect 28700 45266 28756 45278
rect 28532 45052 28644 45108
rect 29148 45108 29204 45118
rect 28476 45014 28532 45052
rect 29148 44994 29204 45052
rect 29148 44942 29150 44994
rect 29202 44942 29204 44994
rect 28364 43540 28420 43550
rect 28364 42754 28420 43484
rect 29148 42980 29204 44942
rect 29372 43708 29428 45836
rect 30156 45890 30212 46172
rect 30156 45838 30158 45890
rect 30210 45838 30212 45890
rect 30156 45826 30212 45838
rect 30156 44996 30212 45006
rect 29372 43652 29540 43708
rect 29148 42924 29428 42980
rect 28364 42702 28366 42754
rect 28418 42702 28420 42754
rect 28364 42196 28420 42702
rect 29148 42756 29204 42766
rect 29148 42662 29204 42700
rect 28476 42532 28532 42542
rect 28588 42532 28644 42542
rect 28476 42530 28588 42532
rect 28476 42478 28478 42530
rect 28530 42478 28588 42530
rect 28476 42476 28588 42478
rect 28476 42466 28532 42476
rect 28588 42308 28644 42476
rect 28700 42532 28756 42542
rect 29260 42532 29316 42542
rect 28700 42530 29316 42532
rect 28700 42478 28702 42530
rect 28754 42478 29262 42530
rect 29314 42478 29316 42530
rect 28700 42476 29316 42478
rect 28700 42466 28756 42476
rect 29260 42466 29316 42476
rect 29372 42308 29428 42924
rect 29484 42530 29540 43652
rect 29820 43652 29876 43662
rect 29820 43558 29876 43596
rect 29708 43538 29764 43550
rect 29708 43486 29710 43538
rect 29762 43486 29764 43538
rect 29708 42868 29764 43486
rect 29932 43540 29988 43550
rect 29932 43446 29988 43484
rect 30156 43540 30212 44940
rect 30716 43708 30772 50316
rect 31052 50260 31108 52780
rect 30380 43652 30772 43708
rect 30828 50204 31108 50260
rect 30156 43474 30212 43484
rect 30268 43538 30324 43550
rect 30268 43486 30270 43538
rect 30322 43486 30324 43538
rect 29708 42802 29764 42812
rect 29484 42478 29486 42530
rect 29538 42478 29540 42530
rect 29484 42466 29540 42478
rect 30044 42754 30100 42766
rect 30044 42702 30046 42754
rect 30098 42702 30100 42754
rect 28588 42252 28756 42308
rect 29372 42252 29652 42308
rect 28476 42196 28532 42206
rect 28420 42194 28532 42196
rect 28420 42142 28478 42194
rect 28530 42142 28532 42194
rect 28420 42140 28532 42142
rect 28364 42102 28420 42140
rect 28476 42130 28532 42140
rect 28588 42084 28644 42094
rect 28588 41970 28644 42028
rect 28588 41918 28590 41970
rect 28642 41918 28644 41970
rect 28588 41906 28644 41918
rect 28700 41970 28756 42252
rect 28700 41918 28702 41970
rect 28754 41918 28756 41970
rect 28588 41748 28644 41758
rect 28588 39956 28644 41692
rect 28700 40964 28756 41918
rect 29036 41970 29092 41982
rect 29036 41918 29038 41970
rect 29090 41918 29092 41970
rect 29036 41186 29092 41918
rect 29484 41972 29540 41982
rect 29484 41878 29540 41916
rect 29036 41134 29038 41186
rect 29090 41134 29092 41186
rect 29036 41122 29092 41134
rect 29372 41074 29428 41086
rect 29372 41022 29374 41074
rect 29426 41022 29428 41074
rect 29260 40964 29316 40974
rect 28700 40962 29316 40964
rect 28700 40910 29262 40962
rect 29314 40910 29316 40962
rect 28700 40908 29316 40910
rect 28924 40628 28980 40638
rect 28924 40402 28980 40572
rect 28924 40350 28926 40402
rect 28978 40350 28980 40402
rect 28924 40338 28980 40350
rect 28588 39890 28644 39900
rect 29148 38276 29204 40908
rect 29260 40898 29316 40908
rect 29372 40628 29428 41022
rect 29260 40572 29428 40628
rect 29260 40402 29316 40572
rect 29260 40350 29262 40402
rect 29314 40350 29316 40402
rect 29260 38612 29316 40350
rect 29372 40404 29428 40414
rect 29372 40290 29428 40348
rect 29372 40238 29374 40290
rect 29426 40238 29428 40290
rect 29372 40226 29428 40238
rect 29260 38546 29316 38556
rect 29260 38276 29316 38286
rect 29148 38274 29316 38276
rect 29148 38222 29262 38274
rect 29314 38222 29316 38274
rect 29148 38220 29316 38222
rect 29260 38210 29316 38220
rect 28588 38052 28644 38062
rect 28476 37996 28588 38052
rect 28364 37828 28420 37838
rect 28364 37734 28420 37772
rect 28364 36596 28420 36606
rect 28476 36596 28532 37996
rect 28588 37958 28644 37996
rect 29148 38052 29204 38062
rect 29148 37266 29204 37996
rect 29260 37940 29316 37950
rect 29260 37846 29316 37884
rect 29372 37938 29428 37950
rect 29372 37886 29374 37938
rect 29426 37886 29428 37938
rect 29148 37214 29150 37266
rect 29202 37214 29204 37266
rect 29148 37202 29204 37214
rect 29260 37268 29316 37278
rect 29372 37268 29428 37886
rect 29316 37212 29428 37268
rect 28364 36594 28532 36596
rect 28364 36542 28366 36594
rect 28418 36542 28532 36594
rect 28364 36540 28532 36542
rect 28364 36530 28420 36540
rect 28364 35924 28420 35934
rect 28252 35922 28420 35924
rect 28252 35870 28366 35922
rect 28418 35870 28420 35922
rect 28252 35868 28420 35870
rect 27356 35810 27636 35812
rect 27356 35758 27358 35810
rect 27410 35758 27636 35810
rect 27356 35756 27636 35758
rect 27356 35588 27412 35756
rect 27356 35522 27412 35532
rect 28364 35028 28420 35868
rect 28364 34934 28420 34972
rect 29148 35028 29204 35038
rect 27916 34914 27972 34926
rect 27916 34862 27918 34914
rect 27970 34862 27972 34914
rect 27580 34692 27636 34702
rect 27916 34692 27972 34862
rect 27468 34690 27972 34692
rect 27468 34638 27582 34690
rect 27634 34638 27972 34690
rect 27468 34636 27972 34638
rect 27468 33236 27524 34636
rect 27580 34626 27636 34636
rect 27916 34356 27972 34636
rect 27916 34290 27972 34300
rect 29148 34354 29204 34972
rect 29148 34302 29150 34354
rect 29202 34302 29204 34354
rect 29148 34290 29204 34302
rect 28364 34132 28420 34142
rect 28364 34130 28532 34132
rect 28364 34078 28366 34130
rect 28418 34078 28532 34130
rect 28364 34076 28532 34078
rect 28364 34066 28420 34076
rect 27580 34020 27636 34030
rect 27580 34018 27972 34020
rect 27580 33966 27582 34018
rect 27634 33966 27972 34018
rect 27580 33964 27972 33966
rect 27580 33954 27636 33964
rect 27916 33458 27972 33964
rect 27916 33406 27918 33458
rect 27970 33406 27972 33458
rect 27916 33394 27972 33406
rect 28364 33684 28420 33694
rect 28140 33348 28196 33358
rect 28140 33254 28196 33292
rect 28364 33346 28420 33628
rect 28364 33294 28366 33346
rect 28418 33294 28420 33346
rect 28364 33282 28420 33294
rect 27468 33170 27524 33180
rect 27804 33234 27860 33246
rect 27804 33182 27806 33234
rect 27858 33182 27860 33234
rect 27580 33124 27636 33134
rect 27804 33124 27860 33182
rect 27580 33122 27804 33124
rect 27580 33070 27582 33122
rect 27634 33070 27804 33122
rect 27580 33068 27804 33070
rect 27580 33058 27636 33068
rect 27804 33058 27860 33068
rect 28476 32452 28532 34076
rect 28700 34130 28756 34142
rect 28700 34078 28702 34130
rect 28754 34078 28756 34130
rect 28700 33124 28756 34078
rect 28924 34132 28980 34142
rect 29260 34132 29316 37212
rect 29596 35252 29652 42252
rect 30044 42084 30100 42702
rect 30044 42018 30100 42028
rect 29708 41970 29764 41982
rect 29708 41918 29710 41970
rect 29762 41918 29764 41970
rect 29708 40628 29764 41918
rect 29708 40562 29764 40572
rect 30268 40516 30324 43486
rect 30380 41970 30436 43652
rect 30380 41918 30382 41970
rect 30434 41918 30436 41970
rect 30380 41906 30436 41918
rect 30604 42642 30660 42654
rect 30604 42590 30606 42642
rect 30658 42590 30660 42642
rect 30604 41412 30660 42590
rect 30604 41346 30660 41356
rect 30268 40450 30324 40460
rect 30828 39844 30884 50204
rect 31164 49924 31220 57820
rect 31276 54404 31332 60620
rect 31612 60676 31668 60686
rect 31948 60676 32004 60734
rect 31612 60674 32004 60676
rect 31612 60622 31614 60674
rect 31666 60622 32004 60674
rect 31612 60620 32004 60622
rect 31388 60004 31444 60014
rect 31612 60004 31668 60620
rect 32060 60564 32116 60574
rect 32060 60114 32116 60508
rect 32060 60062 32062 60114
rect 32114 60062 32116 60114
rect 32060 60050 32116 60062
rect 31388 60002 31668 60004
rect 31388 59950 31390 60002
rect 31442 59950 31668 60002
rect 31388 59948 31668 59950
rect 31388 59108 31444 59948
rect 32284 59668 32340 60958
rect 32508 60226 32564 61292
rect 32620 61282 32676 61292
rect 32508 60174 32510 60226
rect 32562 60174 32564 60226
rect 32508 60162 32564 60174
rect 32844 60002 32900 61404
rect 32844 59950 32846 60002
rect 32898 59950 32900 60002
rect 32844 59938 32900 59950
rect 32396 59892 32452 59902
rect 32396 59798 32452 59836
rect 32508 59778 32564 59790
rect 32508 59726 32510 59778
rect 32562 59726 32564 59778
rect 32508 59668 32564 59726
rect 32284 59612 32564 59668
rect 31388 59042 31444 59052
rect 32284 59108 32340 59118
rect 31612 57540 31668 57550
rect 32060 57540 32116 57550
rect 31612 57538 32116 57540
rect 31612 57486 31614 57538
rect 31666 57486 32062 57538
rect 32114 57486 32116 57538
rect 31612 57484 32116 57486
rect 31612 57474 31668 57484
rect 32060 57474 32116 57484
rect 31612 57316 31668 57326
rect 31612 56978 31668 57260
rect 32284 57092 32340 59052
rect 32956 57876 33012 62188
rect 33740 62132 33908 62188
rect 35868 62356 35924 62366
rect 33404 60788 33460 60798
rect 33292 60786 33460 60788
rect 33292 60734 33406 60786
rect 33458 60734 33460 60786
rect 33292 60732 33460 60734
rect 33180 60674 33236 60686
rect 33180 60622 33182 60674
rect 33234 60622 33236 60674
rect 33180 60340 33236 60622
rect 33180 60274 33236 60284
rect 33292 60564 33348 60732
rect 33404 60722 33460 60732
rect 33292 60116 33348 60508
rect 33068 60060 33348 60116
rect 33404 60340 33460 60350
rect 33068 59890 33124 60060
rect 33068 59838 33070 59890
rect 33122 59838 33124 59890
rect 33068 59826 33124 59838
rect 33180 59892 33236 59902
rect 33404 59892 33460 60284
rect 33628 60004 33684 60014
rect 33628 59910 33684 59948
rect 33180 59890 33460 59892
rect 33180 59838 33182 59890
rect 33234 59838 33460 59890
rect 33180 59836 33460 59838
rect 33180 59826 33236 59836
rect 32956 57820 33460 57876
rect 32396 57652 32452 57690
rect 32396 57586 32452 57596
rect 33180 57652 33236 57662
rect 33180 57538 33236 57596
rect 33180 57486 33182 57538
rect 33234 57486 33236 57538
rect 32284 57026 32340 57036
rect 32396 57426 32452 57438
rect 32396 57374 32398 57426
rect 32450 57374 32452 57426
rect 31612 56926 31614 56978
rect 31666 56926 31668 56978
rect 31612 56914 31668 56926
rect 32396 56980 32452 57374
rect 32396 56914 32452 56924
rect 31836 56196 31892 56206
rect 31724 56194 31892 56196
rect 31724 56142 31838 56194
rect 31890 56142 31892 56194
rect 31724 56140 31892 56142
rect 31388 55970 31444 55982
rect 31388 55918 31390 55970
rect 31442 55918 31444 55970
rect 31388 55858 31444 55918
rect 31388 55806 31390 55858
rect 31442 55806 31444 55858
rect 31388 55794 31444 55806
rect 31724 55298 31780 56140
rect 31836 56130 31892 56140
rect 32508 56196 32564 56206
rect 32508 56102 32564 56140
rect 32284 56082 32340 56094
rect 32284 56030 32286 56082
rect 32338 56030 32340 56082
rect 32284 55522 32340 56030
rect 32284 55470 32286 55522
rect 32338 55470 32340 55522
rect 32284 55458 32340 55470
rect 33068 55410 33124 55422
rect 33068 55358 33070 55410
rect 33122 55358 33124 55410
rect 31724 55246 31726 55298
rect 31778 55246 31780 55298
rect 31724 55234 31780 55246
rect 32956 55298 33012 55310
rect 32956 55246 32958 55298
rect 33010 55246 33012 55298
rect 31388 55186 31444 55198
rect 31388 55134 31390 55186
rect 31442 55134 31444 55186
rect 31388 54740 31444 55134
rect 31612 55188 31668 55198
rect 31500 55076 31556 55086
rect 31500 54982 31556 55020
rect 31388 54674 31444 54684
rect 31500 54628 31556 54638
rect 31612 54628 31668 55132
rect 32284 55188 32340 55198
rect 32284 55094 32340 55132
rect 32396 55188 32452 55198
rect 32956 55188 33012 55246
rect 32396 55186 33012 55188
rect 32396 55134 32398 55186
rect 32450 55134 33012 55186
rect 32396 55132 33012 55134
rect 33068 55188 33124 55358
rect 31500 54626 31668 54628
rect 31500 54574 31502 54626
rect 31554 54574 31668 54626
rect 31500 54572 31668 54574
rect 31948 54628 32004 54638
rect 31500 54562 31556 54572
rect 31948 54534 32004 54572
rect 31276 54348 31556 54404
rect 31276 53956 31332 53966
rect 31276 53172 31332 53900
rect 31276 53078 31332 53116
rect 31500 50428 31556 54348
rect 32396 54292 32452 55132
rect 33068 55122 33124 55132
rect 33180 54964 33236 57486
rect 32396 54226 32452 54236
rect 33068 54908 33236 54964
rect 32172 53172 32228 53182
rect 31612 52948 31668 52958
rect 31612 52946 31892 52948
rect 31612 52894 31614 52946
rect 31666 52894 31892 52946
rect 31612 52892 31892 52894
rect 31612 52882 31668 52892
rect 31836 52164 31892 52892
rect 32172 52946 32228 53116
rect 32172 52894 32174 52946
rect 32226 52894 32228 52946
rect 32172 52882 32228 52894
rect 31948 52836 32004 52846
rect 31948 52742 32004 52780
rect 32508 52724 32564 52734
rect 32508 52722 32788 52724
rect 32508 52670 32510 52722
rect 32562 52670 32788 52722
rect 32508 52668 32788 52670
rect 32508 52658 32564 52668
rect 32508 52500 32564 52510
rect 31836 52098 31892 52108
rect 31948 52276 32004 52286
rect 31948 52162 32004 52220
rect 32396 52276 32452 52286
rect 32396 52182 32452 52220
rect 31948 52110 31950 52162
rect 32002 52110 32004 52162
rect 31948 52098 32004 52110
rect 32284 52164 32340 52174
rect 32284 52070 32340 52108
rect 32508 51602 32564 52444
rect 32732 52162 32788 52668
rect 32732 52110 32734 52162
rect 32786 52110 32788 52162
rect 32732 52098 32788 52110
rect 32508 51550 32510 51602
rect 32562 51550 32564 51602
rect 32508 51538 32564 51550
rect 32284 50932 32340 50942
rect 32284 50594 32340 50876
rect 32284 50542 32286 50594
rect 32338 50542 32340 50594
rect 32284 50428 32340 50542
rect 32508 50594 32564 50606
rect 32508 50542 32510 50594
rect 32562 50542 32564 50594
rect 31500 50372 31892 50428
rect 32284 50372 32452 50428
rect 30940 49868 31220 49924
rect 30940 42978 30996 49868
rect 31500 49810 31556 49822
rect 31500 49758 31502 49810
rect 31554 49758 31556 49810
rect 31164 49700 31220 49710
rect 31164 49606 31220 49644
rect 31500 49028 31556 49758
rect 31276 49026 31556 49028
rect 31276 48974 31502 49026
rect 31554 48974 31556 49026
rect 31276 48972 31556 48974
rect 31164 46786 31220 46798
rect 31164 46734 31166 46786
rect 31218 46734 31220 46786
rect 31164 46228 31220 46734
rect 31164 46162 31220 46172
rect 31052 46004 31108 46014
rect 31052 45910 31108 45948
rect 31164 44324 31220 44334
rect 31164 44210 31220 44268
rect 31164 44158 31166 44210
rect 31218 44158 31220 44210
rect 31164 44146 31220 44158
rect 31276 43652 31332 48972
rect 31500 48962 31556 48972
rect 31388 46564 31444 46574
rect 31724 46564 31780 46574
rect 31388 46562 31780 46564
rect 31388 46510 31390 46562
rect 31442 46510 31726 46562
rect 31778 46510 31780 46562
rect 31388 46508 31780 46510
rect 31388 46498 31444 46508
rect 31724 46498 31780 46508
rect 31836 46340 31892 50372
rect 32060 49810 32116 49822
rect 32060 49758 32062 49810
rect 32114 49758 32116 49810
rect 32060 49028 32116 49758
rect 32396 49698 32452 50372
rect 32508 49924 32564 50542
rect 32508 49858 32564 49868
rect 32396 49646 32398 49698
rect 32450 49646 32452 49698
rect 32396 49634 32452 49646
rect 32732 49812 32788 49822
rect 32732 49140 32788 49756
rect 32956 49140 33012 49150
rect 32396 49138 32788 49140
rect 32396 49086 32734 49138
rect 32786 49086 32788 49138
rect 32396 49084 32788 49086
rect 32172 49028 32228 49038
rect 32060 49026 32340 49028
rect 32060 48974 32174 49026
rect 32226 48974 32340 49026
rect 32060 48972 32340 48974
rect 32172 48962 32228 48972
rect 32060 46900 32116 46910
rect 32060 46674 32116 46844
rect 32060 46622 32062 46674
rect 32114 46622 32116 46674
rect 32060 46610 32116 46622
rect 31612 46284 31892 46340
rect 32060 46450 32116 46462
rect 32060 46398 32062 46450
rect 32114 46398 32116 46450
rect 31388 44322 31444 44334
rect 31388 44270 31390 44322
rect 31442 44270 31444 44322
rect 31388 44212 31444 44270
rect 31388 44146 31444 44156
rect 31276 43586 31332 43596
rect 30940 42926 30942 42978
rect 30994 42926 30996 42978
rect 30940 42914 30996 42926
rect 31276 42868 31332 42878
rect 31332 42812 31444 42868
rect 31276 42774 31332 42812
rect 30940 42754 30996 42766
rect 30940 42702 30942 42754
rect 30994 42702 30996 42754
rect 30940 42532 30996 42702
rect 30940 42466 30996 42476
rect 31164 40516 31220 40526
rect 31164 40290 31220 40460
rect 31388 40402 31444 42812
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 31388 40338 31444 40350
rect 31164 40238 31166 40290
rect 31218 40238 31220 40290
rect 31164 40226 31220 40238
rect 30828 39788 31444 39844
rect 31276 39620 31332 39630
rect 30380 39618 31332 39620
rect 30380 39566 31278 39618
rect 31330 39566 31332 39618
rect 30380 39564 31332 39566
rect 30044 39060 30100 39070
rect 30044 38834 30100 39004
rect 30380 38946 30436 39564
rect 31276 39554 31332 39564
rect 30828 39396 30884 39406
rect 30380 38894 30382 38946
rect 30434 38894 30436 38946
rect 30380 38882 30436 38894
rect 30716 39340 30828 39396
rect 30604 38836 30660 38846
rect 30044 38782 30046 38834
rect 30098 38782 30100 38834
rect 30044 38770 30100 38782
rect 30492 38834 30660 38836
rect 30492 38782 30606 38834
rect 30658 38782 30660 38834
rect 30492 38780 30660 38782
rect 29932 38724 29988 38734
rect 29932 38630 29988 38668
rect 30268 38610 30324 38622
rect 30268 38558 30270 38610
rect 30322 38558 30324 38610
rect 30268 37268 30324 38558
rect 30492 38274 30548 38780
rect 30604 38770 30660 38780
rect 30492 38222 30494 38274
rect 30546 38222 30548 38274
rect 30492 38210 30548 38222
rect 30604 37940 30660 37950
rect 30604 37846 30660 37884
rect 30268 37202 30324 37212
rect 30492 37826 30548 37838
rect 30492 37774 30494 37826
rect 30546 37774 30548 37826
rect 30156 36148 30212 36158
rect 29596 35186 29652 35196
rect 29708 35700 29764 35710
rect 29708 35026 29764 35644
rect 29708 34974 29710 35026
rect 29762 34974 29764 35026
rect 29708 34962 29764 34974
rect 29932 34916 29988 34926
rect 29820 34804 29876 34814
rect 29820 34710 29876 34748
rect 29372 34692 29428 34702
rect 29596 34692 29652 34702
rect 29372 34690 29540 34692
rect 29372 34638 29374 34690
rect 29426 34638 29540 34690
rect 29372 34636 29540 34638
rect 29372 34626 29428 34636
rect 28924 34130 29316 34132
rect 28924 34078 28926 34130
rect 28978 34078 29316 34130
rect 28924 34076 29316 34078
rect 29484 34132 29540 34636
rect 29596 34598 29652 34636
rect 29820 34356 29876 34366
rect 29932 34356 29988 34860
rect 29820 34354 29988 34356
rect 29820 34302 29822 34354
rect 29874 34302 29988 34354
rect 29820 34300 29988 34302
rect 29820 34290 29876 34300
rect 30044 34132 30100 34142
rect 29484 34130 30100 34132
rect 29484 34078 30046 34130
rect 30098 34078 30100 34130
rect 29484 34076 30100 34078
rect 28812 34018 28868 34030
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33684 28868 33966
rect 28812 33618 28868 33628
rect 28924 33348 28980 34076
rect 30044 34066 30100 34076
rect 28924 33282 28980 33292
rect 28700 33058 28756 33068
rect 29372 33124 29428 33134
rect 29484 33124 29540 33134
rect 29428 33122 29540 33124
rect 29428 33070 29486 33122
rect 29538 33070 29540 33122
rect 29428 33068 29540 33070
rect 28588 32452 28644 32462
rect 28476 32450 28644 32452
rect 28476 32398 28590 32450
rect 28642 32398 28644 32450
rect 28476 32396 28644 32398
rect 26796 31892 26852 31902
rect 26796 31798 26852 31836
rect 27244 31554 27300 31566
rect 27244 31502 27246 31554
rect 27298 31502 27300 31554
rect 27244 30884 27300 31502
rect 28140 30996 28196 31006
rect 28588 30996 28644 32396
rect 28812 31668 28868 31678
rect 28140 30994 28644 30996
rect 28140 30942 28142 30994
rect 28194 30942 28644 30994
rect 28140 30940 28644 30942
rect 28700 31612 28812 31668
rect 27692 30884 27748 30894
rect 28140 30884 28196 30940
rect 27244 30882 28196 30884
rect 27244 30830 27694 30882
rect 27746 30830 28196 30882
rect 27244 30828 28196 30830
rect 27692 30818 27748 30828
rect 28140 30212 28196 30828
rect 28588 30324 28644 30334
rect 28700 30324 28756 31612
rect 28812 31602 28868 31612
rect 28812 30884 28868 30894
rect 28812 30882 29204 30884
rect 28812 30830 28814 30882
rect 28866 30830 29204 30882
rect 28812 30828 29204 30830
rect 28812 30818 28868 30828
rect 28588 30322 28756 30324
rect 28588 30270 28590 30322
rect 28642 30270 28756 30322
rect 28588 30268 28756 30270
rect 28588 30258 28644 30268
rect 26460 30098 26516 30110
rect 26460 30046 26462 30098
rect 26514 30046 26516 30098
rect 26460 29316 26516 30046
rect 26460 29250 26516 29260
rect 26908 29652 26964 29662
rect 26348 29026 26404 29036
rect 26908 28980 26964 29596
rect 27804 29652 27860 29662
rect 27804 29558 27860 29596
rect 28028 29652 28084 29662
rect 28028 29558 28084 29596
rect 27580 29538 27636 29550
rect 27580 29486 27582 29538
rect 27634 29486 27636 29538
rect 27580 29428 27636 29486
rect 27692 29540 27748 29550
rect 27692 29446 27748 29484
rect 27580 29362 27636 29372
rect 27692 29316 27748 29326
rect 27692 29222 27748 29260
rect 28140 29316 28196 30156
rect 28700 29650 28756 30268
rect 29148 30322 29204 30828
rect 29148 30270 29150 30322
rect 29202 30270 29204 30322
rect 29148 30258 29204 30270
rect 29372 30100 29428 33068
rect 29484 33058 29540 33068
rect 29708 30884 29764 30894
rect 29596 30324 29652 30334
rect 29148 30044 29428 30100
rect 29484 30098 29540 30110
rect 29484 30046 29486 30098
rect 29538 30046 29540 30098
rect 28700 29598 28702 29650
rect 28754 29598 28756 29650
rect 28700 29586 28756 29598
rect 29036 29652 29092 29662
rect 28476 29540 28532 29550
rect 28476 29446 28532 29484
rect 28812 29426 28868 29438
rect 28812 29374 28814 29426
rect 28866 29374 28868 29426
rect 28812 29316 28868 29374
rect 28140 29250 28196 29260
rect 28364 29260 28868 29316
rect 26908 28914 26964 28924
rect 28364 28868 28420 29260
rect 28252 28084 28308 28094
rect 28252 27990 28308 28028
rect 26348 27748 26404 27758
rect 25900 27746 26404 27748
rect 25900 27694 26350 27746
rect 26402 27694 26404 27746
rect 25900 27692 26404 27694
rect 25788 27682 25844 27692
rect 25900 27074 25956 27086
rect 25900 27022 25902 27074
rect 25954 27022 25956 27074
rect 24668 25554 24724 25564
rect 24780 26852 24836 26862
rect 24556 25454 24558 25506
rect 24610 25454 24612 25506
rect 24556 25442 24612 25454
rect 24668 25396 24724 25406
rect 24780 25396 24836 26796
rect 24724 25340 24836 25396
rect 25004 26852 25172 26908
rect 25676 26962 25732 26974
rect 25676 26910 25678 26962
rect 25730 26910 25732 26962
rect 25676 26908 25732 26910
rect 25900 26908 25956 27022
rect 26124 27074 26180 27086
rect 26124 27022 26126 27074
rect 26178 27022 26180 27074
rect 26124 26908 26180 27022
rect 26348 27076 26404 27692
rect 26348 27010 26404 27020
rect 26796 27076 26852 27086
rect 26796 26982 26852 27020
rect 28028 27076 28084 27086
rect 28028 26982 28084 27020
rect 26460 26962 26516 26974
rect 26460 26910 26462 26962
rect 26514 26910 26516 26962
rect 25340 26852 25396 26862
rect 24668 25302 24724 25340
rect 24332 23828 24388 23838
rect 24332 23734 24388 23772
rect 23492 23324 23716 23380
rect 23436 23286 23492 23324
rect 23660 23154 23716 23324
rect 23660 23102 23662 23154
rect 23714 23102 23716 23154
rect 23660 23090 23716 23102
rect 23884 22260 23940 22270
rect 23884 22166 23940 22204
rect 23996 21588 24052 23324
rect 24332 23380 24388 23390
rect 24444 23380 24500 25228
rect 24892 23938 24948 23950
rect 24892 23886 24894 23938
rect 24946 23886 24948 23938
rect 24892 23604 24948 23886
rect 24892 23538 24948 23548
rect 24332 23378 24500 23380
rect 24332 23326 24334 23378
rect 24386 23326 24500 23378
rect 24332 23324 24500 23326
rect 24332 23314 24388 23324
rect 24108 23154 24164 23166
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 22260 24164 23102
rect 24220 23156 24276 23166
rect 24220 23062 24276 23100
rect 24444 23156 24500 23166
rect 24444 22372 24500 23100
rect 24444 22370 24612 22372
rect 24444 22318 24446 22370
rect 24498 22318 24612 22370
rect 24444 22316 24612 22318
rect 24444 22306 24500 22316
rect 24108 22194 24164 22204
rect 23996 21522 24052 21532
rect 24556 21474 24612 22316
rect 24556 21422 24558 21474
rect 24610 21422 24612 21474
rect 24556 21410 24612 21422
rect 24892 21588 24948 21598
rect 24892 20914 24948 21532
rect 24892 20862 24894 20914
rect 24946 20862 24948 20914
rect 24892 20850 24948 20862
rect 23660 19236 23716 19246
rect 23660 19142 23716 19180
rect 24332 19236 24388 19246
rect 24332 19142 24388 19180
rect 25004 19236 25060 26852
rect 25116 26516 25172 26526
rect 25116 26422 25172 26460
rect 25340 26514 25396 26796
rect 25452 26850 25508 26862
rect 25452 26798 25454 26850
rect 25506 26798 25508 26850
rect 25452 26740 25508 26798
rect 25452 26674 25508 26684
rect 25564 26850 25620 26862
rect 25676 26852 25844 26908
rect 25900 26852 26068 26908
rect 26124 26852 26404 26908
rect 25564 26798 25566 26850
rect 25618 26798 25620 26850
rect 25340 26462 25342 26514
rect 25394 26462 25396 26514
rect 25340 26450 25396 26462
rect 25452 26404 25508 26414
rect 25564 26404 25620 26798
rect 25788 26516 25844 26852
rect 26012 26628 26068 26852
rect 26012 26572 26292 26628
rect 25900 26516 25956 26526
rect 25788 26460 25900 26516
rect 25900 26450 25956 26460
rect 25452 26402 25620 26404
rect 25452 26350 25454 26402
rect 25506 26350 25620 26402
rect 25452 26348 25620 26350
rect 26236 26404 26292 26572
rect 25452 26338 25508 26348
rect 26236 26338 26292 26348
rect 26124 26292 26180 26302
rect 26124 26198 26180 26236
rect 26348 26290 26404 26852
rect 26460 26514 26516 26910
rect 26572 26852 26628 26862
rect 26572 26758 26628 26796
rect 27804 26850 27860 26862
rect 27804 26798 27806 26850
rect 27858 26798 27860 26850
rect 26460 26462 26462 26514
rect 26514 26462 26516 26514
rect 26460 26450 26516 26462
rect 27020 26516 27076 26526
rect 26348 26238 26350 26290
rect 26402 26238 26404 26290
rect 25900 26066 25956 26078
rect 25900 26014 25902 26066
rect 25954 26014 25956 26066
rect 25564 25732 25620 25742
rect 25564 25508 25620 25676
rect 25900 25732 25956 26014
rect 26124 26068 26180 26078
rect 26348 26068 26404 26238
rect 26180 26012 26292 26068
rect 26124 26002 26180 26012
rect 25900 25666 25956 25676
rect 26012 25956 26068 25966
rect 25452 25506 25620 25508
rect 25452 25454 25566 25506
rect 25618 25454 25620 25506
rect 25452 25452 25620 25454
rect 25340 24834 25396 24846
rect 25340 24782 25342 24834
rect 25394 24782 25396 24834
rect 25228 24722 25284 24734
rect 25228 24670 25230 24722
rect 25282 24670 25284 24722
rect 25228 24612 25284 24670
rect 25228 24546 25284 24556
rect 25340 24052 25396 24782
rect 25228 23996 25396 24052
rect 25228 23492 25284 23996
rect 25116 23436 25284 23492
rect 25340 23828 25396 23838
rect 25116 22260 25172 23436
rect 25340 23378 25396 23772
rect 25340 23326 25342 23378
rect 25394 23326 25396 23378
rect 25340 23314 25396 23326
rect 25228 23156 25284 23166
rect 25228 23062 25284 23100
rect 25228 22260 25284 22270
rect 25116 22204 25228 22260
rect 25228 22194 25284 22204
rect 25340 22260 25396 22270
rect 25452 22260 25508 25452
rect 25564 25442 25620 25452
rect 25900 25506 25956 25518
rect 25900 25454 25902 25506
rect 25954 25454 25956 25506
rect 25900 25396 25956 25454
rect 26012 25506 26068 25900
rect 26236 25844 26292 26012
rect 26348 26002 26404 26012
rect 26572 26292 26628 26302
rect 26572 25956 26628 26236
rect 26572 25890 26628 25900
rect 26908 26180 26964 26190
rect 26684 25844 26740 25854
rect 26236 25788 26516 25844
rect 26124 25620 26180 25630
rect 26348 25620 26404 25630
rect 26124 25526 26180 25564
rect 26236 25564 26348 25620
rect 26012 25454 26014 25506
rect 26066 25454 26068 25506
rect 26012 25442 26068 25454
rect 26236 25506 26292 25564
rect 26348 25554 26404 25564
rect 26236 25454 26238 25506
rect 26290 25454 26292 25506
rect 26236 25442 26292 25454
rect 25900 25060 25956 25340
rect 25900 25004 26180 25060
rect 25564 24948 25620 24958
rect 25564 24854 25620 24892
rect 26124 24946 26180 25004
rect 26124 24894 26126 24946
rect 26178 24894 26180 24946
rect 26124 24882 26180 24894
rect 25900 24834 25956 24846
rect 25900 24782 25902 24834
rect 25954 24782 25956 24834
rect 25788 24722 25844 24734
rect 25788 24670 25790 24722
rect 25842 24670 25844 24722
rect 25788 24612 25844 24670
rect 25788 24546 25844 24556
rect 25900 23828 25956 24782
rect 25900 23762 25956 23772
rect 26348 24500 26404 24510
rect 26348 23826 26404 24444
rect 26348 23774 26350 23826
rect 26402 23774 26404 23826
rect 25340 22258 25508 22260
rect 25340 22206 25342 22258
rect 25394 22206 25508 22258
rect 25340 22204 25508 22206
rect 25340 22194 25396 22204
rect 25340 21812 25396 21822
rect 25340 21718 25396 21756
rect 26348 21698 26404 23774
rect 26460 23940 26516 25788
rect 26684 25618 26740 25788
rect 26684 25566 26686 25618
rect 26738 25566 26740 25618
rect 26684 25554 26740 25566
rect 26908 25620 26964 26124
rect 26908 25506 26964 25564
rect 26908 25454 26910 25506
rect 26962 25454 26964 25506
rect 26908 25442 26964 25454
rect 27020 24948 27076 26460
rect 27356 26516 27412 26526
rect 27356 26422 27412 26460
rect 27804 26516 27860 26798
rect 28364 26850 28420 28812
rect 29036 28082 29092 29596
rect 29036 28030 29038 28082
rect 29090 28030 29092 28082
rect 29036 28018 29092 28030
rect 28700 27858 28756 27870
rect 28700 27806 28702 27858
rect 28754 27806 28756 27858
rect 28700 27076 28756 27806
rect 28700 27010 28756 27020
rect 29148 26908 29204 30044
rect 29484 29540 29540 30046
rect 29596 30098 29652 30268
rect 29596 30046 29598 30098
rect 29650 30046 29652 30098
rect 29596 30034 29652 30046
rect 29708 29986 29764 30828
rect 30156 30436 30212 36092
rect 30492 35924 30548 37774
rect 30716 37490 30772 39340
rect 30828 39330 30884 39340
rect 30828 39060 30884 39070
rect 30884 39004 30996 39060
rect 30828 38994 30884 39004
rect 30828 38612 30884 38622
rect 30828 38518 30884 38556
rect 30716 37438 30718 37490
rect 30770 37438 30772 37490
rect 30716 37426 30772 37438
rect 30716 36596 30772 36606
rect 30940 36596 30996 39004
rect 31276 38050 31332 38062
rect 31276 37998 31278 38050
rect 31330 37998 31332 38050
rect 31276 37492 31332 37998
rect 31276 37266 31332 37436
rect 31276 37214 31278 37266
rect 31330 37214 31332 37266
rect 31276 37202 31332 37214
rect 30716 36594 30996 36596
rect 30716 36542 30718 36594
rect 30770 36542 30996 36594
rect 30716 36540 30996 36542
rect 31052 37042 31108 37054
rect 31052 36990 31054 37042
rect 31106 36990 31108 37042
rect 30492 35868 30660 35924
rect 30492 35700 30548 35710
rect 30492 35606 30548 35644
rect 30268 34916 30324 34954
rect 30268 34850 30324 34860
rect 30268 34692 30324 34702
rect 30268 34242 30324 34636
rect 30268 34190 30270 34242
rect 30322 34190 30324 34242
rect 30268 34132 30324 34190
rect 30268 34066 30324 34076
rect 30380 34130 30436 34142
rect 30380 34078 30382 34130
rect 30434 34078 30436 34130
rect 30380 33236 30436 34078
rect 30380 33170 30436 33180
rect 30604 31668 30660 35868
rect 30716 34804 30772 36540
rect 30940 35810 30996 35822
rect 30940 35758 30942 35810
rect 30994 35758 30996 35810
rect 30940 35028 30996 35758
rect 30940 34962 30996 34972
rect 30716 34130 30772 34748
rect 31052 34804 31108 36990
rect 31164 36260 31220 36270
rect 31164 36166 31220 36204
rect 31388 35922 31444 39788
rect 31500 39618 31556 39630
rect 31500 39566 31502 39618
rect 31554 39566 31556 39618
rect 31500 37940 31556 39566
rect 31612 39396 31668 46284
rect 31948 46228 32004 46238
rect 31836 45220 31892 45230
rect 31836 45126 31892 45164
rect 31724 45106 31780 45118
rect 31724 45054 31726 45106
rect 31778 45054 31780 45106
rect 31724 44546 31780 45054
rect 31948 44994 32004 46172
rect 32060 45780 32116 46398
rect 32060 45714 32116 45724
rect 31948 44942 31950 44994
rect 32002 44942 32004 44994
rect 31948 44930 32004 44942
rect 31724 44494 31726 44546
rect 31778 44494 31780 44546
rect 31724 44482 31780 44494
rect 31836 44324 31892 44334
rect 31836 43538 31892 44268
rect 32172 44322 32228 44334
rect 32172 44270 32174 44322
rect 32226 44270 32228 44322
rect 32172 44212 32228 44270
rect 32172 43708 32228 44156
rect 31836 43486 31838 43538
rect 31890 43486 31892 43538
rect 31836 43474 31892 43486
rect 32060 43652 32228 43708
rect 32060 43538 32116 43652
rect 32060 43486 32062 43538
rect 32114 43486 32116 43538
rect 32060 43474 32116 43486
rect 32172 41972 32228 41982
rect 31612 39330 31668 39340
rect 32060 41186 32116 41198
rect 32060 41134 32062 41186
rect 32114 41134 32116 41186
rect 32060 39060 32116 41134
rect 32172 39730 32228 41916
rect 32284 41410 32340 48972
rect 32396 49026 32452 49084
rect 32732 49074 32788 49084
rect 32844 49084 32956 49140
rect 32396 48974 32398 49026
rect 32450 48974 32452 49026
rect 32396 48962 32452 48974
rect 32844 48916 32900 49084
rect 32956 49046 33012 49084
rect 32508 48860 32900 48916
rect 32508 48466 32564 48860
rect 32508 48414 32510 48466
rect 32562 48414 32564 48466
rect 32508 48402 32564 48414
rect 33068 47684 33124 54908
rect 33180 53508 33236 53518
rect 33180 53506 33348 53508
rect 33180 53454 33182 53506
rect 33234 53454 33348 53506
rect 33180 53452 33348 53454
rect 33180 53442 33236 53452
rect 33292 52500 33348 53452
rect 33180 52388 33236 52398
rect 33180 50706 33236 52332
rect 33292 52162 33348 52444
rect 33292 52110 33294 52162
rect 33346 52110 33348 52162
rect 33292 52098 33348 52110
rect 33180 50654 33182 50706
rect 33234 50654 33236 50706
rect 33180 50642 33236 50654
rect 33292 50594 33348 50606
rect 33292 50542 33294 50594
rect 33346 50542 33348 50594
rect 33292 49250 33348 50542
rect 33404 50036 33460 57820
rect 33740 57652 33796 62132
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35868 61682 35924 62300
rect 37212 62354 37268 62366
rect 37212 62302 37214 62354
rect 37266 62302 37268 62354
rect 35868 61630 35870 61682
rect 35922 61630 35924 61682
rect 35868 61618 35924 61630
rect 36764 62244 36820 62254
rect 35644 61570 35700 61582
rect 35644 61518 35646 61570
rect 35698 61518 35700 61570
rect 34412 61458 34468 61470
rect 34412 61406 34414 61458
rect 34466 61406 34468 61458
rect 34412 61124 34468 61406
rect 34972 61458 35028 61470
rect 34972 61406 34974 61458
rect 35026 61406 35028 61458
rect 34524 61346 34580 61358
rect 34524 61294 34526 61346
rect 34578 61294 34580 61346
rect 34524 61236 34580 61294
rect 34748 61348 34804 61358
rect 34748 61346 34916 61348
rect 34748 61294 34750 61346
rect 34802 61294 34916 61346
rect 34748 61292 34916 61294
rect 34748 61282 34804 61292
rect 34524 61170 34580 61180
rect 34412 61058 34468 61068
rect 33852 60900 33908 60910
rect 34748 60900 34804 60910
rect 33908 60844 34020 60900
rect 33852 60834 33908 60844
rect 33964 60452 34020 60844
rect 34748 60786 34804 60844
rect 34748 60734 34750 60786
rect 34802 60734 34804 60786
rect 34748 60722 34804 60734
rect 34076 60676 34132 60686
rect 34524 60676 34580 60686
rect 34076 60674 34580 60676
rect 34076 60622 34078 60674
rect 34130 60622 34526 60674
rect 34578 60622 34580 60674
rect 34076 60620 34580 60622
rect 34076 60610 34132 60620
rect 33964 60396 34244 60452
rect 34188 60114 34244 60396
rect 34412 60226 34468 60620
rect 34524 60610 34580 60620
rect 34412 60174 34414 60226
rect 34466 60174 34468 60226
rect 34412 60162 34468 60174
rect 34748 60564 34804 60574
rect 34748 60226 34804 60508
rect 34748 60174 34750 60226
rect 34802 60174 34804 60226
rect 34748 60162 34804 60174
rect 34188 60062 34190 60114
rect 34242 60062 34244 60114
rect 34188 60050 34244 60062
rect 34860 59220 34916 61292
rect 34972 61124 35028 61406
rect 34972 61058 35028 61068
rect 35084 61346 35140 61358
rect 35084 61294 35086 61346
rect 35138 61294 35140 61346
rect 34860 59154 34916 59164
rect 35084 58996 35140 61294
rect 35196 61346 35252 61358
rect 35196 61294 35198 61346
rect 35250 61294 35252 61346
rect 35196 61236 35252 61294
rect 35196 61170 35252 61180
rect 35420 60900 35476 60910
rect 35420 60806 35476 60844
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35644 59332 35700 61518
rect 35980 61460 36036 61470
rect 35980 61458 36260 61460
rect 35980 61406 35982 61458
rect 36034 61406 36260 61458
rect 35980 61404 36260 61406
rect 35980 61394 36036 61404
rect 36092 61236 36148 61246
rect 35868 61124 35924 61134
rect 35868 60786 35924 61068
rect 35868 60734 35870 60786
rect 35922 60734 35924 60786
rect 35868 60722 35924 60734
rect 36092 60786 36148 61180
rect 36092 60734 36094 60786
rect 36146 60734 36148 60786
rect 36092 60722 36148 60734
rect 35644 59330 36036 59332
rect 35644 59278 35646 59330
rect 35698 59278 36036 59330
rect 35644 59276 36036 59278
rect 35644 59266 35700 59276
rect 35756 58996 35812 59006
rect 35084 58994 35812 58996
rect 35084 58942 35758 58994
rect 35810 58942 35812 58994
rect 35084 58940 35812 58942
rect 35756 58930 35812 58940
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35980 58658 36036 59276
rect 36204 59220 36260 61404
rect 36764 60898 36820 62188
rect 36764 60846 36766 60898
rect 36818 60846 36820 60898
rect 36764 60834 36820 60846
rect 36988 61458 37044 61470
rect 36988 61406 36990 61458
rect 37042 61406 37044 61458
rect 36988 60564 37044 61406
rect 36988 60498 37044 60508
rect 37212 61458 37268 62302
rect 37436 61682 37492 62412
rect 37884 62466 37940 62748
rect 37884 62414 37886 62466
rect 37938 62414 37940 62466
rect 37884 62402 37940 62414
rect 38220 62468 38276 62478
rect 37436 61630 37438 61682
rect 37490 61630 37492 61682
rect 37436 61618 37492 61630
rect 37548 62242 37604 62254
rect 37548 62190 37550 62242
rect 37602 62190 37604 62242
rect 37212 61406 37214 61458
rect 37266 61406 37268 61458
rect 36540 59220 36596 59230
rect 36204 59218 36596 59220
rect 36204 59166 36542 59218
rect 36594 59166 36596 59218
rect 36204 59164 36596 59166
rect 35980 58606 35982 58658
rect 36034 58606 36036 58658
rect 35980 58594 36036 58606
rect 36316 58324 36372 58334
rect 36204 58322 36372 58324
rect 36204 58270 36318 58322
rect 36370 58270 36372 58322
rect 36204 58268 36372 58270
rect 36092 58210 36148 58222
rect 36092 58158 36094 58210
rect 36146 58158 36148 58210
rect 33740 57586 33796 57596
rect 35532 57764 35588 57774
rect 34972 57428 35028 57438
rect 33740 56980 33796 56990
rect 34972 56980 35028 57372
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 33740 56886 33796 56924
rect 34524 56978 35028 56980
rect 34524 56926 34974 56978
rect 35026 56926 35028 56978
rect 34524 56924 35028 56926
rect 34524 56866 34580 56924
rect 34972 56914 35028 56924
rect 34524 56814 34526 56866
rect 34578 56814 34580 56866
rect 34524 56802 34580 56814
rect 35196 56756 35252 56766
rect 35196 56194 35252 56700
rect 35196 56142 35198 56194
rect 35250 56142 35252 56194
rect 35196 56130 35252 56142
rect 33628 56082 33684 56094
rect 33628 56030 33630 56082
rect 33682 56030 33684 56082
rect 33628 55412 33684 56030
rect 33516 52834 33572 52846
rect 33516 52782 33518 52834
rect 33570 52782 33572 52834
rect 33516 52500 33572 52782
rect 33516 52434 33572 52444
rect 33628 52274 33684 55356
rect 34188 56082 34244 56094
rect 34188 56030 34190 56082
rect 34242 56030 34244 56082
rect 33852 55300 33908 55310
rect 34188 55300 34244 56030
rect 35532 56082 35588 57708
rect 36092 57540 36148 58158
rect 36204 57764 36260 58268
rect 36316 58258 36372 58268
rect 36428 57764 36484 57774
rect 36204 57698 36260 57708
rect 36316 57762 36484 57764
rect 36316 57710 36430 57762
rect 36482 57710 36484 57762
rect 36316 57708 36484 57710
rect 36204 57540 36260 57550
rect 36092 57538 36260 57540
rect 36092 57486 36206 57538
rect 36258 57486 36260 57538
rect 36092 57484 36260 57486
rect 35980 56866 36036 56878
rect 35980 56814 35982 56866
rect 36034 56814 36036 56866
rect 35644 56196 35700 56206
rect 35644 56102 35700 56140
rect 35532 56030 35534 56082
rect 35586 56030 35588 56082
rect 35532 56018 35588 56030
rect 35980 56084 36036 56814
rect 36092 56756 36148 56766
rect 36092 56662 36148 56700
rect 36204 56196 36260 57484
rect 36316 56978 36372 57708
rect 36428 57698 36484 57708
rect 36316 56926 36318 56978
rect 36370 56926 36372 56978
rect 36316 56914 36372 56926
rect 36428 56868 36484 56878
rect 36428 56756 36484 56812
rect 36204 56130 36260 56140
rect 36316 56754 36484 56756
rect 36316 56702 36430 56754
rect 36482 56702 36484 56754
rect 36316 56700 36484 56702
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35196 55524 35252 55534
rect 35196 55430 35252 55468
rect 35980 55524 36036 56028
rect 35980 55458 36036 55468
rect 34860 55412 34916 55422
rect 34860 55318 34916 55356
rect 34748 55300 34804 55310
rect 33852 55298 34804 55300
rect 33852 55246 33854 55298
rect 33906 55246 34750 55298
rect 34802 55246 34804 55298
rect 33852 55244 34804 55246
rect 33852 55234 33908 55244
rect 34748 55234 34804 55244
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 36316 53954 36372 56700
rect 36428 56690 36484 56700
rect 36540 56306 36596 59164
rect 37100 59220 37156 59230
rect 37100 59126 37156 59164
rect 37212 58994 37268 61406
rect 37548 61458 37604 62190
rect 38220 62244 38276 62412
rect 39452 62468 39508 62478
rect 39452 62374 39508 62412
rect 38780 62356 38836 62366
rect 38668 62354 38836 62356
rect 38668 62302 38782 62354
rect 38834 62302 38836 62354
rect 38668 62300 38836 62302
rect 38556 62244 38612 62254
rect 38220 62242 38612 62244
rect 38220 62190 38558 62242
rect 38610 62190 38612 62242
rect 38220 62188 38612 62190
rect 38220 61794 38276 62188
rect 38556 62178 38612 62188
rect 38668 62020 38724 62300
rect 38780 62290 38836 62300
rect 38220 61742 38222 61794
rect 38274 61742 38276 61794
rect 38220 61730 38276 61742
rect 38556 61964 38724 62020
rect 37548 61406 37550 61458
rect 37602 61406 37604 61458
rect 37324 61012 37380 61022
rect 37324 60918 37380 60956
rect 37548 60900 37604 61406
rect 38556 61570 38612 61964
rect 38556 61518 38558 61570
rect 38610 61518 38612 61570
rect 37548 60834 37604 60844
rect 37772 61348 37828 61358
rect 37772 60900 37828 61292
rect 38332 61348 38388 61358
rect 38332 61254 38388 61292
rect 37772 60786 37828 60844
rect 37772 60734 37774 60786
rect 37826 60734 37828 60786
rect 37772 60722 37828 60734
rect 37884 61012 37940 61022
rect 37884 60674 37940 60956
rect 37884 60622 37886 60674
rect 37938 60622 37940 60674
rect 37884 60610 37940 60622
rect 38556 60674 38612 61518
rect 38556 60622 38558 60674
rect 38610 60622 38612 60674
rect 38556 60610 38612 60622
rect 38668 61124 38724 61134
rect 38668 60788 38724 61068
rect 39116 60900 39172 60938
rect 39116 60834 39172 60844
rect 39004 60788 39060 60798
rect 38668 60786 39060 60788
rect 38668 60734 39006 60786
rect 39058 60734 39060 60786
rect 38668 60732 39060 60734
rect 37212 58942 37214 58994
rect 37266 58942 37268 58994
rect 37212 58930 37268 58942
rect 38108 60116 38164 60126
rect 37772 58548 37828 58558
rect 37660 57764 37716 57774
rect 37660 57650 37716 57708
rect 37660 57598 37662 57650
rect 37714 57598 37716 57650
rect 37660 57586 37716 57598
rect 37772 57428 37828 58492
rect 37772 57204 37828 57372
rect 37660 57148 37828 57204
rect 36540 56254 36542 56306
rect 36594 56254 36596 56306
rect 36540 56242 36596 56254
rect 36876 57092 36932 57102
rect 36316 53902 36318 53954
rect 36370 53902 36372 53954
rect 36316 53890 36372 53902
rect 36092 53842 36148 53854
rect 36092 53790 36094 53842
rect 36146 53790 36148 53842
rect 34524 53732 34580 53742
rect 34524 53638 34580 53676
rect 35980 53730 36036 53742
rect 35980 53678 35982 53730
rect 36034 53678 36036 53730
rect 35980 53172 36036 53678
rect 35980 53106 36036 53116
rect 35644 53060 35700 53070
rect 33628 52222 33630 52274
rect 33682 52222 33684 52274
rect 33628 52210 33684 52222
rect 33740 52946 33796 52958
rect 33740 52894 33742 52946
rect 33794 52894 33796 52946
rect 33740 52276 33796 52894
rect 34412 52948 34468 52958
rect 34412 52854 34468 52892
rect 35644 52946 35700 53004
rect 35644 52894 35646 52946
rect 35698 52894 35700 52946
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 33740 52050 33796 52220
rect 35644 52388 35700 52894
rect 33740 51998 33742 52050
rect 33794 51998 33796 52050
rect 33740 51986 33796 51998
rect 33852 52164 33908 52174
rect 33404 49980 33572 50036
rect 33404 49812 33460 49822
rect 33404 49718 33460 49756
rect 33292 49198 33294 49250
rect 33346 49198 33348 49250
rect 33292 49186 33348 49198
rect 32508 47628 33124 47684
rect 32508 46900 32564 47628
rect 32508 46806 32564 46844
rect 33180 45780 33236 45790
rect 33180 45686 33236 45724
rect 32508 45106 32564 45118
rect 32508 45054 32510 45106
rect 32562 45054 32564 45106
rect 32396 43764 32452 43774
rect 32508 43764 32564 45054
rect 33292 44994 33348 45006
rect 33292 44942 33294 44994
rect 33346 44942 33348 44994
rect 32620 44324 32676 44334
rect 32620 44230 32676 44268
rect 33292 44324 33348 44942
rect 33292 44258 33348 44268
rect 33068 44212 33124 44222
rect 33068 44118 33124 44156
rect 32396 43762 32564 43764
rect 32396 43710 32398 43762
rect 32450 43710 32564 43762
rect 32396 43708 32564 43710
rect 33516 43708 33572 49980
rect 33740 49698 33796 49710
rect 33740 49646 33742 49698
rect 33794 49646 33796 49698
rect 33740 49140 33796 49646
rect 33740 49046 33796 49084
rect 33628 44322 33684 44334
rect 33628 44270 33630 44322
rect 33682 44270 33684 44322
rect 33628 44212 33684 44270
rect 33628 44146 33684 44156
rect 32396 43698 32452 43708
rect 33404 43652 33572 43708
rect 33628 43988 33684 43998
rect 32620 43092 32676 43102
rect 32620 42194 32676 43036
rect 32620 42142 32622 42194
rect 32674 42142 32676 42194
rect 32620 42130 32676 42142
rect 33180 42530 33236 42542
rect 33180 42478 33182 42530
rect 33234 42478 33236 42530
rect 33180 41748 33236 42478
rect 33404 41972 33460 43652
rect 33516 43092 33572 43102
rect 33516 42866 33572 43036
rect 33516 42814 33518 42866
rect 33570 42814 33572 42866
rect 33516 42196 33572 42814
rect 33628 42420 33684 43932
rect 33852 43708 33908 52108
rect 35644 52162 35700 52332
rect 35980 52948 36036 52958
rect 35980 52274 36036 52892
rect 36092 52386 36148 53790
rect 36204 53844 36260 53854
rect 36204 53058 36260 53788
rect 36428 53732 36484 53742
rect 36204 53006 36206 53058
rect 36258 53006 36260 53058
rect 36204 52994 36260 53006
rect 36316 53172 36372 53182
rect 36092 52334 36094 52386
rect 36146 52334 36148 52386
rect 36092 52322 36148 52334
rect 35980 52222 35982 52274
rect 36034 52222 36036 52274
rect 35980 52210 36036 52222
rect 35644 52110 35646 52162
rect 35698 52110 35700 52162
rect 35644 52098 35700 52110
rect 36316 51602 36372 53116
rect 36428 53170 36484 53676
rect 36428 53118 36430 53170
rect 36482 53118 36484 53170
rect 36428 53106 36484 53118
rect 36652 53060 36708 53070
rect 36652 52966 36708 53004
rect 36764 52948 36820 52958
rect 36764 52854 36820 52892
rect 36316 51550 36318 51602
rect 36370 51550 36372 51602
rect 36316 51538 36372 51550
rect 36204 51380 36260 51390
rect 35532 51378 36260 51380
rect 35532 51326 36206 51378
rect 36258 51326 36260 51378
rect 35532 51324 36260 51326
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 50706 35252 50718
rect 35196 50654 35198 50706
rect 35250 50654 35252 50706
rect 35084 50594 35140 50606
rect 35084 50542 35086 50594
rect 35138 50542 35140 50594
rect 35084 50036 35140 50542
rect 34860 49980 35140 50036
rect 34076 49922 34132 49934
rect 34076 49870 34078 49922
rect 34130 49870 34132 49922
rect 34076 49812 34132 49870
rect 34188 49812 34244 49822
rect 34076 49756 34188 49812
rect 34188 49746 34244 49756
rect 34860 49698 34916 49980
rect 35084 49812 35140 49822
rect 35196 49812 35252 50654
rect 35420 50036 35476 50046
rect 35532 50036 35588 51324
rect 36204 51314 36260 51324
rect 36764 51378 36820 51390
rect 36764 51326 36766 51378
rect 36818 51326 36820 51378
rect 36764 51268 36820 51326
rect 35420 50034 35588 50036
rect 35420 49982 35422 50034
rect 35474 49982 35588 50034
rect 35420 49980 35588 49982
rect 36092 51156 36148 51166
rect 35420 49970 35476 49980
rect 35140 49756 35252 49812
rect 35084 49718 35140 49756
rect 34860 49646 34862 49698
rect 34914 49646 34916 49698
rect 34860 49476 34916 49646
rect 34860 49410 34916 49420
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35084 49028 35140 49038
rect 34636 47572 34692 47582
rect 34636 47478 34692 47516
rect 34972 47572 35028 47582
rect 34748 47458 34804 47470
rect 34748 47406 34750 47458
rect 34802 47406 34804 47458
rect 34748 46788 34804 47406
rect 34748 46694 34804 46732
rect 34972 46674 35028 47516
rect 34972 46622 34974 46674
rect 35026 46622 35028 46674
rect 34972 46610 35028 46622
rect 33964 45890 34020 45902
rect 33964 45838 33966 45890
rect 34018 45838 34020 45890
rect 33964 45668 34020 45838
rect 34412 45668 34468 45678
rect 33964 45666 34468 45668
rect 33964 45614 34414 45666
rect 34466 45614 34468 45666
rect 33964 45612 34468 45614
rect 34412 45332 34468 45612
rect 34412 45266 34468 45276
rect 34076 45220 34132 45230
rect 33964 44996 34020 45006
rect 33964 44098 34020 44940
rect 34076 44212 34132 45164
rect 35084 44436 35140 48972
rect 35980 48244 36036 48254
rect 35532 48242 36036 48244
rect 35532 48190 35982 48242
rect 36034 48190 36036 48242
rect 35532 48188 36036 48190
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35420 47684 35476 47694
rect 35420 47590 35476 47628
rect 35532 47236 35588 48188
rect 35980 48178 36036 48188
rect 36092 48020 36148 51100
rect 36316 50708 36372 50718
rect 36764 50708 36820 51212
rect 36316 50706 36820 50708
rect 36316 50654 36318 50706
rect 36370 50654 36820 50706
rect 36316 50652 36820 50654
rect 36316 50642 36372 50652
rect 35308 47180 35588 47236
rect 35980 47964 36148 48020
rect 36652 48130 36708 48142
rect 36652 48078 36654 48130
rect 36706 48078 36708 48130
rect 35308 46898 35364 47180
rect 35308 46846 35310 46898
rect 35362 46846 35364 46898
rect 35308 46834 35364 46846
rect 35868 46786 35924 46798
rect 35868 46734 35870 46786
rect 35922 46734 35924 46786
rect 35756 46674 35812 46686
rect 35756 46622 35758 46674
rect 35810 46622 35812 46674
rect 35756 46452 35812 46622
rect 35868 46676 35924 46734
rect 35868 46610 35924 46620
rect 35756 46386 35812 46396
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35420 44996 35476 45006
rect 35420 44902 35476 44940
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35644 44436 35700 44446
rect 35084 44380 35644 44436
rect 34300 44324 34356 44334
rect 34748 44324 34804 44334
rect 34300 44322 34804 44324
rect 34300 44270 34302 44322
rect 34354 44270 34750 44322
rect 34802 44270 34804 44322
rect 34300 44268 34804 44270
rect 34300 44258 34356 44268
rect 34748 44258 34804 44268
rect 34076 44118 34132 44156
rect 35084 44210 35140 44380
rect 35644 44342 35700 44380
rect 35084 44158 35086 44210
rect 35138 44158 35140 44210
rect 35084 44146 35140 44158
rect 33964 44046 33966 44098
rect 34018 44046 34020 44098
rect 33964 44034 34020 44046
rect 34636 44100 34692 44110
rect 34636 44006 34692 44044
rect 34860 44100 34916 44110
rect 34860 44006 34916 44044
rect 33628 42354 33684 42364
rect 33740 43652 33908 43708
rect 35084 43764 35140 43774
rect 35980 43708 36036 47964
rect 36652 47684 36708 48078
rect 36652 47618 36708 47628
rect 36428 47460 36484 47470
rect 36092 47348 36148 47358
rect 36092 46898 36148 47292
rect 36092 46846 36094 46898
rect 36146 46846 36148 46898
rect 36092 46834 36148 46846
rect 36428 46898 36484 47404
rect 36428 46846 36430 46898
rect 36482 46846 36484 46898
rect 36428 46834 36484 46846
rect 36652 46676 36708 46686
rect 36652 46582 36708 46620
rect 36316 46452 36372 46462
rect 36316 46358 36372 46396
rect 36204 45332 36260 45342
rect 36204 45106 36260 45276
rect 36652 45332 36708 45342
rect 36652 45238 36708 45276
rect 36204 45054 36206 45106
rect 36258 45054 36260 45106
rect 36204 45042 36260 45054
rect 36876 43708 36932 57036
rect 37100 56868 37156 56878
rect 37100 56196 37156 56812
rect 37324 56866 37380 56878
rect 37324 56814 37326 56866
rect 37378 56814 37380 56866
rect 37324 56756 37380 56814
rect 37324 56690 37380 56700
rect 37100 56130 37156 56140
rect 37212 56084 37268 56094
rect 37212 55990 37268 56028
rect 37660 55298 37716 57148
rect 37996 56868 38052 56878
rect 37996 56774 38052 56812
rect 37660 55246 37662 55298
rect 37714 55246 37716 55298
rect 37660 55234 37716 55246
rect 37100 53844 37156 53854
rect 37100 53750 37156 53788
rect 37996 53844 38052 53854
rect 37324 53730 37380 53742
rect 37324 53678 37326 53730
rect 37378 53678 37380 53730
rect 37324 53172 37380 53678
rect 37996 53730 38052 53788
rect 37996 53678 37998 53730
rect 38050 53678 38052 53730
rect 37996 53666 38052 53678
rect 37324 53106 37380 53116
rect 37660 52052 37716 52062
rect 37324 52050 37716 52052
rect 37324 51998 37662 52050
rect 37714 51998 37716 52050
rect 37324 51996 37716 51998
rect 37324 51490 37380 51996
rect 37660 51986 37716 51996
rect 37324 51438 37326 51490
rect 37378 51438 37380 51490
rect 37324 50428 37380 51438
rect 37996 51938 38052 51950
rect 37996 51886 37998 51938
rect 38050 51886 38052 51938
rect 37996 51378 38052 51886
rect 37996 51326 37998 51378
rect 38050 51326 38052 51378
rect 37996 51314 38052 51326
rect 37772 51268 37828 51278
rect 37772 51174 37828 51212
rect 37212 50372 37380 50428
rect 38108 50428 38164 60060
rect 38668 60114 38724 60732
rect 39004 60722 39060 60732
rect 38668 60062 38670 60114
rect 38722 60062 38724 60114
rect 38668 60050 38724 60062
rect 39452 59668 39508 59678
rect 39228 59108 39284 59118
rect 38556 58548 38612 58558
rect 38556 58434 38612 58492
rect 39228 58546 39284 59052
rect 39228 58494 39230 58546
rect 39282 58494 39284 58546
rect 39228 58482 39284 58494
rect 39452 59106 39508 59612
rect 39452 59054 39454 59106
rect 39506 59054 39508 59106
rect 38556 58382 38558 58434
rect 38610 58382 38612 58434
rect 38556 58370 38612 58382
rect 39004 57764 39060 57774
rect 39452 57764 39508 59054
rect 39004 57762 39508 57764
rect 39004 57710 39006 57762
rect 39058 57710 39508 57762
rect 39004 57708 39508 57710
rect 39004 57698 39060 57708
rect 39564 57092 39620 63868
rect 39900 61348 39956 61358
rect 39900 60786 39956 61292
rect 39900 60734 39902 60786
rect 39954 60734 39956 60786
rect 39900 60722 39956 60734
rect 40012 61010 40068 61022
rect 40012 60958 40014 61010
rect 40066 60958 40068 61010
rect 40012 60788 40068 60958
rect 40012 60722 40068 60732
rect 39900 60564 39956 60574
rect 39900 59218 39956 60508
rect 40012 59780 40068 59790
rect 40012 59686 40068 59724
rect 39900 59166 39902 59218
rect 39954 59166 39956 59218
rect 39900 59154 39956 59166
rect 39564 57036 39732 57092
rect 38220 56756 38276 56766
rect 38220 56082 38276 56700
rect 38220 56030 38222 56082
rect 38274 56030 38276 56082
rect 38220 56018 38276 56030
rect 39004 56084 39060 56094
rect 39004 55990 39060 56028
rect 38332 55188 38388 55198
rect 38332 55094 38388 55132
rect 39564 55188 39620 55198
rect 39564 54738 39620 55132
rect 39564 54686 39566 54738
rect 39618 54686 39620 54738
rect 39564 54674 39620 54686
rect 39452 54628 39508 54638
rect 39452 54534 39508 54572
rect 39564 53620 39620 53630
rect 39452 53564 39564 53620
rect 38556 53060 38612 53070
rect 38444 53004 38556 53060
rect 38444 50428 38500 53004
rect 38556 52994 38612 53004
rect 39452 52274 39508 53564
rect 39564 53526 39620 53564
rect 39452 52222 39454 52274
rect 39506 52222 39508 52274
rect 39452 52210 39508 52222
rect 38892 52164 38948 52174
rect 38668 52162 38948 52164
rect 38668 52110 38894 52162
rect 38946 52110 38948 52162
rect 38668 52108 38948 52110
rect 38668 51490 38724 52108
rect 38892 52098 38948 52108
rect 38668 51438 38670 51490
rect 38722 51438 38724 51490
rect 38668 51426 38724 51438
rect 38556 51268 38612 51278
rect 38612 51212 38724 51268
rect 38556 51202 38612 51212
rect 38556 50706 38612 50718
rect 38556 50654 38558 50706
rect 38610 50654 38612 50706
rect 38556 50428 38612 50654
rect 38108 50372 38276 50428
rect 38444 50372 38612 50428
rect 37212 49698 37268 50372
rect 37772 49924 37828 49934
rect 37772 49830 37828 49868
rect 37212 49646 37214 49698
rect 37266 49646 37268 49698
rect 37212 48354 37268 49646
rect 37212 48302 37214 48354
rect 37266 48302 37268 48354
rect 37212 48290 37268 48302
rect 37100 48242 37156 48254
rect 37100 48190 37102 48242
rect 37154 48190 37156 48242
rect 37100 47236 37156 48190
rect 37436 47684 37492 47694
rect 37436 47570 37492 47628
rect 37436 47518 37438 47570
rect 37490 47518 37492 47570
rect 37436 47506 37492 47518
rect 38108 47572 38164 47582
rect 37100 47170 37156 47180
rect 37660 47458 37716 47470
rect 37660 47406 37662 47458
rect 37714 47406 37716 47458
rect 37660 47236 37716 47406
rect 38108 47458 38164 47516
rect 38108 47406 38110 47458
rect 38162 47406 38164 47458
rect 38108 47394 38164 47406
rect 37660 47170 37716 47180
rect 37548 46900 37604 46910
rect 38220 46900 38276 50372
rect 38556 49924 38612 50372
rect 38556 49858 38612 49868
rect 38668 49810 38724 51212
rect 39340 50036 39396 50046
rect 39340 49922 39396 49980
rect 39340 49870 39342 49922
rect 39394 49870 39396 49922
rect 39340 49858 39396 49870
rect 38668 49758 38670 49810
rect 38722 49758 38724 49810
rect 38668 49746 38724 49758
rect 39676 49364 39732 57036
rect 39900 54628 39956 54638
rect 39788 54514 39844 54526
rect 39788 54462 39790 54514
rect 39842 54462 39844 54514
rect 39788 53508 39844 54462
rect 39900 53730 39956 54572
rect 40012 54514 40068 54526
rect 40012 54462 40014 54514
rect 40066 54462 40068 54514
rect 40012 53842 40068 54462
rect 40124 53956 40180 65212
rect 41356 64818 41412 64830
rect 41356 64766 41358 64818
rect 41410 64766 41412 64818
rect 41356 64708 41412 64766
rect 41692 64708 41748 64718
rect 41356 64706 41748 64708
rect 41356 64654 41694 64706
rect 41746 64654 41748 64706
rect 41356 64652 41748 64654
rect 41692 64642 41748 64652
rect 41580 64148 41636 64158
rect 41580 64054 41636 64092
rect 41244 63138 41300 63150
rect 41244 63086 41246 63138
rect 41298 63086 41300 63138
rect 41020 63028 41076 63038
rect 41020 62934 41076 62972
rect 41244 62356 41300 63086
rect 41804 63028 41860 65324
rect 42028 64148 42084 65324
rect 42700 64930 42756 65436
rect 44380 65492 44436 65502
rect 44828 65492 44884 65502
rect 44380 65490 44996 65492
rect 44380 65438 44382 65490
rect 44434 65438 44830 65490
rect 44882 65438 44996 65490
rect 44380 65436 44996 65438
rect 43708 65380 43764 65390
rect 42700 64878 42702 64930
rect 42754 64878 42756 64930
rect 42700 64866 42756 64878
rect 43596 65378 43764 65380
rect 43596 65326 43710 65378
rect 43762 65326 43764 65378
rect 43596 65324 43764 65326
rect 42028 64146 42196 64148
rect 42028 64094 42030 64146
rect 42082 64094 42196 64146
rect 42028 64092 42196 64094
rect 42028 64082 42084 64092
rect 41804 62962 41860 62972
rect 41916 62916 41972 62926
rect 41916 62466 41972 62860
rect 41916 62414 41918 62466
rect 41970 62414 41972 62466
rect 41916 62402 41972 62414
rect 41244 62262 41300 62300
rect 41020 62244 41076 62254
rect 41020 62150 41076 62188
rect 42028 61460 42084 61470
rect 41356 60788 41412 60798
rect 41356 60786 41636 60788
rect 41356 60734 41358 60786
rect 41410 60734 41636 60786
rect 41356 60732 41636 60734
rect 41356 60722 41412 60732
rect 40460 60676 40516 60686
rect 40460 59778 40516 60620
rect 41468 60564 41524 60574
rect 41468 60470 41524 60508
rect 40796 60004 40852 60014
rect 40796 60002 41524 60004
rect 40796 59950 40798 60002
rect 40850 59950 41524 60002
rect 40796 59948 41524 59950
rect 40796 59938 40852 59948
rect 40460 59726 40462 59778
rect 40514 59726 40516 59778
rect 40348 59106 40404 59118
rect 40348 59054 40350 59106
rect 40402 59054 40404 59106
rect 40348 58996 40404 59054
rect 40348 58930 40404 58940
rect 40460 57204 40516 59726
rect 40684 59778 40740 59790
rect 40908 59780 40964 59790
rect 40684 59726 40686 59778
rect 40738 59726 40740 59778
rect 40684 59556 40740 59726
rect 40684 59490 40740 59500
rect 40796 59778 40964 59780
rect 40796 59726 40910 59778
rect 40962 59726 40964 59778
rect 40796 59724 40964 59726
rect 40796 59218 40852 59724
rect 40908 59714 40964 59724
rect 41468 59330 41524 59948
rect 41468 59278 41470 59330
rect 41522 59278 41524 59330
rect 41468 59266 41524 59278
rect 40796 59166 40798 59218
rect 40850 59166 40852 59218
rect 40796 58996 40852 59166
rect 41244 59220 41300 59230
rect 41244 59126 41300 59164
rect 41020 59108 41076 59118
rect 41580 59108 41636 60732
rect 41916 60676 41972 60686
rect 41916 60582 41972 60620
rect 41804 60564 41860 60574
rect 41020 59014 41076 59052
rect 41356 59052 41636 59108
rect 41692 60002 41748 60014
rect 41692 59950 41694 60002
rect 41746 59950 41748 60002
rect 41692 59780 41748 59950
rect 40796 58930 40852 58940
rect 41020 58548 41076 58558
rect 40460 57148 40628 57204
rect 40460 55410 40516 55422
rect 40460 55358 40462 55410
rect 40514 55358 40516 55410
rect 40460 55076 40516 55358
rect 40460 55010 40516 55020
rect 40124 53890 40180 53900
rect 40012 53790 40014 53842
rect 40066 53790 40068 53842
rect 40012 53778 40068 53790
rect 39900 53678 39902 53730
rect 39954 53678 39956 53730
rect 39900 53666 39956 53678
rect 40572 53730 40628 57148
rect 40796 55186 40852 55198
rect 40796 55134 40798 55186
rect 40850 55134 40852 55186
rect 40796 54628 40852 55134
rect 40796 54562 40852 54572
rect 41020 54738 41076 58492
rect 41356 58546 41412 59052
rect 41356 58494 41358 58546
rect 41410 58494 41412 58546
rect 41356 58482 41412 58494
rect 41692 58324 41748 59724
rect 41804 59108 41860 60508
rect 41916 59668 41972 59678
rect 41916 59220 41972 59612
rect 42028 59444 42084 61404
rect 42140 60116 42196 64092
rect 43372 63924 43428 63934
rect 43372 63830 43428 63868
rect 43036 63700 43092 63710
rect 43372 63700 43428 63710
rect 43596 63700 43652 65324
rect 43708 65314 43764 65324
rect 44380 65380 44436 65436
rect 44828 65426 44884 65436
rect 44380 65314 44436 65324
rect 44940 64820 44996 65436
rect 45612 65380 45668 65390
rect 45500 65378 45668 65380
rect 45500 65326 45614 65378
rect 45666 65326 45668 65378
rect 45500 65324 45668 65326
rect 45388 64820 45444 64830
rect 44940 64818 45444 64820
rect 44940 64766 44942 64818
rect 44994 64766 45390 64818
rect 45442 64766 45444 64818
rect 44940 64764 45444 64766
rect 44940 64754 44996 64764
rect 45388 64754 45444 64764
rect 44940 64260 44996 64270
rect 44828 64036 44884 64046
rect 43036 63698 43316 63700
rect 43036 63646 43038 63698
rect 43090 63646 43316 63698
rect 43036 63644 43316 63646
rect 43036 63634 43092 63644
rect 42252 63026 42308 63038
rect 42252 62974 42254 63026
rect 42306 62974 42308 63026
rect 42252 62244 42308 62974
rect 42252 62178 42308 62188
rect 42476 62914 42532 62926
rect 42476 62862 42478 62914
rect 42530 62862 42532 62914
rect 42476 62356 42532 62862
rect 42924 62916 42980 62926
rect 42924 62822 42980 62860
rect 43260 62466 43316 63644
rect 43372 63698 43652 63700
rect 43372 63646 43374 63698
rect 43426 63646 43652 63698
rect 43372 63644 43652 63646
rect 43820 63924 43876 63934
rect 43372 63634 43428 63644
rect 43484 63140 43540 63150
rect 43484 63046 43540 63084
rect 43260 62414 43262 62466
rect 43314 62414 43316 62466
rect 43260 62402 43316 62414
rect 42700 62356 42756 62366
rect 42476 62300 42700 62356
rect 42476 62242 42532 62300
rect 42700 62290 42756 62300
rect 42812 62356 42868 62366
rect 43484 62356 43540 62366
rect 42812 62354 43204 62356
rect 42812 62302 42814 62354
rect 42866 62302 43204 62354
rect 42812 62300 43204 62302
rect 42812 62290 42868 62300
rect 42476 62190 42478 62242
rect 42530 62190 42532 62242
rect 42476 62178 42532 62190
rect 43148 62188 43204 62300
rect 43484 62262 43540 62300
rect 43596 62244 43652 62254
rect 43148 62132 43428 62188
rect 43372 61794 43428 62132
rect 43372 61742 43374 61794
rect 43426 61742 43428 61794
rect 43372 61730 43428 61742
rect 43372 61572 43428 61582
rect 43596 61572 43652 62188
rect 43372 61570 43652 61572
rect 43372 61518 43374 61570
rect 43426 61518 43652 61570
rect 43372 61516 43652 61518
rect 42700 61012 42756 61022
rect 43372 61012 43428 61516
rect 43708 61460 43764 61470
rect 43708 61366 43764 61404
rect 42700 61010 43428 61012
rect 42700 60958 42702 61010
rect 42754 60958 43428 61010
rect 42700 60956 43428 60958
rect 42700 60946 42756 60956
rect 42476 60786 42532 60798
rect 42476 60734 42478 60786
rect 42530 60734 42532 60786
rect 42476 60564 42532 60734
rect 42476 60498 42532 60508
rect 42812 60562 42868 60574
rect 42812 60510 42814 60562
rect 42866 60510 42868 60562
rect 42476 60116 42532 60126
rect 42140 60114 42532 60116
rect 42140 60062 42478 60114
rect 42530 60062 42532 60114
rect 42140 60060 42532 60062
rect 42252 59444 42308 59454
rect 42028 59442 42308 59444
rect 42028 59390 42254 59442
rect 42306 59390 42308 59442
rect 42028 59388 42308 59390
rect 42252 59378 42308 59388
rect 42364 59332 42420 59342
rect 42364 59238 42420 59276
rect 42028 59220 42084 59230
rect 41916 59218 42084 59220
rect 41916 59166 42030 59218
rect 42082 59166 42084 59218
rect 41916 59164 42084 59166
rect 42028 59154 42084 59164
rect 42140 59218 42196 59230
rect 42140 59166 42142 59218
rect 42194 59166 42196 59218
rect 41804 59052 41972 59108
rect 41916 58996 41972 59052
rect 42140 58996 42196 59166
rect 41916 58940 42196 58996
rect 41804 58548 41860 58558
rect 41804 58454 41860 58492
rect 42364 58548 42420 58558
rect 42476 58548 42532 60060
rect 42812 59668 42868 60510
rect 42812 59602 42868 59612
rect 43036 59332 43092 59342
rect 43092 59276 43204 59332
rect 43036 59238 43092 59276
rect 42420 58492 42532 58548
rect 42588 59220 42644 59230
rect 42924 59220 42980 59230
rect 42588 59218 42980 59220
rect 42588 59166 42590 59218
rect 42642 59166 42926 59218
rect 42978 59166 42980 59218
rect 42588 59164 42980 59166
rect 42364 58482 42420 58492
rect 42588 58324 42644 59164
rect 42924 59154 42980 59164
rect 43148 58658 43204 59276
rect 43260 59220 43316 59230
rect 43260 59126 43316 59164
rect 43820 59220 43876 63868
rect 44044 63140 44100 63150
rect 44044 63046 44100 63084
rect 44156 63028 44212 63038
rect 44156 62934 44212 62972
rect 44380 62916 44436 62926
rect 44380 62914 44772 62916
rect 44380 62862 44382 62914
rect 44434 62862 44772 62914
rect 44380 62860 44772 62862
rect 44380 62850 44436 62860
rect 44044 62580 44100 62590
rect 44044 62578 44660 62580
rect 44044 62526 44046 62578
rect 44098 62526 44660 62578
rect 44044 62524 44660 62526
rect 44044 62514 44100 62524
rect 43932 62356 43988 62366
rect 43932 62262 43988 62300
rect 44156 62354 44212 62366
rect 44156 62302 44158 62354
rect 44210 62302 44212 62354
rect 44156 61460 44212 62302
rect 44604 62356 44660 62524
rect 44716 62578 44772 62860
rect 44716 62526 44718 62578
rect 44770 62526 44772 62578
rect 44716 62514 44772 62526
rect 44828 62356 44884 63980
rect 44940 63140 44996 64204
rect 45164 63924 45220 63934
rect 45164 63250 45220 63868
rect 45500 63252 45556 65324
rect 45612 65314 45668 65324
rect 45164 63198 45166 63250
rect 45218 63198 45220 63250
rect 45164 63186 45220 63198
rect 45388 63196 45556 63252
rect 45612 64148 45668 64158
rect 44940 63046 44996 63084
rect 45052 63028 45108 63038
rect 45052 62934 45108 62972
rect 45276 62916 45332 62926
rect 45276 62822 45332 62860
rect 44604 62354 44884 62356
rect 44604 62302 44606 62354
rect 44658 62302 44884 62354
rect 44604 62300 44884 62302
rect 44940 62356 44996 62366
rect 44604 62290 44660 62300
rect 44940 62262 44996 62300
rect 45052 62354 45108 62366
rect 45052 62302 45054 62354
rect 45106 62302 45108 62354
rect 45052 62188 45108 62302
rect 45388 62356 45444 63196
rect 45612 63140 45668 64092
rect 45500 63084 45668 63140
rect 46060 63140 46116 63150
rect 45500 63026 45556 63084
rect 46060 63046 46116 63084
rect 45836 63028 45892 63038
rect 45500 62974 45502 63026
rect 45554 62974 45556 63026
rect 45500 62962 45556 62974
rect 45612 63026 45892 63028
rect 45612 62974 45838 63026
rect 45890 62974 45892 63026
rect 45612 62972 45892 62974
rect 45612 62804 45668 62972
rect 45500 62748 45668 62804
rect 45500 62578 45556 62748
rect 45836 62692 45892 62972
rect 46172 62804 46228 66108
rect 47404 66274 47460 66286
rect 47404 66222 47406 66274
rect 47458 66222 47460 66274
rect 46508 65380 46564 65390
rect 46508 64148 46564 65324
rect 46396 63924 46452 63934
rect 46396 63830 46452 63868
rect 46508 63140 46564 64092
rect 46732 64148 46788 64158
rect 46732 64054 46788 64092
rect 46844 64036 46900 64046
rect 46844 63942 46900 63980
rect 47068 63922 47124 63934
rect 47068 63870 47070 63922
rect 47122 63870 47124 63922
rect 46508 63138 47012 63140
rect 46508 63086 46510 63138
rect 46562 63086 47012 63138
rect 46508 63084 47012 63086
rect 46508 63074 46564 63084
rect 46172 62748 46452 62804
rect 45836 62636 46340 62692
rect 45500 62526 45502 62578
rect 45554 62526 45556 62578
rect 45500 62514 45556 62526
rect 45612 62580 45668 62590
rect 45612 62486 45668 62524
rect 45724 62356 45780 62366
rect 45948 62356 46004 62366
rect 45388 62300 45668 62356
rect 44156 61394 44212 61404
rect 44940 62132 45108 62188
rect 45612 62188 45668 62300
rect 45780 62354 46004 62356
rect 45780 62302 45950 62354
rect 46002 62302 46004 62354
rect 45780 62300 46004 62302
rect 45724 62262 45780 62300
rect 45948 62290 46004 62300
rect 46284 62354 46340 62636
rect 46284 62302 46286 62354
rect 46338 62302 46340 62354
rect 46284 62290 46340 62302
rect 46172 62244 46228 62254
rect 46060 62242 46228 62244
rect 46060 62190 46174 62242
rect 46226 62190 46228 62242
rect 46060 62188 46228 62190
rect 46396 62188 46452 62748
rect 46508 62580 46564 62590
rect 46508 62354 46564 62524
rect 46508 62302 46510 62354
rect 46562 62302 46564 62354
rect 46508 62290 46564 62302
rect 46956 62354 47012 63084
rect 47068 62692 47124 63870
rect 47292 63140 47348 63150
rect 47180 62916 47236 62926
rect 47180 62822 47236 62860
rect 47068 62636 47236 62692
rect 47180 62578 47236 62636
rect 47180 62526 47182 62578
rect 47234 62526 47236 62578
rect 47180 62514 47236 62526
rect 47292 62466 47348 63084
rect 47292 62414 47294 62466
rect 47346 62414 47348 62466
rect 47292 62402 47348 62414
rect 46956 62302 46958 62354
rect 47010 62302 47012 62354
rect 46956 62290 47012 62302
rect 47404 62188 47460 66222
rect 47516 64930 47572 67172
rect 48412 66500 48468 66510
rect 48412 66406 48468 66444
rect 49084 66500 49140 69200
rect 49084 66434 49140 66444
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 51100 65604 51156 69200
rect 52220 66500 52276 66510
rect 52220 66406 52276 66444
rect 53116 66500 53172 69200
rect 53116 66434 53172 66444
rect 51100 65538 51156 65548
rect 51212 66274 51268 66286
rect 55020 66276 55076 66286
rect 51212 66222 51214 66274
rect 51266 66222 51268 66274
rect 48860 65490 48916 65502
rect 48860 65438 48862 65490
rect 48914 65438 48916 65490
rect 47740 65380 47796 65390
rect 47740 65286 47796 65324
rect 47516 64878 47518 64930
rect 47570 64878 47572 64930
rect 47516 64866 47572 64878
rect 47516 64372 47572 64382
rect 47572 64316 47684 64372
rect 47516 64306 47572 64316
rect 45612 62132 46116 62188
rect 46172 62178 46228 62188
rect 46284 62132 46452 62188
rect 47180 62132 47460 62188
rect 44940 61346 44996 62132
rect 44940 61294 44942 61346
rect 44994 61294 44996 61346
rect 44940 60676 44996 61294
rect 44940 60610 44996 60620
rect 44268 60228 44324 60238
rect 44268 60134 44324 60172
rect 44156 59890 44212 59902
rect 44156 59838 44158 59890
rect 44210 59838 44212 59890
rect 44156 59668 44212 59838
rect 44156 59602 44212 59612
rect 43820 59154 43876 59164
rect 45276 59220 45332 59258
rect 45332 59164 45444 59220
rect 45276 59154 45332 59164
rect 45388 59108 45444 59164
rect 45724 59108 45780 59118
rect 45388 59106 45780 59108
rect 45388 59054 45726 59106
rect 45778 59054 45780 59106
rect 45388 59052 45780 59054
rect 44940 58994 44996 59006
rect 44940 58942 44942 58994
rect 44994 58942 44996 58994
rect 43148 58606 43150 58658
rect 43202 58606 43204 58658
rect 43148 58594 43204 58606
rect 43260 58772 43316 58782
rect 41692 58258 41748 58268
rect 42476 58268 42644 58324
rect 43148 58436 43204 58446
rect 43148 58322 43204 58380
rect 43260 58436 43316 58716
rect 44828 58546 44884 58558
rect 44828 58494 44830 58546
rect 44882 58494 44884 58546
rect 44828 58436 44884 58494
rect 43260 58434 43428 58436
rect 43260 58382 43262 58434
rect 43314 58382 43428 58434
rect 43260 58380 43428 58382
rect 43260 58370 43316 58380
rect 43148 58270 43150 58322
rect 43202 58270 43204 58322
rect 42140 57650 42196 57662
rect 42140 57598 42142 57650
rect 42194 57598 42196 57650
rect 42140 56868 42196 57598
rect 42364 56980 42420 56990
rect 42476 56980 42532 58268
rect 43148 57764 43204 58270
rect 43260 57764 43316 57774
rect 42700 57762 43316 57764
rect 42700 57710 43262 57762
rect 43314 57710 43316 57762
rect 42700 57708 43316 57710
rect 42588 57540 42644 57550
rect 42588 57446 42644 57484
rect 42700 57204 42756 57708
rect 43260 57698 43316 57708
rect 43148 57540 43204 57550
rect 43372 57540 43428 58380
rect 44828 58370 44884 58380
rect 44940 57874 44996 58942
rect 45276 58994 45332 59006
rect 45276 58942 45278 58994
rect 45330 58942 45332 58994
rect 45276 58548 45332 58942
rect 45724 58884 45780 59052
rect 45724 58818 45780 58828
rect 45276 58482 45332 58492
rect 44940 57822 44942 57874
rect 44994 57822 44996 57874
rect 44940 57810 44996 57822
rect 43204 57484 43428 57540
rect 43596 57652 43652 57662
rect 43148 57446 43204 57484
rect 42364 56978 42532 56980
rect 42364 56926 42366 56978
rect 42418 56926 42532 56978
rect 42364 56924 42532 56926
rect 42588 57148 42756 57204
rect 42364 56914 42420 56924
rect 42252 56868 42308 56878
rect 42140 56812 42252 56868
rect 42252 56774 42308 56812
rect 42476 56756 42532 56766
rect 42588 56756 42644 57148
rect 42700 57036 43540 57092
rect 42700 56978 42756 57036
rect 42700 56926 42702 56978
rect 42754 56926 42756 56978
rect 42700 56914 42756 56926
rect 42476 56754 42644 56756
rect 42476 56702 42478 56754
rect 42530 56702 42644 56754
rect 42476 56700 42644 56702
rect 42924 56866 42980 56878
rect 42924 56814 42926 56866
rect 42978 56814 42980 56866
rect 42924 56756 42980 56814
rect 42476 56690 42532 56700
rect 41692 55972 41748 55982
rect 41580 55412 41636 55422
rect 41580 55318 41636 55356
rect 41468 55298 41524 55310
rect 41468 55246 41470 55298
rect 41522 55246 41524 55298
rect 41468 55076 41524 55246
rect 41468 55010 41524 55020
rect 41580 54740 41636 54750
rect 41020 54686 41022 54738
rect 41074 54686 41076 54738
rect 41020 54068 41076 54686
rect 41020 54002 41076 54012
rect 41244 54738 41636 54740
rect 41244 54686 41582 54738
rect 41634 54686 41636 54738
rect 41244 54684 41636 54686
rect 40572 53678 40574 53730
rect 40626 53678 40628 53730
rect 40124 53508 40180 53518
rect 39788 53452 40124 53508
rect 40124 53414 40180 53452
rect 39676 49298 39732 49308
rect 40572 52724 40628 53678
rect 41244 53732 41300 54684
rect 41580 54674 41636 54684
rect 41692 54738 41748 55916
rect 42924 55972 42980 56700
rect 42924 55906 42980 55916
rect 43148 55522 43204 57036
rect 43260 56756 43316 56766
rect 43260 56662 43316 56700
rect 43484 56754 43540 57036
rect 43596 57090 43652 57596
rect 44492 57652 44548 57662
rect 44492 57558 44548 57596
rect 43596 57038 43598 57090
rect 43650 57038 43652 57090
rect 43596 57026 43652 57038
rect 43484 56702 43486 56754
rect 43538 56702 43540 56754
rect 43484 56690 43540 56702
rect 45500 55972 45556 55982
rect 45500 55878 45556 55916
rect 43148 55470 43150 55522
rect 43202 55470 43204 55522
rect 43148 55458 43204 55470
rect 45612 55858 45668 55870
rect 45612 55806 45614 55858
rect 45666 55806 45668 55858
rect 42140 55412 42196 55422
rect 42140 55318 42196 55356
rect 45612 55410 45668 55806
rect 45612 55358 45614 55410
rect 45666 55358 45668 55410
rect 45612 55346 45668 55358
rect 42364 55300 42420 55310
rect 42812 55300 42868 55310
rect 42252 55298 42868 55300
rect 42252 55246 42366 55298
rect 42418 55246 42814 55298
rect 42866 55246 42868 55298
rect 42252 55244 42868 55246
rect 41692 54686 41694 54738
rect 41746 54686 41748 54738
rect 41692 54674 41748 54686
rect 41804 54740 41860 54750
rect 41804 54646 41860 54684
rect 41468 54514 41524 54526
rect 41468 54462 41470 54514
rect 41522 54462 41524 54514
rect 41468 54068 41524 54462
rect 42028 54516 42084 54526
rect 42252 54516 42308 55244
rect 42364 55234 42420 55244
rect 42812 55234 42868 55244
rect 44268 55300 44324 55310
rect 42364 55076 42420 55086
rect 42364 54626 42420 55020
rect 43036 55074 43092 55086
rect 43036 55022 43038 55074
rect 43090 55022 43092 55074
rect 43036 54852 43092 55022
rect 42476 54796 43092 54852
rect 44268 55074 44324 55244
rect 44940 55300 44996 55310
rect 44940 55206 44996 55244
rect 46284 55076 46340 62132
rect 47068 60002 47124 60014
rect 47068 59950 47070 60002
rect 47122 59950 47124 60002
rect 47068 59444 47124 59950
rect 47068 59378 47124 59388
rect 46956 58548 47012 58558
rect 46956 58454 47012 58492
rect 47068 57428 47124 57438
rect 47068 56978 47124 57372
rect 47068 56926 47070 56978
rect 47122 56926 47124 56978
rect 47068 56914 47124 56926
rect 46956 56308 47012 56318
rect 47180 56308 47236 62132
rect 46732 56306 47236 56308
rect 46732 56254 46958 56306
rect 47010 56254 47236 56306
rect 46732 56252 47236 56254
rect 47628 56308 47684 64316
rect 47740 63588 47796 63598
rect 47740 63250 47796 63532
rect 47740 63198 47742 63250
rect 47794 63198 47796 63250
rect 47740 63140 47796 63198
rect 47740 63074 47796 63084
rect 48860 62580 48916 65438
rect 49532 65380 49588 65390
rect 49532 65378 50260 65380
rect 49532 65326 49534 65378
rect 49586 65326 50260 65378
rect 49532 65324 50260 65326
rect 49532 65314 49588 65324
rect 50204 64930 50260 65324
rect 50204 64878 50206 64930
rect 50258 64878 50260 64930
rect 50204 64866 50260 64878
rect 48860 62354 48916 62524
rect 49420 64706 49476 64718
rect 49420 64654 49422 64706
rect 49474 64654 49476 64706
rect 49420 62356 49476 64654
rect 50316 64594 50372 64606
rect 50316 64542 50318 64594
rect 50370 64542 50372 64594
rect 49532 64260 49588 64270
rect 49532 63924 49588 64204
rect 50316 64148 50372 64542
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 51212 64260 51268 66222
rect 54460 66274 55076 66276
rect 54460 66222 55022 66274
rect 55074 66222 55076 66274
rect 54460 66220 55076 66222
rect 52332 65492 52388 65502
rect 51660 65380 51716 65390
rect 50556 64250 50820 64260
rect 50988 64204 51268 64260
rect 51324 65378 51716 65380
rect 51324 65326 51662 65378
rect 51714 65326 51716 65378
rect 51324 65324 51716 65326
rect 50428 64148 50484 64158
rect 50316 64146 50484 64148
rect 50316 64094 50430 64146
rect 50482 64094 50484 64146
rect 50316 64092 50484 64094
rect 50428 64082 50484 64092
rect 50876 64036 50932 64046
rect 50764 64034 50932 64036
rect 50764 63982 50878 64034
rect 50930 63982 50932 64034
rect 50764 63980 50932 63982
rect 49532 63830 49588 63868
rect 49644 63922 49700 63934
rect 49644 63870 49646 63922
rect 49698 63870 49700 63922
rect 49644 63140 49700 63870
rect 49980 63922 50036 63934
rect 49980 63870 49982 63922
rect 50034 63870 50036 63922
rect 49980 63252 50036 63870
rect 49980 63186 50036 63196
rect 50092 63922 50148 63934
rect 50092 63870 50094 63922
rect 50146 63870 50148 63922
rect 49644 63074 49700 63084
rect 48860 62302 48862 62354
rect 48914 62302 48916 62354
rect 48860 62290 48916 62302
rect 49084 62300 49476 62356
rect 49084 62188 49140 62300
rect 49532 62244 49588 62254
rect 48972 62132 49140 62188
rect 49196 62242 49588 62244
rect 49196 62190 49534 62242
rect 49586 62190 49588 62242
rect 49196 62188 49588 62190
rect 48860 61908 48916 61918
rect 48860 60786 48916 61852
rect 48860 60734 48862 60786
rect 48914 60734 48916 60786
rect 48860 60228 48916 60734
rect 48860 60162 48916 60172
rect 47740 59892 47796 59902
rect 47740 59890 48132 59892
rect 47740 59838 47742 59890
rect 47794 59838 48132 59890
rect 47740 59836 48132 59838
rect 47740 59826 47796 59836
rect 48076 59442 48132 59836
rect 48972 59668 49028 62132
rect 49196 61794 49252 62188
rect 49532 62178 49588 62188
rect 50092 62244 50148 63870
rect 49196 61742 49198 61794
rect 49250 61742 49252 61794
rect 49196 61730 49252 61742
rect 49084 61460 49140 61470
rect 49084 61458 49476 61460
rect 49084 61406 49086 61458
rect 49138 61406 49476 61458
rect 49084 61404 49476 61406
rect 49084 61394 49140 61404
rect 49420 61124 49476 61404
rect 49420 61068 49700 61124
rect 48860 59612 49028 59668
rect 49084 61012 49140 61022
rect 48076 59390 48078 59442
rect 48130 59390 48132 59442
rect 48076 59378 48132 59390
rect 48300 59444 48356 59454
rect 48188 59332 48244 59342
rect 48188 59238 48244 59276
rect 48188 58548 48244 58558
rect 48300 58548 48356 59388
rect 48860 59442 48916 59612
rect 48860 59390 48862 59442
rect 48914 59390 48916 59442
rect 48860 58772 48916 59390
rect 48972 59444 49028 59454
rect 49084 59444 49140 60956
rect 49644 61010 49700 61068
rect 49644 60958 49646 61010
rect 49698 60958 49700 61010
rect 49644 60946 49700 60958
rect 49756 61012 49812 61022
rect 48972 59442 49140 59444
rect 48972 59390 48974 59442
rect 49026 59390 49140 59442
rect 48972 59388 49140 59390
rect 49308 60786 49364 60798
rect 49308 60734 49310 60786
rect 49362 60734 49364 60786
rect 48972 59378 49028 59388
rect 48860 58706 48916 58716
rect 49308 59218 49364 60734
rect 49644 60786 49700 60798
rect 49644 60734 49646 60786
rect 49698 60734 49700 60786
rect 49532 60676 49588 60686
rect 49532 60004 49588 60620
rect 49644 60228 49700 60734
rect 49756 60676 49812 60956
rect 50092 60786 50148 62188
rect 50428 63810 50484 63822
rect 50428 63758 50430 63810
rect 50482 63758 50484 63810
rect 50428 61012 50484 63758
rect 50764 63810 50820 63980
rect 50876 63970 50932 63980
rect 50764 63758 50766 63810
rect 50818 63758 50820 63810
rect 50764 63746 50820 63758
rect 50652 63588 50708 63598
rect 50652 63138 50708 63532
rect 50652 63086 50654 63138
rect 50706 63086 50708 63138
rect 50652 63074 50708 63086
rect 50764 63140 50820 63150
rect 50764 63046 50820 63084
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 50988 61908 51044 64204
rect 51324 64148 51380 65324
rect 51660 65314 51716 65324
rect 51772 65380 51828 65390
rect 51772 64930 51828 65324
rect 51772 64878 51774 64930
rect 51826 64878 51828 64930
rect 51772 64866 51828 64878
rect 51996 65378 52052 65390
rect 51996 65326 51998 65378
rect 52050 65326 52052 65378
rect 51212 64092 51380 64148
rect 51660 64594 51716 64606
rect 51660 64542 51662 64594
rect 51714 64542 51716 64594
rect 51212 64034 51268 64092
rect 51212 63982 51214 64034
rect 51266 63982 51268 64034
rect 50988 61842 51044 61852
rect 51100 63252 51156 63262
rect 51100 63138 51156 63196
rect 51100 63086 51102 63138
rect 51154 63086 51156 63138
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50428 60946 50484 60956
rect 50988 61012 51044 61022
rect 50988 60918 51044 60956
rect 50092 60734 50094 60786
rect 50146 60734 50148 60786
rect 50092 60722 50148 60734
rect 50204 60900 50260 60910
rect 49756 60582 49812 60620
rect 49644 60172 49924 60228
rect 49868 60114 49924 60172
rect 49868 60062 49870 60114
rect 49922 60062 49924 60114
rect 49532 59948 49700 60004
rect 49532 59442 49588 59454
rect 49532 59390 49534 59442
rect 49586 59390 49588 59442
rect 49532 59332 49588 59390
rect 49532 59266 49588 59276
rect 49308 59166 49310 59218
rect 49362 59166 49364 59218
rect 47740 58546 48356 58548
rect 47740 58494 48190 58546
rect 48242 58494 48356 58546
rect 47740 58492 48356 58494
rect 47740 58434 47796 58492
rect 48188 58482 48244 58492
rect 47740 58382 47742 58434
rect 47794 58382 47796 58434
rect 47740 58370 47796 58382
rect 48188 57428 48244 57438
rect 48076 57372 48188 57428
rect 46396 55972 46452 55982
rect 46452 55916 46676 55972
rect 46396 55906 46452 55916
rect 44268 55022 44270 55074
rect 44322 55022 44324 55074
rect 42476 54740 42532 54796
rect 42476 54646 42532 54684
rect 42364 54574 42366 54626
rect 42418 54574 42420 54626
rect 42364 54562 42420 54574
rect 42028 54514 42308 54516
rect 42028 54462 42030 54514
rect 42082 54462 42308 54514
rect 42028 54460 42308 54462
rect 41468 54012 41860 54068
rect 41244 53676 41524 53732
rect 40908 53620 40964 53630
rect 40908 53526 40964 53564
rect 41244 53618 41300 53676
rect 41244 53566 41246 53618
rect 41298 53566 41300 53618
rect 41244 53554 41300 53566
rect 41468 53620 41524 53676
rect 41580 53620 41636 53630
rect 41468 53618 41636 53620
rect 41468 53566 41582 53618
rect 41634 53566 41636 53618
rect 41468 53564 41636 53566
rect 41580 53554 41636 53564
rect 41692 53620 41748 53630
rect 41804 53620 41860 54012
rect 42028 53844 42084 54460
rect 42028 53778 42084 53788
rect 42476 54068 42532 54078
rect 41692 53618 41860 53620
rect 41692 53566 41694 53618
rect 41746 53566 41860 53618
rect 41692 53564 41860 53566
rect 41020 53506 41076 53518
rect 41020 53454 41022 53506
rect 41074 53454 41076 53506
rect 41020 53060 41076 53454
rect 41356 53508 41412 53518
rect 41356 53414 41412 53452
rect 41020 52994 41076 53004
rect 41020 52834 41076 52846
rect 41020 52782 41022 52834
rect 41074 52782 41076 52834
rect 41020 52724 41076 52782
rect 40572 52668 41076 52724
rect 38444 47460 38500 47470
rect 38444 47366 38500 47404
rect 39004 47458 39060 47470
rect 39004 47406 39006 47458
rect 39058 47406 39060 47458
rect 39004 47348 39060 47406
rect 39004 47282 39060 47292
rect 39116 47346 39172 47358
rect 39116 47294 39118 47346
rect 39170 47294 39172 47346
rect 38556 47236 38612 47246
rect 38556 47142 38612 47180
rect 38332 46900 38388 46910
rect 38220 46844 38332 46900
rect 37436 46786 37492 46798
rect 37436 46734 37438 46786
rect 37490 46734 37492 46786
rect 37436 46676 37492 46734
rect 37100 46562 37156 46574
rect 37100 46510 37102 46562
rect 37154 46510 37156 46562
rect 37100 46452 37156 46510
rect 37100 46386 37156 46396
rect 33628 42196 33684 42206
rect 33516 42140 33628 42196
rect 33628 42102 33684 42140
rect 33740 42084 33796 43652
rect 33740 42018 33796 42028
rect 33852 43540 33908 43550
rect 33404 41916 33572 41972
rect 33404 41748 33460 41758
rect 33180 41692 33404 41748
rect 33404 41654 33460 41692
rect 32284 41358 32286 41410
rect 32338 41358 32340 41410
rect 32284 41346 32340 41358
rect 32508 41300 32564 41310
rect 32508 39732 32564 41244
rect 33180 41188 33236 41198
rect 33180 41094 33236 41132
rect 32172 39678 32174 39730
rect 32226 39678 32228 39730
rect 32172 39666 32228 39678
rect 32284 39730 32564 39732
rect 32284 39678 32510 39730
rect 32562 39678 32564 39730
rect 32284 39676 32564 39678
rect 32060 38994 32116 39004
rect 31500 37156 31556 37884
rect 31836 38780 32228 38836
rect 31836 37938 31892 38780
rect 32172 38724 32228 38780
rect 32284 38724 32340 39676
rect 32508 39666 32564 39676
rect 33068 39394 33124 39406
rect 33068 39342 33070 39394
rect 33122 39342 33124 39394
rect 32172 38722 32340 38724
rect 32172 38670 32174 38722
rect 32226 38670 32340 38722
rect 32172 38668 32340 38670
rect 32508 38834 32564 38846
rect 32508 38782 32510 38834
rect 32562 38782 32564 38834
rect 32508 38668 32564 38782
rect 32172 38658 32228 38668
rect 31836 37886 31838 37938
rect 31890 37886 31892 37938
rect 31836 37874 31892 37886
rect 31948 38610 32004 38622
rect 32508 38612 33012 38668
rect 31948 38558 31950 38610
rect 32002 38558 32004 38610
rect 31948 38500 32004 38558
rect 31500 37090 31556 37100
rect 31388 35870 31390 35922
rect 31442 35870 31444 35922
rect 31388 35858 31444 35870
rect 31388 35698 31444 35710
rect 31388 35646 31390 35698
rect 31442 35646 31444 35698
rect 31052 34738 31108 34748
rect 31164 35588 31220 35598
rect 30716 34078 30718 34130
rect 30770 34078 30772 34130
rect 30716 34066 30772 34078
rect 30940 34242 30996 34254
rect 30940 34190 30942 34242
rect 30994 34190 30996 34242
rect 30940 34132 30996 34190
rect 30940 33122 30996 34076
rect 30940 33070 30942 33122
rect 30994 33070 30996 33122
rect 30828 31892 30884 31902
rect 30828 31798 30884 31836
rect 30604 31602 30660 31612
rect 30940 31444 30996 33070
rect 30380 31388 30996 31444
rect 31164 31778 31220 35532
rect 31388 34242 31444 35646
rect 31388 34190 31390 34242
rect 31442 34190 31444 34242
rect 31388 34178 31444 34190
rect 31500 35252 31556 35262
rect 31276 33122 31332 33134
rect 31276 33070 31278 33122
rect 31330 33070 31332 33122
rect 31276 31892 31332 33070
rect 31500 33122 31556 35196
rect 31612 35028 31668 35038
rect 31612 34018 31668 34972
rect 31836 34132 31892 34142
rect 31836 34038 31892 34076
rect 31612 33966 31614 34018
rect 31666 33966 31668 34018
rect 31612 33954 31668 33966
rect 31836 33908 31892 33918
rect 31836 33346 31892 33852
rect 31836 33294 31838 33346
rect 31890 33294 31892 33346
rect 31836 33282 31892 33294
rect 31500 33070 31502 33122
rect 31554 33070 31556 33122
rect 31500 33058 31556 33070
rect 31836 32676 31892 32686
rect 31276 31826 31332 31836
rect 31612 32562 31668 32574
rect 31612 32510 31614 32562
rect 31666 32510 31668 32562
rect 31164 31726 31166 31778
rect 31218 31726 31220 31778
rect 30156 30380 30324 30436
rect 30044 30324 30100 30334
rect 30044 30212 30100 30268
rect 30156 30212 30212 30222
rect 30044 30210 30212 30212
rect 30044 30158 30158 30210
rect 30210 30158 30212 30210
rect 30044 30156 30212 30158
rect 30156 30146 30212 30156
rect 29708 29934 29710 29986
rect 29762 29934 29764 29986
rect 29708 29540 29764 29934
rect 29932 29986 29988 29998
rect 30268 29988 30324 30380
rect 30380 30098 30436 31388
rect 31052 31220 31108 31230
rect 31164 31220 31220 31726
rect 31052 31218 31220 31220
rect 31052 31166 31054 31218
rect 31106 31166 31220 31218
rect 31052 31164 31220 31166
rect 31052 31154 31108 31164
rect 31276 30212 31332 30222
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 30380 30034 30436 30046
rect 30492 30100 30548 30110
rect 29932 29934 29934 29986
rect 29986 29934 29988 29986
rect 29932 29652 29988 29934
rect 29932 29586 29988 29596
rect 30044 29932 30324 29988
rect 29484 29474 29540 29484
rect 29596 29484 29764 29540
rect 29260 29316 29316 29326
rect 29596 29316 29652 29484
rect 29260 29314 29652 29316
rect 29260 29262 29262 29314
rect 29314 29262 29652 29314
rect 29260 29260 29652 29262
rect 29708 29316 29764 29326
rect 29260 29250 29316 29260
rect 29708 28644 29764 29260
rect 29708 28578 29764 28588
rect 30044 28420 30100 29932
rect 30492 28868 30548 30044
rect 31164 30100 31220 30110
rect 31164 30006 31220 30044
rect 31276 30098 31332 30156
rect 31276 30046 31278 30098
rect 31330 30046 31332 30098
rect 31276 30034 31332 30046
rect 31500 29988 31556 29998
rect 31388 29986 31556 29988
rect 31388 29934 31502 29986
rect 31554 29934 31556 29986
rect 31388 29932 31556 29934
rect 31388 29764 31444 29932
rect 31500 29922 31556 29932
rect 31164 29708 31444 29764
rect 30604 29652 30660 29662
rect 30660 29596 30772 29652
rect 30604 29586 30660 29596
rect 30716 29540 30772 29596
rect 30716 29538 30884 29540
rect 30716 29486 30718 29538
rect 30770 29486 30884 29538
rect 30716 29484 30884 29486
rect 30716 29474 30772 29484
rect 30716 29092 30772 29102
rect 30604 28868 30660 28878
rect 30492 28812 30604 28868
rect 30380 28756 30436 28766
rect 30268 28644 30324 28654
rect 30268 28550 30324 28588
rect 28364 26798 28366 26850
rect 28418 26798 28420 26850
rect 28364 26786 28420 26798
rect 28924 26852 29204 26908
rect 29372 28364 30100 28420
rect 29372 27186 29428 28364
rect 30380 27972 30436 28700
rect 30604 28642 30660 28812
rect 30604 28590 30606 28642
rect 30658 28590 30660 28642
rect 30604 28578 30660 28590
rect 30716 28530 30772 29036
rect 30716 28478 30718 28530
rect 30770 28478 30772 28530
rect 30716 28466 30772 28478
rect 30828 28082 30884 29484
rect 30940 29538 30996 29550
rect 30940 29486 30942 29538
rect 30994 29486 30996 29538
rect 30940 29316 30996 29486
rect 31164 29426 31220 29708
rect 31612 29652 31668 32510
rect 31836 32562 31892 32620
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32498 31892 32510
rect 31948 30322 32004 38444
rect 32956 38050 33012 38612
rect 32956 37998 32958 38050
rect 33010 37998 33012 38050
rect 32620 37044 32676 37054
rect 32060 36370 32116 36382
rect 32060 36318 32062 36370
rect 32114 36318 32116 36370
rect 32060 36260 32116 36318
rect 32060 32786 32116 36204
rect 32396 35812 32452 35822
rect 32284 35810 32452 35812
rect 32284 35758 32398 35810
rect 32450 35758 32452 35810
rect 32284 35756 32452 35758
rect 32060 32734 32062 32786
rect 32114 32734 32116 32786
rect 32060 32722 32116 32734
rect 32172 32788 32228 32798
rect 32172 32450 32228 32732
rect 32172 32398 32174 32450
rect 32226 32398 32228 32450
rect 32172 32386 32228 32398
rect 32284 32676 32340 35756
rect 32396 35746 32452 35756
rect 32508 35700 32564 35710
rect 32620 35700 32676 36988
rect 32956 36258 33012 37998
rect 33068 37828 33124 39342
rect 33068 37762 33124 37772
rect 33068 37268 33124 37278
rect 33068 36932 33124 37212
rect 33404 37268 33460 37278
rect 33404 37174 33460 37212
rect 33404 36932 33460 36942
rect 33068 36876 33404 36932
rect 33068 36482 33124 36876
rect 33404 36866 33460 36876
rect 33292 36596 33348 36606
rect 33292 36502 33348 36540
rect 33068 36430 33070 36482
rect 33122 36430 33124 36482
rect 33068 36418 33124 36430
rect 32956 36206 32958 36258
rect 33010 36206 33012 36258
rect 32956 36194 33012 36206
rect 32508 35698 32676 35700
rect 32508 35646 32510 35698
rect 32562 35646 32676 35698
rect 32508 35644 32676 35646
rect 32508 35634 32564 35644
rect 32396 35474 32452 35486
rect 32396 35422 32398 35474
rect 32450 35422 32452 35474
rect 32396 33234 32452 35422
rect 32396 33182 32398 33234
rect 32450 33182 32452 33234
rect 32396 33170 32452 33182
rect 32284 32116 32340 32620
rect 32284 32050 32340 32060
rect 31948 30270 31950 30322
rect 32002 30270 32004 30322
rect 31948 30258 32004 30270
rect 32508 31892 32564 31902
rect 32508 30322 32564 31836
rect 32620 31890 32676 35644
rect 33292 35364 33348 35374
rect 32620 31838 32622 31890
rect 32674 31838 32676 31890
rect 32620 31826 32676 31838
rect 33180 32788 33236 32798
rect 32956 31780 33012 31790
rect 32956 31686 33012 31724
rect 32508 30270 32510 30322
rect 32562 30270 32564 30322
rect 32508 30258 32564 30270
rect 33180 30100 33236 32732
rect 33292 31778 33348 35308
rect 33292 31726 33294 31778
rect 33346 31726 33348 31778
rect 33292 31714 33348 31726
rect 33292 30100 33348 30110
rect 33180 30098 33348 30100
rect 33180 30046 33294 30098
rect 33346 30046 33348 30098
rect 33180 30044 33348 30046
rect 33292 30034 33348 30044
rect 31388 29596 31612 29652
rect 31276 29540 31332 29550
rect 31276 29446 31332 29484
rect 31164 29374 31166 29426
rect 31218 29374 31220 29426
rect 31164 29362 31220 29374
rect 30940 29250 30996 29260
rect 31388 29092 31444 29596
rect 31612 29558 31668 29596
rect 31500 29316 31556 29326
rect 31948 29316 32004 29326
rect 31500 29314 31892 29316
rect 31500 29262 31502 29314
rect 31554 29262 31892 29314
rect 31500 29260 31892 29262
rect 31500 29250 31556 29260
rect 31388 29026 31444 29036
rect 31052 28812 31332 28868
rect 30940 28644 30996 28654
rect 31052 28644 31108 28812
rect 30940 28642 31108 28644
rect 30940 28590 30942 28642
rect 30994 28590 31108 28642
rect 30940 28588 31108 28590
rect 31164 28644 31220 28654
rect 30940 28578 30996 28588
rect 31164 28196 31220 28588
rect 30828 28030 30830 28082
rect 30882 28030 30884 28082
rect 30828 28018 30884 28030
rect 30940 28140 31220 28196
rect 30380 27906 30436 27916
rect 29372 27134 29374 27186
rect 29426 27134 29428 27186
rect 27804 26450 27860 26460
rect 28476 26516 28532 26526
rect 28476 26422 28532 26460
rect 27468 26404 27524 26414
rect 27132 26290 27188 26302
rect 27132 26238 27134 26290
rect 27186 26238 27188 26290
rect 27132 25396 27188 26238
rect 27468 26290 27524 26348
rect 28812 26404 28868 26414
rect 28812 26310 28868 26348
rect 27468 26238 27470 26290
rect 27522 26238 27524 26290
rect 27468 26226 27524 26238
rect 28252 26292 28308 26302
rect 28252 26198 28308 26236
rect 28588 26292 28644 26302
rect 27244 26178 27300 26190
rect 27244 26126 27246 26178
rect 27298 26126 27300 26178
rect 27244 25508 27300 26126
rect 27804 26066 27860 26078
rect 27804 26014 27806 26066
rect 27858 26014 27860 26066
rect 27804 25732 27860 26014
rect 27804 25666 27860 25676
rect 27692 25620 27748 25630
rect 27692 25526 27748 25564
rect 27916 25620 27972 25630
rect 27244 25442 27300 25452
rect 27804 25508 27860 25518
rect 27916 25508 27972 25564
rect 28588 25620 28644 26236
rect 28588 25526 28644 25564
rect 27804 25506 28196 25508
rect 27804 25454 27806 25506
rect 27858 25454 28196 25506
rect 27804 25452 28196 25454
rect 27132 25330 27188 25340
rect 27356 25394 27412 25406
rect 27356 25342 27358 25394
rect 27410 25342 27412 25394
rect 27132 24948 27188 24958
rect 27020 24946 27188 24948
rect 27020 24894 27134 24946
rect 27186 24894 27188 24946
rect 27020 24892 27188 24894
rect 27020 24500 27076 24892
rect 27132 24882 27188 24892
rect 27356 24948 27412 25342
rect 27804 25284 27860 25452
rect 27356 24882 27412 24892
rect 27468 25228 27860 25284
rect 28028 25284 28084 25294
rect 27468 24724 27524 25228
rect 27692 24948 27748 24958
rect 27692 24836 27748 24892
rect 27692 24834 27972 24836
rect 27692 24782 27694 24834
rect 27746 24782 27972 24834
rect 27692 24780 27972 24782
rect 27692 24770 27748 24780
rect 27468 24722 27636 24724
rect 27468 24670 27470 24722
rect 27522 24670 27636 24722
rect 27468 24668 27636 24670
rect 27468 24658 27524 24668
rect 27020 24434 27076 24444
rect 27580 24052 27636 24668
rect 27692 24052 27748 24062
rect 27580 24050 27748 24052
rect 27580 23998 27694 24050
rect 27746 23998 27748 24050
rect 27580 23996 27748 23998
rect 27692 23986 27748 23996
rect 26908 23940 26964 23950
rect 26460 23938 26964 23940
rect 26460 23886 26910 23938
rect 26962 23886 26964 23938
rect 26460 23884 26964 23886
rect 26460 22372 26516 23884
rect 26908 23874 26964 23884
rect 26796 23714 26852 23726
rect 26796 23662 26798 23714
rect 26850 23662 26852 23714
rect 26796 23268 26852 23662
rect 26796 23202 26852 23212
rect 26908 23604 26964 23614
rect 26460 22370 26852 22372
rect 26460 22318 26462 22370
rect 26514 22318 26852 22370
rect 26460 22316 26852 22318
rect 26460 22306 26516 22316
rect 26348 21646 26350 21698
rect 26402 21646 26404 21698
rect 26348 21634 26404 21646
rect 26796 21586 26852 22316
rect 26796 21534 26798 21586
rect 26850 21534 26852 21586
rect 26796 21522 26852 21534
rect 26908 22370 26964 23548
rect 27580 23380 27636 23390
rect 27580 23286 27636 23324
rect 26908 22318 26910 22370
rect 26962 22318 26964 22370
rect 26908 21588 26964 22318
rect 27356 23268 27412 23278
rect 27244 21588 27300 21598
rect 26908 21586 27300 21588
rect 26908 21534 27246 21586
rect 27298 21534 27300 21586
rect 26908 21532 27300 21534
rect 27244 21522 27300 21532
rect 27356 20804 27412 23212
rect 27916 23042 27972 24780
rect 28028 23938 28084 25228
rect 28140 24946 28196 25452
rect 28924 25060 28980 26852
rect 29036 26516 29092 26526
rect 29036 26514 29316 26516
rect 29036 26462 29038 26514
rect 29090 26462 29316 26514
rect 29036 26460 29316 26462
rect 29036 26450 29092 26460
rect 29148 26292 29204 26302
rect 29148 26198 29204 26236
rect 29260 26068 29316 26460
rect 29372 26292 29428 27134
rect 30156 27748 30212 27758
rect 30156 26908 30212 27692
rect 30604 27076 30660 27086
rect 30940 27076 30996 28140
rect 30604 27074 30996 27076
rect 30604 27022 30606 27074
rect 30658 27022 30942 27074
rect 30994 27022 30996 27074
rect 30604 27020 30996 27022
rect 30604 27010 30660 27020
rect 30940 27010 30996 27020
rect 31052 27972 31108 27982
rect 31052 26908 31108 27916
rect 31276 27858 31332 28812
rect 31836 28756 31892 29260
rect 31948 29222 32004 29260
rect 31948 28756 32004 28766
rect 31836 28754 32004 28756
rect 31836 28702 31950 28754
rect 32002 28702 32004 28754
rect 31836 28700 32004 28702
rect 31948 28690 32004 28700
rect 32060 27972 32116 27982
rect 32060 27878 32116 27916
rect 31276 27806 31278 27858
rect 31330 27806 31332 27858
rect 31276 27794 31332 27806
rect 31500 27860 31556 27870
rect 31500 27766 31556 27804
rect 32508 27860 32564 27870
rect 32508 27766 32564 27804
rect 33404 27860 33460 27870
rect 31612 27748 31668 27758
rect 31612 27746 31780 27748
rect 31612 27694 31614 27746
rect 31666 27694 31780 27746
rect 31612 27692 31780 27694
rect 31612 27682 31668 27692
rect 31724 27186 31780 27692
rect 31724 27134 31726 27186
rect 31778 27134 31780 27186
rect 31724 27122 31780 27134
rect 29820 26852 30324 26908
rect 29820 26850 29876 26852
rect 29820 26798 29822 26850
rect 29874 26798 29876 26850
rect 29596 26516 29652 26526
rect 29820 26516 29876 26798
rect 29652 26460 29876 26516
rect 30268 26516 30324 26852
rect 30940 26852 31108 26908
rect 30828 26516 30884 26526
rect 30268 26514 30884 26516
rect 30268 26462 30270 26514
rect 30322 26462 30830 26514
rect 30882 26462 30884 26514
rect 30268 26460 30884 26462
rect 29596 26402 29652 26460
rect 30268 26450 30324 26460
rect 30828 26450 30884 26460
rect 29596 26350 29598 26402
rect 29650 26350 29652 26402
rect 29596 26338 29652 26350
rect 30156 26292 30212 26302
rect 29372 26226 29428 26236
rect 29708 26290 30212 26292
rect 29708 26238 30158 26290
rect 30210 26238 30212 26290
rect 29708 26236 30212 26238
rect 29484 26068 29540 26078
rect 29260 26066 29540 26068
rect 29260 26014 29486 26066
rect 29538 26014 29540 26066
rect 29260 26012 29540 26014
rect 29484 25394 29540 26012
rect 29484 25342 29486 25394
rect 29538 25342 29540 25394
rect 29484 25330 29540 25342
rect 29708 25506 29764 26236
rect 30156 26226 30212 26236
rect 30268 26068 30324 26078
rect 30268 25974 30324 26012
rect 29708 25454 29710 25506
rect 29762 25454 29764 25506
rect 29708 25284 29764 25454
rect 29708 25218 29764 25228
rect 29820 25394 29876 25406
rect 29820 25342 29822 25394
rect 29874 25342 29876 25394
rect 28140 24894 28142 24946
rect 28194 24894 28196 24946
rect 28140 24882 28196 24894
rect 28812 25004 28980 25060
rect 29484 25060 29540 25070
rect 28700 24724 28756 24734
rect 28028 23886 28030 23938
rect 28082 23886 28084 23938
rect 28028 23874 28084 23886
rect 28252 24722 28756 24724
rect 28252 24670 28702 24722
rect 28754 24670 28756 24722
rect 28252 24668 28756 24670
rect 28252 23940 28308 24668
rect 28700 24658 28756 24668
rect 28252 23826 28308 23884
rect 28252 23774 28254 23826
rect 28306 23774 28308 23826
rect 28252 23762 28308 23774
rect 28812 23268 28868 25004
rect 29036 24948 29092 24958
rect 28924 24892 29036 24948
rect 28924 24834 28980 24892
rect 29036 24882 29092 24892
rect 28924 24782 28926 24834
rect 28978 24782 28980 24834
rect 28924 24770 28980 24782
rect 29148 24836 29204 24846
rect 29148 24722 29204 24780
rect 29148 24670 29150 24722
rect 29202 24670 29204 24722
rect 29148 24658 29204 24670
rect 29484 24722 29540 25004
rect 29820 24836 29876 25342
rect 30940 25394 30996 26852
rect 33292 26180 33348 26190
rect 32396 25956 32452 25966
rect 32396 25506 32452 25900
rect 33180 25732 33236 25742
rect 33180 25638 33236 25676
rect 32396 25454 32398 25506
rect 32450 25454 32452 25506
rect 32396 25442 32452 25454
rect 32620 25508 32676 25518
rect 30940 25342 30942 25394
rect 30994 25342 30996 25394
rect 30940 25330 30996 25342
rect 32620 25394 32676 25452
rect 32732 25508 32788 25518
rect 33292 25508 33348 26124
rect 32732 25506 33348 25508
rect 32732 25454 32734 25506
rect 32786 25454 33294 25506
rect 33346 25454 33348 25506
rect 32732 25452 33348 25454
rect 32732 25442 32788 25452
rect 32620 25342 32622 25394
rect 32674 25342 32676 25394
rect 32620 25330 32676 25342
rect 31276 25282 31332 25294
rect 31276 25230 31278 25282
rect 31330 25230 31332 25282
rect 29932 25060 29988 25070
rect 29932 24946 29988 25004
rect 29932 24894 29934 24946
rect 29986 24894 29988 24946
rect 29932 24882 29988 24894
rect 31276 24948 31332 25230
rect 33180 25284 33236 25294
rect 33180 25190 33236 25228
rect 31388 24948 31444 24958
rect 31276 24946 31444 24948
rect 31276 24894 31390 24946
rect 31442 24894 31444 24946
rect 31276 24892 31444 24894
rect 29820 24770 29876 24780
rect 29484 24670 29486 24722
rect 29538 24670 29540 24722
rect 29484 24658 29540 24670
rect 29036 24610 29092 24622
rect 29036 24558 29038 24610
rect 29090 24558 29092 24610
rect 28812 23202 28868 23212
rect 28924 24388 28980 24398
rect 27916 22990 27918 23042
rect 27970 22990 27972 23042
rect 27916 22978 27972 22990
rect 27804 22260 27860 22270
rect 27916 22260 27972 22270
rect 27860 22258 27972 22260
rect 27860 22206 27918 22258
rect 27970 22206 27972 22258
rect 27860 22204 27972 22206
rect 27804 21698 27860 22204
rect 27916 22194 27972 22204
rect 28476 22146 28532 22158
rect 28476 22094 28478 22146
rect 28530 22094 28532 22146
rect 28476 21812 28532 22094
rect 28476 21746 28532 21756
rect 27804 21646 27806 21698
rect 27858 21646 27860 21698
rect 27804 21634 27860 21646
rect 27916 20804 27972 20814
rect 27356 20802 27972 20804
rect 27356 20750 27918 20802
rect 27970 20750 27972 20802
rect 27356 20748 27972 20750
rect 26796 20132 26852 20142
rect 26684 20076 26796 20132
rect 26572 20020 26628 20030
rect 26572 19926 26628 19964
rect 26236 19348 26292 19358
rect 26236 19254 26292 19292
rect 25004 19170 25060 19180
rect 26572 19236 26628 19246
rect 26684 19236 26740 20076
rect 26796 20038 26852 20076
rect 27132 20132 27188 20142
rect 27132 19908 27188 20076
rect 27244 20020 27300 20030
rect 27356 20020 27412 20748
rect 27916 20738 27972 20748
rect 27580 20580 27636 20590
rect 27468 20132 27524 20142
rect 27468 20038 27524 20076
rect 27244 20018 27356 20020
rect 27244 19966 27246 20018
rect 27298 19966 27356 20018
rect 27244 19964 27356 19966
rect 27244 19954 27300 19964
rect 27356 19954 27412 19964
rect 27580 19908 27636 20524
rect 28252 20578 28308 20590
rect 28252 20526 28254 20578
rect 28306 20526 28308 20578
rect 27916 20020 27972 20030
rect 28252 20020 28308 20526
rect 28924 20468 28980 24332
rect 29036 24052 29092 24558
rect 31276 24612 31332 24622
rect 29148 24052 29204 24062
rect 29036 24050 29204 24052
rect 29036 23998 29150 24050
rect 29202 23998 29204 24050
rect 29036 23996 29204 23998
rect 29148 23986 29204 23996
rect 29260 23716 29316 23726
rect 29260 23714 30100 23716
rect 29260 23662 29262 23714
rect 29314 23662 30100 23714
rect 29260 23660 30100 23662
rect 29260 23650 29316 23660
rect 30044 23266 30100 23660
rect 30044 23214 30046 23266
rect 30098 23214 30100 23266
rect 30044 23202 30100 23214
rect 30716 23380 30772 23390
rect 30716 23154 30772 23324
rect 30716 23102 30718 23154
rect 30770 23102 30772 23154
rect 30716 23090 30772 23102
rect 29260 20916 29316 20926
rect 28924 20402 28980 20412
rect 29036 20914 29316 20916
rect 29036 20862 29262 20914
rect 29314 20862 29316 20914
rect 29036 20860 29316 20862
rect 29036 20244 29092 20860
rect 29260 20850 29316 20860
rect 29372 20916 29428 20926
rect 29372 20802 29428 20860
rect 30156 20916 30212 20926
rect 30156 20822 30212 20860
rect 29372 20750 29374 20802
rect 29426 20750 29428 20802
rect 29372 20738 29428 20750
rect 30716 20804 30772 20814
rect 30772 20748 30996 20804
rect 30716 20710 30772 20748
rect 28588 20188 29092 20244
rect 29148 20690 29204 20702
rect 29148 20638 29150 20690
rect 29202 20638 29204 20690
rect 27916 20018 28084 20020
rect 27916 19966 27918 20018
rect 27970 19966 28084 20018
rect 27916 19964 28084 19966
rect 27916 19954 27972 19964
rect 27132 19842 27188 19852
rect 27468 19852 27636 19908
rect 27692 19908 27748 19918
rect 26572 19234 26740 19236
rect 26572 19182 26574 19234
rect 26626 19182 26740 19234
rect 26572 19180 26740 19182
rect 26796 19348 26852 19358
rect 26796 19234 26852 19292
rect 26796 19182 26798 19234
rect 26850 19182 26852 19234
rect 26572 19170 26628 19180
rect 26796 19170 26852 19182
rect 27132 19122 27188 19134
rect 27132 19070 27134 19122
rect 27186 19070 27188 19122
rect 23996 19010 24052 19022
rect 23996 18958 23998 19010
rect 24050 18958 24052 19010
rect 23996 18564 24052 18958
rect 26684 19010 26740 19022
rect 26684 18958 26686 19010
rect 26738 18958 26740 19010
rect 26684 18676 26740 18958
rect 26012 18620 26740 18676
rect 24220 18564 24276 18574
rect 23996 18508 24220 18564
rect 24220 18450 24276 18508
rect 24220 18398 24222 18450
rect 24274 18398 24276 18450
rect 24220 18386 24276 18398
rect 24444 18562 24500 18574
rect 24444 18510 24446 18562
rect 24498 18510 24500 18562
rect 23772 18340 23828 18350
rect 23772 18246 23828 18284
rect 24444 18340 24500 18510
rect 26012 18562 26068 18620
rect 26012 18510 26014 18562
rect 26066 18510 26068 18562
rect 26012 18498 26068 18510
rect 24444 18116 24500 18284
rect 25340 18450 25396 18462
rect 25340 18398 25342 18450
rect 25394 18398 25396 18450
rect 24444 18050 24500 18060
rect 25004 18228 25060 18238
rect 23100 17388 23380 17444
rect 22988 16100 23044 16110
rect 22876 16098 23044 16100
rect 22876 16046 22990 16098
rect 23042 16046 23044 16098
rect 22876 16044 23044 16046
rect 22988 16034 23044 16044
rect 22988 15876 23044 15886
rect 22988 15782 23044 15820
rect 23100 15148 23156 17388
rect 24668 16212 24724 16222
rect 23324 15988 23380 15998
rect 24444 15988 24500 15998
rect 18732 14084 18788 15092
rect 22204 15090 22260 15102
rect 22428 15092 22596 15148
rect 22652 15092 22820 15148
rect 22204 15038 22206 15090
rect 22258 15038 22260 15090
rect 22204 14532 22260 15038
rect 22260 14476 22484 14532
rect 22204 14466 22260 14476
rect 18844 14308 18900 14318
rect 18844 14306 19012 14308
rect 18844 14254 18846 14306
rect 18898 14254 19012 14306
rect 18844 14252 19012 14254
rect 18844 14242 18900 14252
rect 18732 14018 18788 14028
rect 18732 13746 18788 13758
rect 18732 13694 18734 13746
rect 18786 13694 18788 13746
rect 18732 13636 18788 13694
rect 18844 13748 18900 13758
rect 18844 13654 18900 13692
rect 18956 13748 19012 14252
rect 22092 14306 22148 14318
rect 22092 14254 22094 14306
rect 22146 14254 22148 14306
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20748 13972 20804 13982
rect 20748 13878 20804 13916
rect 21308 13972 21364 13982
rect 21084 13860 21140 13870
rect 19404 13748 19460 13758
rect 18956 13746 19460 13748
rect 18956 13694 18958 13746
rect 19010 13694 19406 13746
rect 19458 13694 19460 13746
rect 18956 13692 19460 13694
rect 18956 13682 19012 13692
rect 19404 13682 19460 13692
rect 19628 13746 19684 13758
rect 19628 13694 19630 13746
rect 19682 13694 19684 13746
rect 18732 13570 18788 13580
rect 19516 13524 19572 13534
rect 18620 12910 18622 12962
rect 18674 12910 18676 12962
rect 18620 12898 18676 12910
rect 18732 13076 18788 13086
rect 19180 13076 19236 13086
rect 18732 13074 19236 13076
rect 18732 13022 18734 13074
rect 18786 13022 19182 13074
rect 19234 13022 19236 13074
rect 18732 13020 19236 13022
rect 18732 12964 18788 13020
rect 19180 13010 19236 13020
rect 18732 12898 18788 12908
rect 18844 12852 18900 12862
rect 18844 12850 19236 12852
rect 18844 12798 18846 12850
rect 18898 12798 19236 12850
rect 18844 12796 19236 12798
rect 18844 12740 18900 12796
rect 18508 12684 18900 12740
rect 18340 11452 18452 11508
rect 18508 12516 18564 12526
rect 18284 11442 18340 11452
rect 18060 10670 18062 10722
rect 18114 10670 18116 10722
rect 18060 10658 18116 10670
rect 18172 10834 18228 10846
rect 18172 10782 18174 10834
rect 18226 10782 18228 10834
rect 17724 10050 17836 10052
rect 17724 9998 17726 10050
rect 17778 9998 17836 10050
rect 17724 9996 17836 9998
rect 17724 9986 17780 9996
rect 17836 9958 17892 9996
rect 17948 10610 18004 10622
rect 17948 10558 17950 10610
rect 18002 10558 18004 10610
rect 17948 9828 18004 10558
rect 18060 10052 18116 10062
rect 18172 10052 18228 10782
rect 18396 10724 18452 10734
rect 18396 10630 18452 10668
rect 18060 10050 18228 10052
rect 18060 9998 18062 10050
rect 18114 9998 18228 10050
rect 18060 9996 18228 9998
rect 18060 9986 18116 9996
rect 17948 9762 18004 9772
rect 17500 9214 17502 9266
rect 17554 9214 17556 9266
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 15484 6692 15540 6702
rect 15484 6598 15540 6636
rect 17500 6692 17556 9214
rect 18172 9268 18228 9996
rect 18172 9202 18228 9212
rect 18284 9826 18340 9838
rect 18284 9774 18286 9826
rect 18338 9774 18340 9826
rect 18284 9044 18340 9774
rect 18284 8978 18340 8988
rect 18508 8428 18564 12460
rect 18732 11844 18788 11854
rect 18620 11788 18732 11844
rect 18620 10724 18676 11788
rect 18732 11778 18788 11788
rect 18732 11508 18788 11518
rect 19180 11508 19236 12796
rect 18788 11452 19124 11508
rect 18732 11394 18788 11452
rect 18732 11342 18734 11394
rect 18786 11342 18788 11394
rect 18732 11330 18788 11342
rect 18956 11282 19012 11294
rect 18956 11230 18958 11282
rect 19010 11230 19012 11282
rect 18844 11172 18900 11182
rect 18844 11078 18900 11116
rect 18732 10724 18788 10734
rect 18620 10722 18788 10724
rect 18620 10670 18734 10722
rect 18786 10670 18788 10722
rect 18620 10668 18788 10670
rect 18732 10658 18788 10668
rect 18956 10612 19012 11230
rect 18844 10556 19012 10612
rect 18844 10388 18900 10556
rect 19068 10500 19124 11452
rect 19292 12738 19348 12750
rect 19292 12686 19294 12738
rect 19346 12686 19348 12738
rect 19292 11508 19348 12686
rect 19404 12740 19460 12750
rect 19404 12646 19460 12684
rect 19516 12290 19572 13468
rect 19628 13412 19684 13694
rect 19852 13746 19908 13758
rect 20860 13748 20916 13758
rect 19852 13694 19854 13746
rect 19906 13694 19908 13746
rect 19852 13636 19908 13694
rect 20524 13746 20916 13748
rect 20524 13694 20862 13746
rect 20914 13694 20916 13746
rect 20524 13692 20916 13694
rect 20412 13636 20468 13646
rect 19908 13580 20132 13636
rect 19852 13570 19908 13580
rect 19628 13346 19684 13356
rect 19964 13188 20020 13198
rect 19516 12238 19518 12290
rect 19570 12238 19572 12290
rect 19516 11732 19572 12238
rect 19516 11666 19572 11676
rect 19628 13186 20020 13188
rect 19628 13134 19966 13186
rect 20018 13134 20020 13186
rect 19628 13132 20020 13134
rect 20076 13188 20132 13580
rect 20412 13522 20468 13580
rect 20412 13470 20414 13522
rect 20466 13470 20468 13522
rect 20412 13458 20468 13470
rect 20076 13132 20356 13188
rect 19628 11618 19684 13132
rect 19964 13122 20020 13132
rect 19852 12964 19908 12974
rect 19852 12870 19908 12908
rect 20300 12852 20356 13132
rect 20524 13186 20580 13692
rect 20860 13682 20916 13692
rect 21084 13746 21140 13804
rect 21084 13694 21086 13746
rect 21138 13694 21140 13746
rect 21084 13682 21140 13694
rect 21308 13746 21364 13916
rect 22092 13860 22148 14254
rect 22092 13794 22148 13804
rect 22204 13972 22260 13982
rect 21308 13694 21310 13746
rect 21362 13694 21364 13746
rect 21308 13682 21364 13694
rect 21420 13746 21476 13758
rect 21420 13694 21422 13746
rect 21474 13694 21476 13746
rect 20524 13134 20526 13186
rect 20578 13134 20580 13186
rect 20524 13122 20580 13134
rect 21196 13636 21252 13646
rect 21196 13188 21252 13580
rect 21308 13188 21364 13198
rect 21196 13186 21364 13188
rect 21196 13134 21310 13186
rect 21362 13134 21364 13186
rect 21196 13132 21364 13134
rect 21308 13122 21364 13132
rect 21420 13074 21476 13694
rect 21756 13748 21812 13758
rect 21756 13654 21812 13692
rect 22204 13634 22260 13916
rect 22428 13746 22484 14476
rect 22540 14420 22596 15092
rect 22652 14420 22708 14430
rect 22540 14364 22652 14420
rect 22652 14326 22708 14364
rect 22428 13694 22430 13746
rect 22482 13694 22484 13746
rect 22428 13682 22484 13694
rect 22652 13748 22708 13758
rect 22652 13654 22708 13692
rect 22764 13746 22820 15092
rect 22876 15092 23156 15148
rect 23212 15986 23380 15988
rect 23212 15934 23326 15986
rect 23378 15934 23380 15986
rect 23212 15932 23380 15934
rect 23212 15148 23268 15932
rect 23324 15922 23380 15932
rect 24220 15986 24500 15988
rect 24220 15934 24446 15986
rect 24498 15934 24500 15986
rect 24220 15932 24500 15934
rect 23660 15876 23716 15886
rect 23660 15202 23716 15820
rect 24220 15426 24276 15932
rect 24444 15922 24500 15932
rect 24668 15986 24724 16156
rect 24668 15934 24670 15986
rect 24722 15934 24724 15986
rect 24668 15922 24724 15934
rect 24220 15374 24222 15426
rect 24274 15374 24276 15426
rect 24220 15362 24276 15374
rect 24556 15874 24612 15886
rect 24556 15822 24558 15874
rect 24610 15822 24612 15874
rect 23660 15150 23662 15202
rect 23714 15150 23716 15202
rect 23212 15092 23380 15148
rect 23660 15138 23716 15150
rect 23772 15314 23828 15326
rect 23772 15262 23774 15314
rect 23826 15262 23828 15314
rect 22876 13972 22932 15092
rect 23324 14644 23380 15092
rect 23324 14578 23380 14588
rect 23548 14530 23604 14542
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 22876 13906 22932 13916
rect 23212 14308 23268 14318
rect 23548 14308 23604 14478
rect 23212 14306 23604 14308
rect 23212 14254 23214 14306
rect 23266 14254 23604 14306
rect 23212 14252 23604 14254
rect 22988 13748 23044 13758
rect 22764 13694 22766 13746
rect 22818 13694 22820 13746
rect 22764 13682 22820 13694
rect 22876 13746 23044 13748
rect 22876 13694 22990 13746
rect 23042 13694 23044 13746
rect 22876 13692 23044 13694
rect 22204 13582 22206 13634
rect 22258 13582 22260 13634
rect 22204 13524 22260 13582
rect 22204 13468 22708 13524
rect 21420 13022 21422 13074
rect 21474 13022 21476 13074
rect 21420 13010 21476 13022
rect 21644 12962 21700 12974
rect 21644 12910 21646 12962
rect 21698 12910 21700 12962
rect 20412 12852 20468 12862
rect 20300 12850 20468 12852
rect 20300 12798 20414 12850
rect 20466 12798 20468 12850
rect 20300 12796 20468 12798
rect 21644 12852 21700 12910
rect 22092 12852 22148 12862
rect 22428 12852 22484 12862
rect 21644 12850 22484 12852
rect 21644 12798 22094 12850
rect 22146 12798 22430 12850
rect 22482 12798 22484 12850
rect 21644 12796 22484 12798
rect 19964 12740 20020 12750
rect 19964 12738 20244 12740
rect 19964 12686 19966 12738
rect 20018 12686 20244 12738
rect 19964 12684 20244 12686
rect 19964 12674 20020 12684
rect 20188 12628 20244 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20188 12562 20244 12572
rect 19836 12506 20100 12516
rect 20188 11844 20244 11854
rect 20300 11844 20356 12796
rect 20412 12786 20468 12796
rect 22092 12786 22148 12796
rect 20860 12628 20916 12638
rect 20860 12402 20916 12572
rect 20860 12350 20862 12402
rect 20914 12350 20916 12402
rect 20860 12338 20916 12350
rect 22428 12404 22484 12796
rect 22540 12852 22596 12862
rect 22540 12758 22596 12796
rect 22428 12338 22484 12348
rect 21196 12068 21252 12078
rect 21196 11974 21252 12012
rect 20244 11788 20356 11844
rect 20188 11778 20244 11788
rect 19628 11566 19630 11618
rect 19682 11566 19684 11618
rect 19628 11554 19684 11566
rect 22652 11620 22708 13468
rect 22652 11554 22708 11564
rect 22764 12852 22820 12862
rect 22876 12852 22932 13692
rect 22988 13682 23044 13692
rect 23212 13524 23268 14252
rect 23212 13458 23268 13468
rect 23324 13748 23380 13758
rect 23660 13748 23716 13758
rect 23324 12962 23380 13692
rect 23548 13746 23716 13748
rect 23548 13694 23662 13746
rect 23714 13694 23716 13746
rect 23548 13692 23716 13694
rect 23548 13636 23604 13692
rect 23660 13682 23716 13692
rect 23548 13186 23604 13580
rect 23772 13636 23828 15262
rect 24332 14644 24388 14654
rect 24556 14644 24612 15822
rect 24332 14642 24612 14644
rect 24332 14590 24334 14642
rect 24386 14590 24612 14642
rect 24332 14588 24612 14590
rect 24332 14578 24388 14588
rect 24332 14308 24388 14318
rect 23884 13972 23940 13982
rect 24332 13972 24388 14252
rect 23884 13970 24388 13972
rect 23884 13918 23886 13970
rect 23938 13918 24334 13970
rect 24386 13918 24388 13970
rect 23884 13916 24388 13918
rect 23884 13906 23940 13916
rect 24332 13906 24388 13916
rect 23772 13634 24276 13636
rect 23772 13582 23774 13634
rect 23826 13582 24276 13634
rect 23772 13580 24276 13582
rect 23772 13570 23828 13580
rect 23548 13134 23550 13186
rect 23602 13134 23604 13186
rect 23548 13122 23604 13134
rect 23324 12910 23326 12962
rect 23378 12910 23380 12962
rect 23324 12898 23380 12910
rect 23772 12964 23828 12974
rect 23828 12908 24052 12964
rect 23772 12870 23828 12908
rect 22764 12850 22932 12852
rect 22764 12798 22766 12850
rect 22818 12798 22932 12850
rect 22764 12796 22932 12798
rect 22988 12850 23044 12862
rect 22988 12798 22990 12850
rect 23042 12798 23044 12850
rect 19516 11508 19572 11518
rect 19292 11506 19572 11508
rect 19292 11454 19518 11506
rect 19570 11454 19572 11506
rect 19292 11452 19572 11454
rect 19180 11442 19236 11452
rect 19516 11442 19572 11452
rect 21308 11508 21364 11518
rect 18732 9828 18788 9838
rect 18844 9828 18900 10332
rect 18956 10444 19124 10500
rect 19292 11282 19348 11294
rect 19292 11230 19294 11282
rect 19346 11230 19348 11282
rect 18956 10386 19012 10444
rect 18956 10334 18958 10386
rect 19010 10334 19012 10386
rect 18956 10322 19012 10334
rect 19180 10386 19236 10398
rect 19180 10334 19182 10386
rect 19234 10334 19236 10386
rect 18956 9828 19012 9838
rect 18844 9826 19012 9828
rect 18844 9774 18958 9826
rect 19010 9774 19012 9826
rect 18844 9772 19012 9774
rect 18732 9734 18788 9772
rect 18956 9762 19012 9772
rect 19180 9828 19236 10334
rect 19180 9762 19236 9772
rect 19292 9716 19348 11230
rect 21308 11282 21364 11452
rect 21308 11230 21310 11282
rect 21362 11230 21364 11282
rect 21308 11218 21364 11230
rect 21532 11394 21588 11406
rect 21532 11342 21534 11394
rect 21586 11342 21588 11394
rect 20188 11170 20244 11182
rect 20188 11118 20190 11170
rect 20242 11118 20244 11170
rect 20188 11060 20244 11118
rect 20300 11060 20356 11070
rect 19836 11004 20100 11014
rect 20188 11004 20300 11060
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20300 10612 20356 11004
rect 20076 10556 20356 10612
rect 21532 10724 21588 11342
rect 19292 9622 19348 9660
rect 19404 10386 19460 10398
rect 19404 10334 19406 10386
rect 19458 10334 19460 10386
rect 18844 9604 18900 9614
rect 18844 9510 18900 9548
rect 18732 9268 18788 9278
rect 18956 9268 19012 9278
rect 18732 9174 18788 9212
rect 18844 9212 18956 9268
rect 18844 9154 18900 9212
rect 18956 9202 19012 9212
rect 18844 9102 18846 9154
rect 18898 9102 18900 9154
rect 18844 9090 18900 9102
rect 18956 9044 19012 9054
rect 18956 8950 19012 8988
rect 19292 9042 19348 9054
rect 19292 8990 19294 9042
rect 19346 8990 19348 9042
rect 18508 8372 19012 8428
rect 18844 7924 18900 7934
rect 18844 7474 18900 7868
rect 18956 7586 19012 8372
rect 19292 8036 19348 8990
rect 19292 7970 19348 7980
rect 19404 7924 19460 10334
rect 19852 10386 19908 10398
rect 19852 10334 19854 10386
rect 19906 10334 19908 10386
rect 19516 10052 19572 10062
rect 19516 9958 19572 9996
rect 19628 9826 19684 9838
rect 19628 9774 19630 9826
rect 19682 9774 19684 9826
rect 19628 9268 19684 9774
rect 19852 9716 19908 10334
rect 20076 10388 20132 10556
rect 20076 9938 20132 10332
rect 20076 9886 20078 9938
rect 20130 9886 20132 9938
rect 20076 9874 20132 9886
rect 19852 9650 19908 9660
rect 20412 9604 20468 9614
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 9202 19684 9212
rect 19404 7858 19460 7868
rect 19516 9044 19572 9054
rect 18956 7534 18958 7586
rect 19010 7534 19012 7586
rect 18956 7522 19012 7534
rect 19068 7698 19124 7710
rect 19068 7646 19070 7698
rect 19122 7646 19124 7698
rect 19068 7588 19124 7646
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 17724 6804 17780 6814
rect 16156 6580 16212 6590
rect 16156 6486 16212 6524
rect 17388 6580 17444 6590
rect 17388 6130 17444 6524
rect 17388 6078 17390 6130
rect 17442 6078 17444 6130
rect 17388 6066 17444 6078
rect 17500 6132 17556 6636
rect 17500 6066 17556 6076
rect 17612 6748 17724 6804
rect 17500 5908 17556 5918
rect 17612 5908 17668 6748
rect 17724 6738 17780 6748
rect 18284 6804 18340 6814
rect 18620 6804 18676 6814
rect 18284 6802 18564 6804
rect 18284 6750 18286 6802
rect 18338 6750 18564 6802
rect 18284 6748 18564 6750
rect 18284 6738 18340 6748
rect 18508 6580 18564 6748
rect 18620 6710 18676 6748
rect 18732 6692 18788 6702
rect 18844 6692 18900 7422
rect 18732 6690 18900 6692
rect 18732 6638 18734 6690
rect 18786 6638 18900 6690
rect 18732 6636 18900 6638
rect 18732 6580 18788 6636
rect 18508 6524 18788 6580
rect 18956 6580 19012 6590
rect 18956 6486 19012 6524
rect 17500 5906 17668 5908
rect 17500 5854 17502 5906
rect 17554 5854 17668 5906
rect 17500 5852 17668 5854
rect 18396 6132 18452 6142
rect 17500 5842 17556 5852
rect 18396 5794 18452 6076
rect 19068 5906 19124 7532
rect 19404 7476 19460 7486
rect 19404 7382 19460 7420
rect 19292 7252 19348 7262
rect 19180 6468 19236 6478
rect 19180 6374 19236 6412
rect 19068 5854 19070 5906
rect 19122 5854 19124 5906
rect 19068 5842 19124 5854
rect 19292 5906 19348 7196
rect 19292 5854 19294 5906
rect 19346 5854 19348 5906
rect 19292 5842 19348 5854
rect 19516 6914 19572 8988
rect 20300 8036 20356 8046
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19628 7588 19684 7598
rect 19628 7494 19684 7532
rect 19852 7474 19908 7486
rect 19852 7422 19854 7474
rect 19906 7422 19908 7474
rect 19740 7362 19796 7374
rect 19740 7310 19742 7362
rect 19794 7310 19796 7362
rect 19516 6862 19518 6914
rect 19570 6862 19572 6914
rect 18396 5742 18398 5794
rect 18450 5742 18452 5794
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 18396 5236 18452 5742
rect 18732 5684 18788 5694
rect 19516 5684 19572 6862
rect 19628 6916 19684 6926
rect 19740 6916 19796 7310
rect 19852 7252 19908 7422
rect 19852 7186 19908 7196
rect 20300 7474 20356 7980
rect 20300 7422 20302 7474
rect 20354 7422 20356 7474
rect 19628 6914 19796 6916
rect 19628 6862 19630 6914
rect 19682 6862 19796 6914
rect 19628 6860 19796 6862
rect 19628 6850 19684 6860
rect 20188 6804 20244 6814
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 18732 5682 19572 5684
rect 18732 5630 18734 5682
rect 18786 5630 19572 5682
rect 18732 5628 19572 5630
rect 18732 5618 18788 5628
rect 18396 4338 18452 5180
rect 20188 5234 20244 6748
rect 20300 6466 20356 7422
rect 20300 6414 20302 6466
rect 20354 6414 20356 6466
rect 20300 6356 20356 6414
rect 20412 6468 20468 9548
rect 21420 9604 21476 9614
rect 21420 9510 21476 9548
rect 21532 9268 21588 10668
rect 21644 10498 21700 10510
rect 21644 10446 21646 10498
rect 21698 10446 21700 10498
rect 21644 10388 21700 10446
rect 21644 10322 21700 10332
rect 22764 10388 22820 12796
rect 22988 12740 23044 12798
rect 23436 12740 23492 12750
rect 22988 12738 23492 12740
rect 22988 12686 23438 12738
rect 23490 12686 23492 12738
rect 22988 12684 23492 12686
rect 23436 12674 23492 12684
rect 23996 12628 24052 12908
rect 24108 12962 24164 12974
rect 24108 12910 24110 12962
rect 24162 12910 24164 12962
rect 24108 12852 24164 12910
rect 24220 12964 24276 13580
rect 24556 13524 24612 13534
rect 24444 12964 24500 12974
rect 24220 12962 24500 12964
rect 24220 12910 24446 12962
rect 24498 12910 24500 12962
rect 24220 12908 24500 12910
rect 24444 12898 24500 12908
rect 24108 12786 24164 12796
rect 24332 12738 24388 12750
rect 24332 12686 24334 12738
rect 24386 12686 24388 12738
rect 23996 12572 24276 12628
rect 23324 12404 23380 12414
rect 23324 12310 23380 12348
rect 24220 12402 24276 12572
rect 24220 12350 24222 12402
rect 24274 12350 24276 12402
rect 24220 12338 24276 12350
rect 24332 11620 24388 12686
rect 24556 12404 24612 13468
rect 24780 12850 24836 12862
rect 24780 12798 24782 12850
rect 24834 12798 24836 12850
rect 24780 12740 24836 12798
rect 24780 12674 24836 12684
rect 23772 11564 24388 11620
rect 24444 12402 24612 12404
rect 24444 12350 24558 12402
rect 24610 12350 24612 12402
rect 24444 12348 24612 12350
rect 23772 10722 23828 11564
rect 24332 11396 24388 11406
rect 24444 11396 24500 12348
rect 24556 12338 24612 12348
rect 24332 11394 24500 11396
rect 24332 11342 24334 11394
rect 24386 11342 24500 11394
rect 24332 11340 24500 11342
rect 24668 11506 24724 11518
rect 24668 11454 24670 11506
rect 24722 11454 24724 11506
rect 24332 11330 24388 11340
rect 23772 10670 23774 10722
rect 23826 10670 23828 10722
rect 23772 10658 23828 10670
rect 23996 11170 24052 11182
rect 23996 11118 23998 11170
rect 24050 11118 24052 11170
rect 22764 10322 22820 10332
rect 21756 9940 21812 9950
rect 21756 9826 21812 9884
rect 22204 9940 22260 9950
rect 22204 9846 22260 9884
rect 21756 9774 21758 9826
rect 21810 9774 21812 9826
rect 21756 9762 21812 9774
rect 23436 9716 23492 9726
rect 23436 9622 23492 9660
rect 22092 9268 22148 9278
rect 21532 9266 22148 9268
rect 21532 9214 22094 9266
rect 22146 9214 22148 9266
rect 21532 9212 22148 9214
rect 21532 7476 21588 9212
rect 22092 9202 22148 9212
rect 22428 9042 22484 9054
rect 22428 8990 22430 9042
rect 22482 8990 22484 9042
rect 22428 8484 22484 8990
rect 22428 8418 22484 8428
rect 23996 8428 24052 11118
rect 24556 10612 24612 10622
rect 24556 10518 24612 10556
rect 24668 10164 24724 11454
rect 24668 8428 24724 10108
rect 25004 9940 25060 18172
rect 25340 17444 25396 18398
rect 27132 18452 27188 19070
rect 27132 18386 27188 18396
rect 25340 17378 25396 17388
rect 25228 16212 25284 16222
rect 25228 16118 25284 16156
rect 27468 15988 27524 19852
rect 27580 16996 27636 17006
rect 27580 16902 27636 16940
rect 27692 16882 27748 19852
rect 27916 18340 27972 18350
rect 27916 18116 27972 18284
rect 27916 18050 27972 18060
rect 28028 17444 28084 19964
rect 28252 19954 28308 19964
rect 28476 20132 28532 20142
rect 28476 19012 28532 20076
rect 28588 20130 28644 20188
rect 28588 20078 28590 20130
rect 28642 20078 28644 20130
rect 28588 20066 28644 20078
rect 29148 19908 29204 20638
rect 29708 20692 29764 20702
rect 29708 20690 30100 20692
rect 29708 20638 29710 20690
rect 29762 20638 30100 20690
rect 29708 20636 30100 20638
rect 29708 20626 29764 20636
rect 29148 19842 29204 19852
rect 30044 19346 30100 20636
rect 30044 19294 30046 19346
rect 30098 19294 30100 19346
rect 30044 19282 30100 19294
rect 30492 20020 30548 20030
rect 28476 18674 28532 18956
rect 29932 19012 29988 19022
rect 29932 18918 29988 18956
rect 30156 19012 30212 19022
rect 30156 18918 30212 18956
rect 28476 18622 28478 18674
rect 28530 18622 28532 18674
rect 28476 18610 28532 18622
rect 29372 18676 29428 18686
rect 28700 18562 28756 18574
rect 28700 18510 28702 18562
rect 28754 18510 28756 18562
rect 28588 18452 28644 18462
rect 28588 18358 28644 18396
rect 28140 18340 28196 18350
rect 28140 18246 28196 18284
rect 28700 18340 28756 18510
rect 28364 17444 28420 17454
rect 28084 17442 28420 17444
rect 28084 17390 28366 17442
rect 28418 17390 28420 17442
rect 28084 17388 28420 17390
rect 28028 17350 28084 17388
rect 28364 17108 28420 17388
rect 28700 17220 28756 18284
rect 29148 18450 29204 18462
rect 29148 18398 29150 18450
rect 29202 18398 29204 18450
rect 29148 18340 29204 18398
rect 29148 18116 29204 18284
rect 29148 18050 29204 18060
rect 28924 17668 28980 17678
rect 28700 17154 28756 17164
rect 28812 17612 28924 17668
rect 28364 17042 28420 17052
rect 28812 17108 28868 17612
rect 28924 17602 28980 17612
rect 28812 17052 29204 17108
rect 28140 16996 28196 17006
rect 28140 16902 28196 16940
rect 28700 16996 28756 17006
rect 28812 16996 28868 17052
rect 28700 16994 28868 16996
rect 28700 16942 28702 16994
rect 28754 16942 28868 16994
rect 28700 16940 28868 16942
rect 28700 16930 28756 16940
rect 27692 16830 27694 16882
rect 27746 16830 27748 16882
rect 27692 16098 27748 16830
rect 28252 16882 28308 16894
rect 28252 16830 28254 16882
rect 28306 16830 28308 16882
rect 27916 16772 27972 16782
rect 28252 16772 28308 16830
rect 28924 16882 28980 16894
rect 28924 16830 28926 16882
rect 28978 16830 28980 16882
rect 27916 16770 28084 16772
rect 27916 16718 27918 16770
rect 27970 16718 28084 16770
rect 27916 16716 28084 16718
rect 27916 16706 27972 16716
rect 27692 16046 27694 16098
rect 27746 16046 27748 16098
rect 27692 16034 27748 16046
rect 27468 15894 27524 15932
rect 27916 15874 27972 15886
rect 27916 15822 27918 15874
rect 27970 15822 27972 15874
rect 27916 15540 27972 15822
rect 27356 15484 27972 15540
rect 27356 15426 27412 15484
rect 27356 15374 27358 15426
rect 27410 15374 27412 15426
rect 27356 15362 27412 15374
rect 26684 15314 26740 15326
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 15204 26740 15262
rect 26684 15148 26964 15204
rect 26908 15092 27076 15148
rect 25788 14644 25844 14654
rect 25228 12740 25284 12750
rect 25228 12646 25284 12684
rect 25340 10612 25396 10650
rect 25340 10546 25396 10556
rect 25004 9874 25060 9884
rect 25340 10388 25396 10398
rect 24892 9826 24948 9838
rect 24892 9774 24894 9826
rect 24946 9774 24948 9826
rect 24892 8428 24948 9774
rect 25340 9826 25396 10332
rect 25340 9774 25342 9826
rect 25394 9774 25396 9826
rect 25340 9762 25396 9774
rect 25788 9716 25844 14588
rect 26460 14644 26516 14654
rect 26460 14550 26516 14588
rect 26796 14420 26852 14430
rect 26796 14326 26852 14364
rect 27020 13748 27076 15092
rect 27580 14644 27636 14654
rect 27580 14550 27636 14588
rect 27132 14308 27188 14318
rect 27188 14252 27300 14308
rect 27132 14214 27188 14252
rect 27132 13748 27188 13758
rect 27020 13746 27188 13748
rect 27020 13694 27134 13746
rect 27186 13694 27188 13746
rect 27020 13692 27188 13694
rect 27020 12740 27076 12750
rect 26908 12684 27020 12740
rect 26796 11282 26852 11294
rect 26796 11230 26798 11282
rect 26850 11230 26852 11282
rect 25900 10836 25956 10846
rect 26236 10836 26292 10846
rect 25900 10834 26236 10836
rect 25900 10782 25902 10834
rect 25954 10782 26236 10834
rect 25900 10780 26236 10782
rect 25900 10770 25956 10780
rect 26236 10742 26292 10780
rect 26348 10780 26740 10836
rect 26348 10722 26404 10780
rect 26348 10670 26350 10722
rect 26402 10670 26404 10722
rect 26348 10658 26404 10670
rect 26572 10610 26628 10622
rect 26572 10558 26574 10610
rect 26626 10558 26628 10610
rect 26236 10388 26292 10398
rect 26572 10388 26628 10558
rect 26236 10386 26628 10388
rect 26236 10334 26238 10386
rect 26290 10334 26628 10386
rect 26236 10332 26628 10334
rect 26236 10322 26292 10332
rect 26572 9828 26628 9838
rect 25900 9716 25956 9726
rect 25788 9714 25956 9716
rect 25788 9662 25902 9714
rect 25954 9662 25956 9714
rect 25788 9660 25956 9662
rect 25900 9650 25956 9660
rect 23996 8372 24276 8428
rect 23548 7532 23828 7588
rect 21308 7362 21364 7374
rect 21308 7310 21310 7362
rect 21362 7310 21364 7362
rect 20748 7252 20804 7262
rect 20748 7158 20804 7196
rect 21084 7252 21140 7262
rect 21084 7250 21252 7252
rect 21084 7198 21086 7250
rect 21138 7198 21252 7250
rect 21084 7196 21252 7198
rect 21084 7186 21140 7196
rect 20524 7028 20580 7038
rect 20524 6690 20580 6972
rect 20524 6638 20526 6690
rect 20578 6638 20580 6690
rect 20524 6626 20580 6638
rect 20636 6802 20692 6814
rect 20636 6750 20638 6802
rect 20690 6750 20692 6802
rect 20636 6692 20692 6750
rect 20636 6626 20692 6636
rect 20412 6402 20468 6412
rect 20748 6466 20804 6478
rect 20748 6414 20750 6466
rect 20802 6414 20804 6466
rect 20748 6356 20804 6414
rect 21196 6356 21252 7196
rect 21308 7028 21364 7310
rect 21308 6962 21364 6972
rect 21420 7252 21476 7262
rect 21420 6914 21476 7196
rect 21420 6862 21422 6914
rect 21474 6862 21476 6914
rect 21420 6850 21476 6862
rect 21308 6802 21364 6814
rect 21308 6750 21310 6802
rect 21362 6750 21364 6802
rect 21308 6692 21364 6750
rect 21308 6626 21364 6636
rect 20748 6300 21364 6356
rect 20300 6290 20356 6300
rect 20188 5182 20190 5234
rect 20242 5182 20244 5234
rect 20188 5170 20244 5182
rect 21196 5908 21252 5918
rect 20076 4900 20132 4910
rect 19068 4898 20132 4900
rect 19068 4846 20078 4898
rect 20130 4846 20132 4898
rect 19068 4844 20132 4846
rect 19068 4450 19124 4844
rect 20076 4834 20132 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4398 19070 4450
rect 19122 4398 19124 4450
rect 19068 4386 19124 4398
rect 18396 4286 18398 4338
rect 18450 4286 18452 4338
rect 18396 4274 18452 4286
rect 21196 4226 21252 5852
rect 21308 5796 21364 6300
rect 21532 6018 21588 7420
rect 23324 7476 23380 7486
rect 23548 7476 23604 7532
rect 23324 7474 23604 7476
rect 23324 7422 23326 7474
rect 23378 7422 23604 7474
rect 23324 7420 23604 7422
rect 23324 7410 23380 7420
rect 23660 7362 23716 7374
rect 23660 7310 23662 7362
rect 23714 7310 23716 7362
rect 22764 7250 22820 7262
rect 22764 7198 22766 7250
rect 22818 7198 22820 7250
rect 22764 7028 22820 7198
rect 23100 7252 23156 7262
rect 23100 7250 23268 7252
rect 23100 7198 23102 7250
rect 23154 7198 23268 7250
rect 23100 7196 23268 7198
rect 23100 7186 23156 7196
rect 23212 7028 23268 7196
rect 23548 7028 23604 7038
rect 23212 6972 23380 7028
rect 22764 6962 22820 6972
rect 22204 6804 22260 6842
rect 22204 6738 22260 6748
rect 23212 6804 23268 6814
rect 21980 6580 22036 6590
rect 21980 6486 22036 6524
rect 22204 6578 22260 6590
rect 22204 6526 22206 6578
rect 22258 6526 22260 6578
rect 21756 6468 21812 6478
rect 21756 6374 21812 6412
rect 22204 6468 22260 6526
rect 21532 5966 21534 6018
rect 21586 5966 21588 6018
rect 21532 5954 21588 5966
rect 21756 5906 21812 5918
rect 21756 5854 21758 5906
rect 21810 5854 21812 5906
rect 21644 5796 21700 5806
rect 21308 5794 21700 5796
rect 21308 5742 21646 5794
rect 21698 5742 21700 5794
rect 21308 5740 21700 5742
rect 21644 5730 21700 5740
rect 21756 5572 21812 5854
rect 21980 5908 22036 5918
rect 22204 5908 22260 6412
rect 22036 5852 22260 5908
rect 21980 5814 22036 5852
rect 21756 5506 21812 5516
rect 21420 5236 21476 5246
rect 21420 4340 21476 5180
rect 23212 5234 23268 6748
rect 23324 6580 23380 6972
rect 23548 6914 23604 6972
rect 23548 6862 23550 6914
rect 23602 6862 23604 6914
rect 23548 6850 23604 6862
rect 23324 6020 23380 6524
rect 23436 6690 23492 6702
rect 23436 6638 23438 6690
rect 23490 6638 23492 6690
rect 23436 6132 23492 6638
rect 23660 6468 23716 7310
rect 23660 6402 23716 6412
rect 23772 7252 23828 7532
rect 24108 7476 24164 7486
rect 24108 7382 24164 7420
rect 23660 6132 23716 6142
rect 23436 6130 23716 6132
rect 23436 6078 23662 6130
rect 23714 6078 23716 6130
rect 23436 6076 23716 6078
rect 23660 6066 23716 6076
rect 23772 6130 23828 7196
rect 23884 7250 23940 7262
rect 23884 7198 23886 7250
rect 23938 7198 23940 7250
rect 23884 6916 23940 7198
rect 23884 6850 23940 6860
rect 24108 6692 24164 6702
rect 24108 6598 24164 6636
rect 23884 6468 23940 6478
rect 23884 6374 23940 6412
rect 23772 6078 23774 6130
rect 23826 6078 23828 6130
rect 23772 6066 23828 6078
rect 24220 6356 24276 8372
rect 24332 8372 24724 8428
rect 24780 8372 24948 8428
rect 25452 8484 25508 8494
rect 24332 7474 24388 8372
rect 24780 7698 24836 8372
rect 24780 7646 24782 7698
rect 24834 7646 24836 7698
rect 24780 7634 24836 7646
rect 24332 7422 24334 7474
rect 24386 7422 24388 7474
rect 24332 7410 24388 7422
rect 24444 6916 24500 6926
rect 24332 6804 24388 6842
rect 24332 6738 24388 6748
rect 23324 5964 23604 6020
rect 23548 5906 23604 5964
rect 23548 5854 23550 5906
rect 23602 5854 23604 5906
rect 23548 5842 23604 5854
rect 24108 5908 24164 5918
rect 24220 5908 24276 6300
rect 24108 5906 24276 5908
rect 24108 5854 24110 5906
rect 24162 5854 24276 5906
rect 24108 5852 24276 5854
rect 24444 6690 24500 6860
rect 24444 6638 24446 6690
rect 24498 6638 24500 6690
rect 24444 6580 24500 6638
rect 25116 6690 25172 6702
rect 25116 6638 25118 6690
rect 25170 6638 25172 6690
rect 24780 6580 24836 6590
rect 24444 6578 24836 6580
rect 24444 6526 24782 6578
rect 24834 6526 24836 6578
rect 24444 6524 24836 6526
rect 24108 5842 24164 5852
rect 23212 5182 23214 5234
rect 23266 5182 23268 5234
rect 23212 5170 23268 5182
rect 23100 4900 23156 4910
rect 22316 4898 23156 4900
rect 22316 4846 23102 4898
rect 23154 4846 23156 4898
rect 22316 4844 23156 4846
rect 22316 4450 22372 4844
rect 23100 4834 23156 4844
rect 22316 4398 22318 4450
rect 22370 4398 22372 4450
rect 22316 4386 22372 4398
rect 21532 4340 21588 4350
rect 21420 4338 21588 4340
rect 21420 4286 21534 4338
rect 21586 4286 21588 4338
rect 21420 4284 21588 4286
rect 21196 4174 21198 4226
rect 21250 4174 21252 4226
rect 21196 4162 21252 4174
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 21532 3666 21588 4284
rect 24444 4226 24500 6524
rect 24780 6514 24836 6524
rect 25116 6244 25172 6638
rect 25452 6690 25508 8428
rect 26572 8484 26628 9772
rect 26348 8036 26404 8046
rect 26348 7474 26404 7980
rect 26348 7422 26350 7474
rect 26402 7422 26404 7474
rect 26348 7410 26404 7422
rect 26572 7474 26628 8428
rect 26684 9604 26740 10780
rect 26796 10834 26852 11230
rect 26796 10782 26798 10834
rect 26850 10782 26852 10834
rect 26796 10770 26852 10782
rect 26908 10500 26964 12684
rect 27020 12674 27076 12684
rect 27132 12404 27188 13692
rect 27132 12338 27188 12348
rect 27132 12180 27188 12190
rect 27020 12178 27188 12180
rect 27020 12126 27134 12178
rect 27186 12126 27188 12178
rect 27020 12124 27188 12126
rect 27020 10722 27076 12124
rect 27132 12114 27188 12124
rect 27244 11396 27300 14252
rect 27916 13860 27972 13870
rect 28028 13860 28084 16716
rect 28252 16706 28308 16716
rect 28812 16772 28868 16782
rect 28812 16678 28868 16716
rect 28140 15988 28196 15998
rect 28140 15894 28196 15932
rect 28364 15988 28420 15998
rect 28364 15894 28420 15932
rect 27916 13858 28084 13860
rect 27916 13806 27918 13858
rect 27970 13806 28084 13858
rect 27916 13804 28084 13806
rect 28476 14756 28532 14766
rect 27916 13794 27972 13804
rect 28476 12628 28532 14700
rect 28924 13972 28980 16830
rect 29148 16100 29204 17052
rect 29372 16884 29428 18620
rect 30492 17668 30548 19964
rect 30716 19906 30772 19918
rect 30716 19854 30718 19906
rect 30770 19854 30772 19906
rect 30604 19234 30660 19246
rect 30604 19182 30606 19234
rect 30658 19182 30660 19234
rect 30604 18676 30660 19182
rect 30716 19012 30772 19854
rect 30716 18946 30772 18956
rect 30940 19346 30996 20748
rect 31276 20580 31332 24556
rect 31388 24164 31444 24892
rect 32956 24722 33012 24734
rect 32956 24670 32958 24722
rect 33010 24670 33012 24722
rect 31836 24612 31892 24622
rect 31836 24518 31892 24556
rect 31500 24164 31556 24174
rect 31388 24162 31556 24164
rect 31388 24110 31502 24162
rect 31554 24110 31556 24162
rect 31388 24108 31556 24110
rect 31500 24098 31556 24108
rect 31612 23826 31668 23838
rect 31612 23774 31614 23826
rect 31666 23774 31668 23826
rect 31612 23716 31668 23774
rect 32060 23716 32116 23726
rect 31612 23714 32116 23716
rect 31612 23662 32062 23714
rect 32114 23662 32116 23714
rect 31612 23660 32116 23662
rect 31276 20514 31332 20524
rect 31388 20690 31444 20702
rect 31388 20638 31390 20690
rect 31442 20638 31444 20690
rect 31276 20244 31332 20254
rect 31388 20244 31444 20638
rect 31276 20242 31444 20244
rect 31276 20190 31278 20242
rect 31330 20190 31444 20242
rect 31276 20188 31444 20190
rect 31276 20178 31332 20188
rect 31612 20132 31668 20142
rect 31612 20038 31668 20076
rect 31052 20020 31108 20030
rect 31052 19926 31108 19964
rect 31388 20020 31444 20030
rect 31388 19926 31444 19964
rect 30940 19294 30942 19346
rect 30994 19294 30996 19346
rect 30604 18610 30660 18620
rect 30492 17574 30548 17612
rect 30828 18116 30884 18126
rect 30828 17780 30884 18060
rect 30828 17666 30884 17724
rect 30828 17614 30830 17666
rect 30882 17614 30884 17666
rect 30828 17602 30884 17614
rect 30716 17442 30772 17454
rect 30716 17390 30718 17442
rect 30770 17390 30772 17442
rect 29708 17108 29764 17118
rect 30716 17108 30772 17390
rect 29708 16884 29764 17052
rect 30380 17052 30772 17108
rect 30940 17108 30996 19294
rect 31500 19124 31556 19134
rect 30380 16994 30436 17052
rect 30940 17042 30996 17052
rect 31052 19012 31108 19022
rect 30380 16942 30382 16994
rect 30434 16942 30436 16994
rect 30380 16930 30436 16942
rect 29372 16882 29652 16884
rect 29372 16830 29374 16882
rect 29426 16830 29652 16882
rect 29372 16828 29652 16830
rect 29372 16818 29428 16828
rect 29260 16100 29316 16110
rect 29148 16098 29316 16100
rect 29148 16046 29262 16098
rect 29314 16046 29316 16098
rect 29148 16044 29316 16046
rect 29260 16034 29316 16044
rect 29372 15988 29428 15998
rect 29596 15988 29652 16828
rect 29708 16882 29988 16884
rect 29708 16830 29710 16882
rect 29762 16830 29988 16882
rect 29708 16828 29988 16830
rect 29708 16818 29764 16828
rect 29708 15988 29764 15998
rect 29596 15986 29764 15988
rect 29596 15934 29710 15986
rect 29762 15934 29764 15986
rect 29596 15932 29764 15934
rect 29372 15894 29428 15932
rect 29708 15922 29764 15932
rect 29484 15874 29540 15886
rect 29484 15822 29486 15874
rect 29538 15822 29540 15874
rect 29484 15202 29540 15822
rect 29484 15150 29486 15202
rect 29538 15150 29540 15202
rect 29484 15148 29540 15150
rect 29932 15538 29988 16828
rect 29932 15486 29934 15538
rect 29986 15486 29988 15538
rect 29484 15092 29652 15148
rect 28924 13906 28980 13916
rect 28476 12562 28532 12572
rect 29372 13860 29428 13870
rect 27580 12404 27636 12414
rect 27244 11330 27300 11340
rect 27356 12290 27412 12302
rect 27356 12238 27358 12290
rect 27410 12238 27412 12290
rect 27020 10670 27022 10722
rect 27074 10670 27076 10722
rect 27020 10658 27076 10670
rect 27132 10610 27188 10622
rect 27132 10558 27134 10610
rect 27186 10558 27188 10610
rect 27132 10500 27188 10558
rect 26908 10444 27300 10500
rect 26684 8428 26740 9548
rect 27020 9828 27076 9838
rect 27020 9602 27076 9772
rect 27020 9550 27022 9602
rect 27074 9550 27076 9602
rect 27020 9538 27076 9550
rect 27244 9380 27300 10444
rect 27356 10164 27412 12238
rect 27468 12178 27524 12190
rect 27468 12126 27470 12178
rect 27522 12126 27524 12178
rect 27468 12068 27524 12126
rect 27468 12002 27524 12012
rect 27580 11394 27636 12348
rect 28364 12404 28420 12414
rect 28364 12310 28420 12348
rect 27916 12068 27972 12078
rect 27916 11974 27972 12012
rect 29372 11508 29428 13804
rect 29484 13076 29540 13086
rect 29484 12962 29540 13020
rect 29484 12910 29486 12962
rect 29538 12910 29540 12962
rect 29484 12404 29540 12910
rect 29484 12338 29540 12348
rect 29372 11442 29428 11452
rect 27580 11342 27582 11394
rect 27634 11342 27636 11394
rect 27580 10724 27636 11342
rect 28252 11396 28308 11406
rect 28252 11302 28308 11340
rect 29260 11396 29316 11406
rect 29260 11302 29316 11340
rect 27580 10658 27636 10668
rect 27916 11170 27972 11182
rect 27916 11118 27918 11170
rect 27970 11118 27972 11170
rect 27580 10500 27636 10510
rect 27580 10498 27748 10500
rect 27580 10446 27582 10498
rect 27634 10446 27748 10498
rect 27580 10444 27748 10446
rect 27580 10434 27636 10444
rect 27356 9828 27412 10108
rect 27468 9828 27524 9838
rect 27356 9826 27524 9828
rect 27356 9774 27470 9826
rect 27522 9774 27524 9826
rect 27356 9772 27524 9774
rect 27468 9762 27524 9772
rect 27692 9716 27748 10444
rect 27692 9650 27748 9660
rect 27580 9604 27636 9614
rect 27580 9510 27636 9548
rect 27244 9324 27636 9380
rect 27580 9266 27636 9324
rect 27580 9214 27582 9266
rect 27634 9214 27636 9266
rect 27580 9202 27636 9214
rect 26684 8372 26964 8428
rect 26908 8260 26964 8372
rect 26908 8166 26964 8204
rect 27356 8260 27412 8270
rect 27356 8166 27412 8204
rect 26572 7422 26574 7474
rect 26626 7422 26628 7474
rect 26572 7410 26628 7422
rect 26684 8034 26740 8046
rect 26684 7982 26686 8034
rect 26738 7982 26740 8034
rect 26684 7588 26740 7982
rect 26796 8034 26852 8046
rect 26796 7982 26798 8034
rect 26850 7982 26852 8034
rect 26796 7812 26852 7982
rect 27916 7812 27972 11118
rect 28028 9828 28084 9838
rect 28028 9734 28084 9772
rect 28588 9716 28644 9726
rect 28588 9622 28644 9660
rect 29596 9492 29652 15092
rect 29932 13076 29988 15486
rect 30044 13972 30100 13982
rect 30044 13634 30100 13916
rect 30044 13582 30046 13634
rect 30098 13582 30100 13634
rect 30044 13570 30100 13582
rect 30156 13748 30212 13758
rect 29932 13010 29988 13020
rect 30156 12516 30212 13692
rect 30492 13636 30548 13646
rect 30268 12962 30324 12974
rect 30268 12910 30270 12962
rect 30322 12910 30324 12962
rect 30268 12852 30324 12910
rect 30380 12852 30436 12862
rect 30268 12796 30380 12852
rect 30380 12786 30436 12796
rect 30156 12450 30212 12460
rect 30380 12404 30436 12414
rect 30492 12404 30548 13580
rect 30436 12348 30548 12404
rect 30156 12180 30212 12190
rect 30156 12086 30212 12124
rect 30380 11172 30436 12348
rect 30828 12066 30884 12078
rect 30828 12014 30830 12066
rect 30882 12014 30884 12066
rect 30716 11172 30772 11182
rect 30828 11172 30884 12014
rect 30380 11170 30884 11172
rect 30380 11118 30718 11170
rect 30770 11118 30884 11170
rect 30380 11116 30884 11118
rect 30380 10612 30436 11116
rect 30716 11106 30772 11116
rect 30940 10612 30996 10622
rect 30268 10610 30436 10612
rect 30268 10558 30382 10610
rect 30434 10558 30436 10610
rect 30268 10556 30436 10558
rect 29708 10498 29764 10510
rect 29708 10446 29710 10498
rect 29762 10446 29764 10498
rect 29708 9940 29764 10446
rect 29708 9874 29764 9884
rect 29932 9716 29988 9726
rect 29932 9622 29988 9660
rect 30044 9604 30100 9614
rect 30044 9510 30100 9548
rect 29708 9492 29764 9502
rect 29596 9436 29708 9492
rect 29708 9426 29764 9436
rect 29820 8036 29876 8046
rect 28028 7812 28084 7822
rect 26796 7756 26964 7812
rect 27916 7756 28028 7812
rect 26796 7588 26852 7598
rect 26684 7586 26852 7588
rect 26684 7534 26798 7586
rect 26850 7534 26852 7586
rect 26684 7532 26852 7534
rect 25788 7252 25844 7262
rect 25788 7158 25844 7196
rect 26124 7250 26180 7262
rect 26124 7198 26126 7250
rect 26178 7198 26180 7250
rect 26124 7140 26180 7198
rect 26684 7140 26740 7532
rect 26796 7522 26852 7532
rect 26124 7084 26740 7140
rect 26796 7252 26852 7262
rect 26796 6914 26852 7196
rect 26796 6862 26798 6914
rect 26850 6862 26852 6914
rect 26796 6850 26852 6862
rect 26908 6914 26964 7756
rect 27020 7474 27076 7486
rect 27020 7422 27022 7474
rect 27074 7422 27076 7474
rect 27020 7364 27076 7422
rect 27244 7476 27300 7486
rect 27244 7382 27300 7420
rect 27020 7298 27076 7308
rect 27692 7364 27748 7374
rect 27692 7270 27748 7308
rect 26908 6862 26910 6914
rect 26962 6862 26964 6914
rect 26908 6850 26964 6862
rect 25452 6638 25454 6690
rect 25506 6638 25508 6690
rect 25452 6626 25508 6638
rect 25900 6802 25956 6814
rect 25900 6750 25902 6802
rect 25954 6750 25956 6802
rect 25228 6580 25284 6590
rect 25228 6486 25284 6524
rect 25116 6178 25172 6188
rect 25900 5234 25956 6750
rect 26236 6692 26292 6702
rect 26236 6598 26292 6636
rect 27244 6692 27300 6702
rect 26012 6578 26068 6590
rect 26012 6526 26014 6578
rect 26066 6526 26068 6578
rect 26012 6356 26068 6526
rect 26572 6580 26628 6590
rect 26572 6486 26628 6524
rect 27244 6578 27300 6636
rect 27580 6692 27636 6702
rect 28028 6692 28084 7756
rect 29820 7586 29876 7980
rect 30268 7812 30324 10556
rect 30380 10546 30436 10556
rect 30716 10610 30996 10612
rect 30716 10558 30942 10610
rect 30994 10558 30996 10610
rect 30716 10556 30996 10558
rect 30492 9940 30548 9950
rect 30492 9846 30548 9884
rect 30716 9714 30772 10556
rect 30940 10546 30996 10556
rect 31052 10052 31108 18956
rect 31388 18338 31444 18350
rect 31388 18286 31390 18338
rect 31442 18286 31444 18338
rect 31388 18116 31444 18286
rect 31388 18050 31444 18060
rect 31500 17666 31556 19068
rect 31500 17614 31502 17666
rect 31554 17614 31556 17666
rect 31500 17602 31556 17614
rect 31164 17556 31220 17566
rect 31164 17554 31332 17556
rect 31164 17502 31166 17554
rect 31218 17502 31332 17554
rect 31164 17500 31332 17502
rect 31164 17490 31220 17500
rect 31276 17444 31332 17500
rect 31612 17444 31668 17454
rect 31276 17442 31668 17444
rect 31276 17390 31614 17442
rect 31666 17390 31668 17442
rect 31276 17388 31668 17390
rect 31612 17378 31668 17388
rect 31724 17442 31780 17454
rect 31724 17390 31726 17442
rect 31778 17390 31780 17442
rect 31500 17220 31556 17230
rect 31500 15314 31556 17164
rect 31724 16772 31780 17390
rect 31724 16706 31780 16716
rect 31500 15262 31502 15314
rect 31554 15262 31556 15314
rect 31500 15250 31556 15262
rect 31724 15204 31780 15242
rect 31724 15138 31780 15148
rect 31500 12852 31556 12862
rect 31500 11170 31556 12796
rect 31612 12404 31668 12414
rect 31612 11394 31668 12348
rect 31836 11732 31892 23660
rect 32060 23650 32116 23660
rect 31948 22820 32004 22830
rect 31948 21700 32004 22764
rect 31948 20244 32004 21644
rect 31948 20178 32004 20188
rect 32060 20132 32116 20142
rect 32396 20132 32452 20142
rect 32060 20038 32116 20076
rect 32284 20130 32452 20132
rect 32284 20078 32398 20130
rect 32450 20078 32452 20130
rect 32284 20076 32452 20078
rect 31948 20018 32004 20030
rect 31948 19966 31950 20018
rect 32002 19966 32004 20018
rect 31948 19124 32004 19966
rect 31948 19058 32004 19068
rect 32172 20018 32228 20030
rect 32172 19966 32174 20018
rect 32226 19966 32228 20018
rect 32172 18452 32228 19966
rect 32172 18386 32228 18396
rect 32284 18340 32340 20076
rect 32396 20066 32452 20076
rect 32172 17668 32228 17678
rect 32284 17668 32340 18284
rect 32172 17666 32340 17668
rect 32172 17614 32174 17666
rect 32226 17614 32340 17666
rect 32172 17612 32340 17614
rect 32172 17602 32228 17612
rect 32508 16772 32564 16782
rect 32060 16100 32116 16110
rect 32060 16006 32116 16044
rect 32396 16098 32452 16110
rect 32396 16046 32398 16098
rect 32450 16046 32452 16098
rect 32396 15204 32452 16046
rect 32508 15876 32564 16716
rect 32508 15810 32564 15820
rect 32620 16098 32676 16110
rect 32620 16046 32622 16098
rect 32674 16046 32676 16098
rect 32396 15138 32452 15148
rect 32620 15764 32676 16046
rect 32060 15092 32116 15102
rect 32060 15090 32228 15092
rect 32060 15038 32062 15090
rect 32114 15038 32228 15090
rect 32060 15036 32228 15038
rect 32060 15026 32116 15036
rect 32060 13636 32116 13646
rect 32060 13542 32116 13580
rect 32172 13076 32228 15036
rect 32620 14644 32676 15708
rect 32956 15148 33012 24670
rect 33292 24722 33348 25452
rect 33292 24670 33294 24722
rect 33346 24670 33348 24722
rect 33292 24658 33348 24670
rect 33180 23380 33236 23390
rect 33068 23042 33124 23054
rect 33068 22990 33070 23042
rect 33122 22990 33124 23042
rect 33068 18788 33124 22990
rect 33180 22484 33236 23324
rect 33180 22390 33236 22428
rect 33068 16884 33124 18732
rect 33404 22148 33460 27804
rect 33516 25060 33572 41916
rect 33740 41860 33796 41870
rect 33740 41766 33796 41804
rect 33628 41300 33684 41310
rect 33628 41206 33684 41244
rect 33852 40964 33908 43484
rect 34076 42532 34132 42542
rect 33964 42530 34132 42532
rect 33964 42478 34078 42530
rect 34130 42478 34132 42530
rect 33964 42476 34132 42478
rect 33964 41860 34020 42476
rect 34076 42466 34132 42476
rect 34076 42196 34132 42206
rect 34076 42082 34132 42140
rect 34076 42030 34078 42082
rect 34130 42030 34132 42082
rect 34076 42018 34132 42030
rect 34412 41860 34468 41870
rect 33964 41858 34468 41860
rect 33964 41806 34414 41858
rect 34466 41806 34468 41858
rect 33964 41804 34468 41806
rect 33964 41748 34020 41804
rect 34412 41794 34468 41804
rect 33964 41682 34020 41692
rect 34636 41748 34692 41758
rect 34636 41746 34916 41748
rect 34636 41694 34638 41746
rect 34690 41694 34916 41746
rect 34636 41692 34916 41694
rect 34636 41682 34692 41692
rect 34076 41412 34132 41422
rect 33740 40908 33908 40964
rect 33964 41186 34020 41198
rect 33964 41134 33966 41186
rect 34018 41134 34020 41186
rect 33740 38668 33796 40908
rect 33740 38612 33908 38668
rect 33628 37266 33684 37278
rect 33628 37214 33630 37266
rect 33682 37214 33684 37266
rect 33628 37044 33684 37214
rect 33628 36978 33684 36988
rect 33628 35586 33684 35598
rect 33628 35534 33630 35586
rect 33682 35534 33684 35586
rect 33628 34132 33684 35534
rect 33852 34916 33908 38612
rect 33964 37940 34020 41134
rect 34076 40962 34132 41356
rect 34076 40910 34078 40962
rect 34130 40910 34132 40962
rect 34076 40898 34132 40910
rect 34524 41356 34804 41412
rect 34524 41188 34580 41356
rect 34524 40404 34580 41132
rect 34636 41186 34692 41198
rect 34636 41134 34638 41186
rect 34690 41134 34692 41186
rect 34636 40516 34692 41134
rect 34748 41186 34804 41356
rect 34860 41298 34916 41692
rect 34860 41246 34862 41298
rect 34914 41246 34916 41298
rect 34860 41234 34916 41246
rect 34748 41134 34750 41186
rect 34802 41134 34804 41186
rect 34748 41122 34804 41134
rect 35084 41188 35140 43708
rect 35644 43652 36036 43708
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35532 42084 35588 42094
rect 35532 41990 35588 42028
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35644 41412 35700 43652
rect 36652 43650 36708 43662
rect 36652 43598 36654 43650
rect 36706 43598 36708 43650
rect 36428 43316 36484 43326
rect 36428 42866 36484 43260
rect 36428 42814 36430 42866
rect 36482 42814 36484 42866
rect 36428 42802 36484 42814
rect 35420 41356 35700 41412
rect 35868 41972 35924 41982
rect 36652 41972 36708 43598
rect 35868 41970 36708 41972
rect 35868 41918 35870 41970
rect 35922 41918 36708 41970
rect 35868 41916 36708 41918
rect 36764 43652 36932 43708
rect 35084 41132 35252 41188
rect 34972 40962 35028 40974
rect 34972 40910 34974 40962
rect 35026 40910 35028 40962
rect 34860 40516 34916 40526
rect 34636 40514 34916 40516
rect 34636 40462 34862 40514
rect 34914 40462 34916 40514
rect 34636 40460 34916 40462
rect 34524 40402 34692 40404
rect 34524 40350 34526 40402
rect 34578 40350 34692 40402
rect 34524 40348 34692 40350
rect 34524 40338 34580 40348
rect 34636 39618 34692 40348
rect 34636 39566 34638 39618
rect 34690 39566 34692 39618
rect 34076 38834 34132 38846
rect 34076 38782 34078 38834
rect 34130 38782 34132 38834
rect 34076 38500 34132 38782
rect 34076 38434 34132 38444
rect 34300 38722 34356 38734
rect 34300 38670 34302 38722
rect 34354 38670 34356 38722
rect 33964 37874 34020 37884
rect 33852 34850 33908 34860
rect 33964 37604 34020 37614
rect 33964 34244 34020 37548
rect 34300 37268 34356 38670
rect 34300 37202 34356 37212
rect 34412 38050 34468 38062
rect 34412 37998 34414 38050
rect 34466 37998 34468 38050
rect 34076 37156 34132 37166
rect 34076 34354 34132 37100
rect 34412 37044 34468 37998
rect 34636 37380 34692 39566
rect 34860 39620 34916 40460
rect 34972 40516 35028 40910
rect 35084 40964 35140 40974
rect 35084 40870 35140 40908
rect 35196 40740 35252 41132
rect 34972 40450 35028 40460
rect 35084 40684 35252 40740
rect 34860 39618 35028 39620
rect 34860 39566 34862 39618
rect 34914 39566 35028 39618
rect 34860 39564 35028 39566
rect 34860 39554 34916 39564
rect 34636 37314 34692 37324
rect 34748 38834 34804 38846
rect 34748 38782 34750 38834
rect 34802 38782 34804 38834
rect 34748 38724 34804 38782
rect 34412 36978 34468 36988
rect 34188 35588 34244 35598
rect 34188 35494 34244 35532
rect 34748 35028 34804 38668
rect 34972 38722 35028 39564
rect 34972 38670 34974 38722
rect 35026 38670 35028 38722
rect 34972 38658 35028 38670
rect 35084 38276 35140 40684
rect 35420 40180 35476 41356
rect 35532 41186 35588 41198
rect 35532 41134 35534 41186
rect 35586 41134 35588 41186
rect 35532 40516 35588 41134
rect 35756 41186 35812 41198
rect 35756 41134 35758 41186
rect 35810 41134 35812 41186
rect 35644 40964 35700 40974
rect 35756 40964 35812 41134
rect 35700 40908 35812 40964
rect 35644 40898 35700 40908
rect 35644 40516 35700 40526
rect 35532 40460 35644 40516
rect 35644 40422 35700 40460
rect 35756 40402 35812 40908
rect 35756 40350 35758 40402
rect 35810 40350 35812 40402
rect 35756 40338 35812 40350
rect 35868 40290 35924 41916
rect 36652 41412 36708 41422
rect 36764 41412 36820 43652
rect 37100 43538 37156 43550
rect 37100 43486 37102 43538
rect 37154 43486 37156 43538
rect 37100 42978 37156 43486
rect 37100 42926 37102 42978
rect 37154 42926 37156 42978
rect 37100 42914 37156 42926
rect 37212 42642 37268 42654
rect 37212 42590 37214 42642
rect 37266 42590 37268 42642
rect 37100 42530 37156 42542
rect 37100 42478 37102 42530
rect 37154 42478 37156 42530
rect 36876 41972 36932 41982
rect 37100 41972 37156 42478
rect 36876 41970 37156 41972
rect 36876 41918 36878 41970
rect 36930 41918 37156 41970
rect 36876 41916 37156 41918
rect 36876 41860 36932 41916
rect 37212 41860 37268 42590
rect 37436 42532 37492 46620
rect 37548 46002 37604 46844
rect 38332 46834 38388 46844
rect 37548 45950 37550 46002
rect 37602 45950 37604 46002
rect 37548 45444 37604 45950
rect 37548 45378 37604 45388
rect 37660 46676 37716 46686
rect 37660 43762 37716 46620
rect 38892 46676 38948 46686
rect 39116 46676 39172 47294
rect 39900 46788 39956 46798
rect 39900 46694 39956 46732
rect 38948 46620 39172 46676
rect 38892 46582 38948 46620
rect 39564 46452 39620 46462
rect 39564 46002 39620 46396
rect 39564 45950 39566 46002
rect 39618 45950 39620 46002
rect 39564 45938 39620 45950
rect 37996 45890 38052 45902
rect 37996 45838 37998 45890
rect 38050 45838 38052 45890
rect 37996 45668 38052 45838
rect 38892 45890 38948 45902
rect 38892 45838 38894 45890
rect 38946 45838 38948 45890
rect 38052 45612 38500 45668
rect 37996 45602 38052 45612
rect 38332 45444 38388 45454
rect 37660 43710 37662 43762
rect 37714 43710 37716 43762
rect 37660 43698 37716 43710
rect 37884 44098 37940 44110
rect 37884 44046 37886 44098
rect 37938 44046 37940 44098
rect 37884 43708 37940 44046
rect 37884 43652 38164 43708
rect 37772 43538 37828 43550
rect 37772 43486 37774 43538
rect 37826 43486 37828 43538
rect 37772 42980 37828 43486
rect 37772 42914 37828 42924
rect 38108 43316 38164 43652
rect 38220 43426 38276 43438
rect 38220 43374 38222 43426
rect 38274 43374 38276 43426
rect 38220 43316 38276 43374
rect 38164 43260 38276 43316
rect 37772 42754 37828 42766
rect 37772 42702 37774 42754
rect 37826 42702 37828 42754
rect 37660 42532 37716 42542
rect 37436 42530 37716 42532
rect 37436 42478 37662 42530
rect 37714 42478 37716 42530
rect 37436 42476 37716 42478
rect 37660 42466 37716 42476
rect 36876 41794 36932 41804
rect 36988 41858 37268 41860
rect 36988 41806 37214 41858
rect 37266 41806 37268 41858
rect 36988 41804 37268 41806
rect 36708 41356 36820 41412
rect 36652 41346 36708 41356
rect 36988 41298 37044 41804
rect 37212 41794 37268 41804
rect 36988 41246 36990 41298
rect 37042 41246 37044 41298
rect 36988 41234 37044 41246
rect 36092 41188 36148 41198
rect 36092 41094 36148 41132
rect 37100 41186 37156 41198
rect 37100 41134 37102 41186
rect 37154 41134 37156 41186
rect 35868 40238 35870 40290
rect 35922 40238 35924 40290
rect 35868 40226 35924 40238
rect 35420 40124 35588 40180
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 39732 35252 39742
rect 35196 39638 35252 39676
rect 35532 38612 35588 40124
rect 37100 39732 37156 41134
rect 37436 41188 37492 41198
rect 37436 41094 37492 41132
rect 37100 38724 37156 39676
rect 37772 39060 37828 42702
rect 38108 42756 38164 43260
rect 38108 42754 38276 42756
rect 38108 42702 38110 42754
rect 38162 42702 38276 42754
rect 38108 42700 38276 42702
rect 38108 42690 38164 42700
rect 38220 41972 38276 42700
rect 38220 41906 38276 41916
rect 38108 41860 38164 41870
rect 38108 41766 38164 41804
rect 37660 39004 37828 39060
rect 37996 40402 38052 40414
rect 37996 40350 37998 40402
rect 38050 40350 38052 40402
rect 37548 38948 37604 38958
rect 37548 38854 37604 38892
rect 37660 38668 37716 39004
rect 37100 38658 37156 38668
rect 35532 38546 35588 38556
rect 37548 38612 37716 38668
rect 37884 38946 37940 38958
rect 37884 38894 37886 38946
rect 37938 38894 37940 38946
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34860 38220 35140 38276
rect 34860 37826 34916 38220
rect 36316 38164 36372 38174
rect 36316 38070 36372 38108
rect 37324 38164 37380 38174
rect 35308 38052 35364 38062
rect 35308 37958 35364 37996
rect 36540 38050 36596 38062
rect 36540 37998 36542 38050
rect 36594 37998 36596 38050
rect 34860 37774 34862 37826
rect 34914 37774 34916 37826
rect 34860 37762 34916 37774
rect 35084 37938 35140 37950
rect 35084 37886 35086 37938
rect 35138 37886 35140 37938
rect 35084 36708 35140 37886
rect 35644 37940 35700 37950
rect 35980 37940 36036 37950
rect 35644 37938 35924 37940
rect 35644 37886 35646 37938
rect 35698 37886 35924 37938
rect 35644 37884 35924 37886
rect 35644 37874 35700 37884
rect 35532 37826 35588 37838
rect 35532 37774 35534 37826
rect 35586 37774 35588 37826
rect 35532 37604 35588 37774
rect 35532 37538 35588 37548
rect 35756 37380 35812 37390
rect 35756 37286 35812 37324
rect 35644 37268 35700 37278
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 36652 35252 36708
rect 35196 36596 35252 36652
rect 35644 36706 35700 37212
rect 35644 36654 35646 36706
rect 35698 36654 35700 36706
rect 35644 36642 35700 36654
rect 35756 36932 35812 36942
rect 34972 35810 35028 35822
rect 34972 35758 34974 35810
rect 35026 35758 35028 35810
rect 34972 35588 35028 35758
rect 35196 35812 35252 36540
rect 35532 36594 35588 36606
rect 35532 36542 35534 36594
rect 35586 36542 35588 36594
rect 35420 36484 35476 36494
rect 35420 36390 35476 36428
rect 35196 35746 35252 35756
rect 35532 35700 35588 36542
rect 35532 35634 35588 35644
rect 34972 35364 35028 35532
rect 34972 35298 35028 35308
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35756 35252 35812 36876
rect 35196 35242 35460 35252
rect 34748 34962 34804 34972
rect 35644 35196 35812 35252
rect 34076 34302 34078 34354
rect 34130 34302 34132 34354
rect 34076 34290 34132 34302
rect 34972 34916 35028 34926
rect 34972 34802 35028 34860
rect 34972 34750 34974 34802
rect 35026 34750 35028 34802
rect 33628 33346 33684 34076
rect 33628 33294 33630 33346
rect 33682 33294 33684 33346
rect 33628 33282 33684 33294
rect 33740 34188 34020 34244
rect 33740 30212 33796 34188
rect 33964 34132 34020 34188
rect 34636 34244 34692 34254
rect 34636 34242 34804 34244
rect 34636 34190 34638 34242
rect 34690 34190 34804 34242
rect 34636 34188 34804 34190
rect 34636 34178 34692 34188
rect 34076 34132 34132 34142
rect 33964 34130 34132 34132
rect 33964 34078 34078 34130
rect 34130 34078 34132 34130
rect 33964 34076 34132 34078
rect 34076 34066 34132 34076
rect 33852 34018 33908 34030
rect 33852 33966 33854 34018
rect 33906 33966 33908 34018
rect 33852 33348 33908 33966
rect 34300 33348 34356 33358
rect 33852 33346 34356 33348
rect 33852 33294 34302 33346
rect 34354 33294 34356 33346
rect 33852 33292 34356 33294
rect 33852 31892 33908 33292
rect 34300 33282 34356 33292
rect 34524 33236 34580 33246
rect 34524 32564 34580 33180
rect 34748 32788 34804 34188
rect 34748 32722 34804 32732
rect 34860 33572 34916 33582
rect 33852 31826 33908 31836
rect 34300 32562 34804 32564
rect 34300 32510 34526 32562
rect 34578 32510 34804 32562
rect 34300 32508 34804 32510
rect 33740 30146 33796 30156
rect 34300 30210 34356 32508
rect 34524 32498 34580 32508
rect 34636 32116 34692 32126
rect 34524 31780 34580 31790
rect 34300 30158 34302 30210
rect 34354 30158 34356 30210
rect 34300 30146 34356 30158
rect 34412 31724 34524 31780
rect 34412 29652 34468 31724
rect 34524 31686 34580 31724
rect 34524 31556 34580 31566
rect 34524 31218 34580 31500
rect 34524 31166 34526 31218
rect 34578 31166 34580 31218
rect 34524 31154 34580 31166
rect 34636 30212 34692 32060
rect 34748 31890 34804 32508
rect 34860 32562 34916 33516
rect 34860 32510 34862 32562
rect 34914 32510 34916 32562
rect 34860 32498 34916 32510
rect 34748 31838 34750 31890
rect 34802 31838 34804 31890
rect 34748 31826 34804 31838
rect 34860 32340 34916 32350
rect 33852 29650 34468 29652
rect 33852 29598 34414 29650
rect 34466 29598 34468 29650
rect 33852 29596 34468 29598
rect 33852 27186 33908 29596
rect 34412 29586 34468 29596
rect 34524 30210 34692 30212
rect 34524 30158 34638 30210
rect 34690 30158 34692 30210
rect 34524 30156 34692 30158
rect 34524 29428 34580 30156
rect 34636 30146 34692 30156
rect 34748 29652 34804 29662
rect 34860 29652 34916 32284
rect 34804 29596 34916 29652
rect 34748 29558 34804 29596
rect 34076 29372 34580 29428
rect 34076 28754 34132 29372
rect 34076 28702 34078 28754
rect 34130 28702 34132 28754
rect 34076 28690 34132 28702
rect 34860 28642 34916 28654
rect 34860 28590 34862 28642
rect 34914 28590 34916 28642
rect 34524 27860 34580 27870
rect 34524 27766 34580 27804
rect 34860 27636 34916 28590
rect 34972 28084 35028 34750
rect 35084 34804 35140 34814
rect 35084 33908 35140 34748
rect 35084 33346 35140 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33294 35086 33346
rect 35138 33294 35140 33346
rect 35084 33282 35140 33294
rect 35084 32788 35140 32798
rect 35084 31556 35140 32732
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 31892 35252 31902
rect 35196 31778 35252 31836
rect 35196 31726 35198 31778
rect 35250 31726 35252 31778
rect 35196 31668 35252 31726
rect 35420 31780 35476 31790
rect 35420 31686 35476 31724
rect 35196 31602 35252 31612
rect 35084 31490 35140 31500
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 30322 35140 30334
rect 35084 30270 35086 30322
rect 35138 30270 35140 30322
rect 35084 30212 35140 30270
rect 35644 30212 35700 35196
rect 35756 35028 35812 35038
rect 35756 34934 35812 34972
rect 35868 34916 35924 37884
rect 35980 37846 36036 37884
rect 36204 37828 36260 37838
rect 36204 37268 36260 37772
rect 36204 37202 36260 37212
rect 36092 37044 36148 37054
rect 35980 35700 36036 35710
rect 35980 35606 36036 35644
rect 36092 35140 36148 36988
rect 36204 36820 36260 36830
rect 36204 36482 36260 36764
rect 36204 36430 36206 36482
rect 36258 36430 36260 36482
rect 36204 35364 36260 36430
rect 36540 35924 36596 37998
rect 36988 38052 37044 38062
rect 37100 38052 37156 38062
rect 37044 38050 37156 38052
rect 37044 37998 37102 38050
rect 37154 37998 37156 38050
rect 37044 37996 37156 37998
rect 36652 37268 36708 37278
rect 36708 37212 36820 37268
rect 36652 37174 36708 37212
rect 36540 35858 36596 35868
rect 36316 35812 36372 35822
rect 36316 35718 36372 35756
rect 36428 35698 36484 35710
rect 36428 35646 36430 35698
rect 36482 35646 36484 35698
rect 36428 35588 36484 35646
rect 36428 35522 36484 35532
rect 36652 35698 36708 35710
rect 36652 35646 36654 35698
rect 36706 35646 36708 35698
rect 36652 35476 36708 35646
rect 36652 35410 36708 35420
rect 36204 35298 36260 35308
rect 36092 35084 36372 35140
rect 36204 34916 36260 34926
rect 35868 34860 36204 34916
rect 36204 34822 36260 34860
rect 36092 34132 36148 34170
rect 35980 34076 36092 34132
rect 35756 32004 35812 32014
rect 35980 32004 36036 34076
rect 36092 34066 36148 34076
rect 36316 34130 36372 35084
rect 36316 34078 36318 34130
rect 36370 34078 36372 34130
rect 36092 33908 36148 33918
rect 36092 33814 36148 33852
rect 35756 32002 36036 32004
rect 35756 31950 35758 32002
rect 35810 31950 36036 32002
rect 35756 31948 36036 31950
rect 36204 33122 36260 33134
rect 36204 33070 36206 33122
rect 36258 33070 36260 33122
rect 35756 31938 35812 31948
rect 36204 31556 36260 33070
rect 36316 32450 36372 34078
rect 36652 34020 36708 34030
rect 36764 34020 36820 37212
rect 36876 36708 36932 36718
rect 36876 36614 36932 36652
rect 36988 36484 37044 37996
rect 37100 37986 37156 37996
rect 37324 37938 37380 38108
rect 37324 37886 37326 37938
rect 37378 37886 37380 37938
rect 37100 37492 37156 37530
rect 37100 37426 37156 37436
rect 37212 37378 37268 37390
rect 37212 37326 37214 37378
rect 37266 37326 37268 37378
rect 37100 37266 37156 37278
rect 37100 37214 37102 37266
rect 37154 37214 37156 37266
rect 37100 36820 37156 37214
rect 37100 36754 37156 36764
rect 37100 36484 37156 36494
rect 36988 36482 37156 36484
rect 36988 36430 37102 36482
rect 37154 36430 37156 36482
rect 36988 36428 37156 36430
rect 37100 36418 37156 36428
rect 37212 36484 37268 37326
rect 36708 33964 36820 34020
rect 36988 35364 37044 35374
rect 36988 34802 37044 35308
rect 37212 35028 37268 36428
rect 37324 36372 37380 37886
rect 37548 36708 37604 38612
rect 37884 38164 37940 38894
rect 37996 38948 38052 40350
rect 37996 38882 38052 38892
rect 38108 40290 38164 40302
rect 38108 40238 38110 40290
rect 38162 40238 38164 40290
rect 38108 39620 38164 40238
rect 38108 38164 38164 39564
rect 38332 38668 38388 45388
rect 38444 45330 38500 45612
rect 38444 45278 38446 45330
rect 38498 45278 38500 45330
rect 38444 45266 38500 45278
rect 38892 45332 38948 45838
rect 40572 45332 40628 52668
rect 41692 52500 41748 53564
rect 41580 52444 41748 52500
rect 42476 52946 42532 54012
rect 44268 54068 44324 55022
rect 45948 55020 46340 55076
rect 42476 52894 42478 52946
rect 42530 52894 42532 52946
rect 41020 51490 41076 51502
rect 41020 51438 41022 51490
rect 41074 51438 41076 51490
rect 40908 51156 40964 51166
rect 40684 51154 40964 51156
rect 40684 51102 40910 51154
rect 40962 51102 40964 51154
rect 40684 51100 40964 51102
rect 40684 50706 40740 51100
rect 40908 51090 40964 51100
rect 41020 50820 41076 51438
rect 41580 51490 41636 52444
rect 42476 51604 42532 52894
rect 43148 53956 43204 53966
rect 43148 52052 43204 53900
rect 44268 53732 44324 54012
rect 44268 53666 44324 53676
rect 45500 54740 45556 54750
rect 45948 54740 46004 55020
rect 45500 54738 46004 54740
rect 45500 54686 45502 54738
rect 45554 54686 45950 54738
rect 46002 54686 46004 54738
rect 45500 54684 46004 54686
rect 45500 53620 45556 54684
rect 45948 54674 46004 54684
rect 46620 54738 46676 55916
rect 46732 55412 46788 56252
rect 46956 56242 47012 56252
rect 47628 56242 47684 56252
rect 47964 56308 48020 56318
rect 47068 56082 47124 56094
rect 47068 56030 47070 56082
rect 47122 56030 47124 56082
rect 47068 55636 47124 56030
rect 46732 55346 46788 55356
rect 46844 55580 47124 55636
rect 47180 56082 47236 56094
rect 47180 56030 47182 56082
rect 47234 56030 47236 56082
rect 46620 54686 46622 54738
rect 46674 54686 46676 54738
rect 46620 54674 46676 54686
rect 46060 54628 46116 54638
rect 46060 54514 46116 54572
rect 46844 54628 46900 55580
rect 47180 55524 47236 56030
rect 46844 54562 46900 54572
rect 46956 55468 47236 55524
rect 47628 56082 47684 56094
rect 47628 56030 47630 56082
rect 47682 56030 47684 56082
rect 46956 55188 47012 55468
rect 47628 55412 47684 56030
rect 47852 55970 47908 55982
rect 47852 55918 47854 55970
rect 47906 55918 47908 55970
rect 47740 55412 47796 55422
rect 47628 55410 47796 55412
rect 47628 55358 47742 55410
rect 47794 55358 47796 55410
rect 47628 55356 47796 55358
rect 46060 54462 46062 54514
rect 46114 54462 46116 54514
rect 45500 53554 45556 53564
rect 45836 53732 45892 53742
rect 45836 53170 45892 53676
rect 45836 53118 45838 53170
rect 45890 53118 45892 53170
rect 45836 53106 45892 53118
rect 43260 52834 43316 52846
rect 43260 52782 43262 52834
rect 43314 52782 43316 52834
rect 43260 52274 43316 52782
rect 43260 52222 43262 52274
rect 43314 52222 43316 52274
rect 43260 52210 43316 52222
rect 43820 52836 43876 52846
rect 43820 52162 43876 52780
rect 45388 52834 45444 52846
rect 45388 52782 45390 52834
rect 45442 52782 45444 52834
rect 45388 52724 45444 52782
rect 45612 52724 45668 52734
rect 45388 52722 45668 52724
rect 45388 52670 45614 52722
rect 45666 52670 45668 52722
rect 45388 52668 45668 52670
rect 45612 52658 45668 52668
rect 43820 52110 43822 52162
rect 43874 52110 43876 52162
rect 43820 52098 43876 52110
rect 45500 52276 45556 52286
rect 43148 51958 43204 51996
rect 44156 52052 44212 52062
rect 43372 51938 43428 51950
rect 43372 51886 43374 51938
rect 43426 51886 43428 51938
rect 42476 51538 42532 51548
rect 43260 51604 43316 51614
rect 43260 51510 43316 51548
rect 41580 51438 41582 51490
rect 41634 51438 41636 51490
rect 41580 51380 41636 51438
rect 41692 51492 41748 51502
rect 41692 51490 41860 51492
rect 41692 51438 41694 51490
rect 41746 51438 41860 51490
rect 41692 51436 41860 51438
rect 41692 51426 41748 51436
rect 41020 50754 41076 50764
rect 41132 51324 41636 51380
rect 40684 50654 40686 50706
rect 40738 50654 40740 50706
rect 40684 50642 40740 50654
rect 41132 50428 41188 51324
rect 41804 51268 41860 51436
rect 43260 51380 43316 51390
rect 41244 51212 41636 51268
rect 41244 51154 41300 51212
rect 41244 51102 41246 51154
rect 41298 51102 41300 51154
rect 41244 51090 41300 51102
rect 41580 51156 41636 51212
rect 41804 51202 41860 51212
rect 42252 51268 42308 51278
rect 42252 51174 42308 51212
rect 41692 51156 41748 51166
rect 41580 51154 41748 51156
rect 41580 51102 41694 51154
rect 41746 51102 41748 51154
rect 41580 51100 41748 51102
rect 41692 51090 41748 51100
rect 41804 50820 41860 50830
rect 41804 50726 41860 50764
rect 41468 50596 41524 50606
rect 41468 50502 41524 50540
rect 41916 50594 41972 50606
rect 41916 50542 41918 50594
rect 41970 50542 41972 50594
rect 41916 50428 41972 50542
rect 41132 50372 41412 50428
rect 41020 50036 41076 50046
rect 41020 49942 41076 49980
rect 41244 49810 41300 49822
rect 41244 49758 41246 49810
rect 41298 49758 41300 49810
rect 41244 49588 41300 49758
rect 41356 49810 41412 50372
rect 41804 50372 41972 50428
rect 42140 50594 42196 50606
rect 42140 50542 42142 50594
rect 42194 50542 42196 50594
rect 41356 49758 41358 49810
rect 41410 49758 41412 49810
rect 41356 49746 41412 49758
rect 41468 49812 41524 49822
rect 41468 49718 41524 49756
rect 41804 49698 41860 50372
rect 42140 50036 42196 50542
rect 42140 49970 42196 49980
rect 42252 50594 42308 50606
rect 42252 50542 42254 50594
rect 42306 50542 42308 50594
rect 41804 49646 41806 49698
rect 41858 49646 41860 49698
rect 41804 49588 41860 49646
rect 41244 49532 41860 49588
rect 41916 49922 41972 49934
rect 41916 49870 41918 49922
rect 41970 49870 41972 49922
rect 41916 49028 41972 49870
rect 42252 49812 42308 50542
rect 42812 50596 42868 50606
rect 42812 50428 42868 50540
rect 42812 50372 42980 50428
rect 42140 49700 42196 49710
rect 41692 49026 41972 49028
rect 41692 48974 41918 49026
rect 41970 48974 41972 49026
rect 41692 48972 41972 48974
rect 41692 48466 41748 48972
rect 41916 48962 41972 48972
rect 42028 49644 42140 49700
rect 42028 49026 42084 49644
rect 42140 49606 42196 49644
rect 42252 49364 42308 49756
rect 42140 49308 42308 49364
rect 42140 49138 42196 49308
rect 42140 49086 42142 49138
rect 42194 49086 42196 49138
rect 42140 49074 42196 49086
rect 42028 48974 42030 49026
rect 42082 48974 42084 49026
rect 41692 48414 41694 48466
rect 41746 48414 41748 48466
rect 41692 48402 41748 48414
rect 41580 48132 41636 48142
rect 41356 47234 41412 47246
rect 41356 47182 41358 47234
rect 41410 47182 41412 47234
rect 41020 46786 41076 46798
rect 41020 46734 41022 46786
rect 41074 46734 41076 46786
rect 40908 46452 40964 46462
rect 41020 46452 41076 46734
rect 41244 46788 41300 46798
rect 41356 46788 41412 47182
rect 41244 46786 41412 46788
rect 41244 46734 41246 46786
rect 41298 46734 41412 46786
rect 41244 46732 41412 46734
rect 41244 46722 41300 46732
rect 41468 46452 41524 46462
rect 41020 46450 41524 46452
rect 41020 46398 41470 46450
rect 41522 46398 41524 46450
rect 41020 46396 41524 46398
rect 40908 46358 40964 46396
rect 41468 46386 41524 46396
rect 41580 46004 41636 48076
rect 41692 47572 41748 47582
rect 41692 47460 41748 47516
rect 42028 47460 42084 48974
rect 42252 49028 42308 49038
rect 42812 49028 42868 49038
rect 42252 49026 42868 49028
rect 42252 48974 42254 49026
rect 42306 48974 42814 49026
rect 42866 48974 42868 49026
rect 42252 48972 42868 48974
rect 42252 48962 42308 48972
rect 42364 48802 42420 48814
rect 42364 48750 42366 48802
rect 42418 48750 42420 48802
rect 42364 48356 42420 48750
rect 42476 48466 42532 48972
rect 42812 48962 42868 48972
rect 42476 48414 42478 48466
rect 42530 48414 42532 48466
rect 42476 48402 42532 48414
rect 42364 48262 42420 48300
rect 42588 48132 42644 48142
rect 42476 48018 42532 48030
rect 42476 47966 42478 48018
rect 42530 47966 42532 48018
rect 41692 47458 42084 47460
rect 41692 47406 41694 47458
rect 41746 47406 42084 47458
rect 41692 47404 42084 47406
rect 42140 47572 42196 47582
rect 41692 47394 41748 47404
rect 41692 46564 41748 46574
rect 41692 46562 41860 46564
rect 41692 46510 41694 46562
rect 41746 46510 41860 46562
rect 41692 46508 41860 46510
rect 41692 46498 41748 46508
rect 41804 46450 41860 46508
rect 41804 46398 41806 46450
rect 41858 46398 41860 46450
rect 41692 46004 41748 46014
rect 41580 46002 41748 46004
rect 41580 45950 41694 46002
rect 41746 45950 41748 46002
rect 41580 45948 41748 45950
rect 41692 45938 41748 45948
rect 40684 45332 40740 45342
rect 40572 45276 40684 45332
rect 38892 44324 38948 45276
rect 40684 45266 40740 45276
rect 40236 44884 40292 44894
rect 38892 44258 38948 44268
rect 39116 44436 39172 44446
rect 38556 43650 38612 43662
rect 38556 43598 38558 43650
rect 38610 43598 38612 43650
rect 38556 42642 38612 43598
rect 38556 42590 38558 42642
rect 38610 42590 38612 42642
rect 38444 41972 38500 41982
rect 38556 41972 38612 42590
rect 39004 42980 39060 42990
rect 38780 41972 38836 41982
rect 38556 41970 38836 41972
rect 38556 41918 38782 41970
rect 38834 41918 38836 41970
rect 38556 41916 38836 41918
rect 38444 41300 38500 41916
rect 38556 41300 38612 41310
rect 38444 41298 38612 41300
rect 38444 41246 38558 41298
rect 38610 41246 38612 41298
rect 38444 41244 38612 41246
rect 38556 41234 38612 41244
rect 38780 40514 38836 41916
rect 38892 41972 38948 41982
rect 38892 41858 38948 41916
rect 38892 41806 38894 41858
rect 38946 41806 38948 41858
rect 38892 41794 38948 41806
rect 39004 41746 39060 42924
rect 39004 41694 39006 41746
rect 39058 41694 39060 41746
rect 39004 41682 39060 41694
rect 38780 40462 38782 40514
rect 38834 40462 38836 40514
rect 38780 40450 38836 40462
rect 39116 38948 39172 44380
rect 39676 43538 39732 43550
rect 39676 43486 39678 43538
rect 39730 43486 39732 43538
rect 39340 42756 39396 42766
rect 39676 42756 39732 43486
rect 40236 42866 40292 44828
rect 40796 44324 40852 44334
rect 40796 44230 40852 44268
rect 41468 44210 41524 44222
rect 41468 44158 41470 44210
rect 41522 44158 41524 44210
rect 41468 43708 41524 44158
rect 41804 43708 41860 46398
rect 42140 46002 42196 47516
rect 42476 47458 42532 47966
rect 42476 47406 42478 47458
rect 42530 47406 42532 47458
rect 42476 47394 42532 47406
rect 42588 47346 42644 48076
rect 42588 47294 42590 47346
rect 42642 47294 42644 47346
rect 42588 47282 42644 47294
rect 42700 47908 42756 47918
rect 42140 45950 42142 46002
rect 42194 45950 42196 46002
rect 41356 43652 41524 43708
rect 41580 43652 41860 43708
rect 41916 45332 41972 45342
rect 41020 43540 41076 43550
rect 41020 43446 41076 43484
rect 40348 43428 40404 43438
rect 40348 43334 40404 43372
rect 40236 42814 40238 42866
rect 40290 42814 40292 42866
rect 40236 42802 40292 42814
rect 40796 42980 40852 42990
rect 39340 42754 39732 42756
rect 39340 42702 39342 42754
rect 39394 42702 39732 42754
rect 39340 42700 39732 42702
rect 39788 42754 39844 42766
rect 39788 42702 39790 42754
rect 39842 42702 39844 42754
rect 39340 42084 39396 42700
rect 39788 42644 39844 42702
rect 40796 42754 40852 42924
rect 41356 42978 41412 43652
rect 41468 43540 41524 43550
rect 41468 43446 41524 43484
rect 41356 42926 41358 42978
rect 41410 42926 41412 42978
rect 41356 42914 41412 42926
rect 40796 42702 40798 42754
rect 40850 42702 40852 42754
rect 40796 42690 40852 42702
rect 39788 42578 39844 42588
rect 40572 42644 40628 42654
rect 40572 42550 40628 42588
rect 41468 42532 41524 42542
rect 41580 42532 41636 43652
rect 41692 42644 41748 42654
rect 41692 42550 41748 42588
rect 41468 42530 41636 42532
rect 41468 42478 41470 42530
rect 41522 42478 41636 42530
rect 41468 42476 41636 42478
rect 41468 42466 41524 42476
rect 39340 42018 39396 42028
rect 39452 42420 39508 42430
rect 39116 38892 39396 38948
rect 39228 38722 39284 38734
rect 39228 38670 39230 38722
rect 39282 38670 39284 38722
rect 38332 38612 38500 38668
rect 38332 38164 38388 38174
rect 38108 38162 38388 38164
rect 38108 38110 38334 38162
rect 38386 38110 38388 38162
rect 38108 38108 38388 38110
rect 37548 36642 37604 36652
rect 37660 37938 37716 37950
rect 37660 37886 37662 37938
rect 37714 37886 37716 37938
rect 37660 36482 37716 37886
rect 37772 37604 37828 37614
rect 37772 37378 37828 37548
rect 37772 37326 37774 37378
rect 37826 37326 37828 37378
rect 37772 37314 37828 37326
rect 37884 36594 37940 38108
rect 38332 38098 38388 38108
rect 37884 36542 37886 36594
rect 37938 36542 37940 36594
rect 37884 36530 37940 36542
rect 37660 36430 37662 36482
rect 37714 36430 37716 36482
rect 37436 36372 37492 36382
rect 37324 36370 37492 36372
rect 37324 36318 37438 36370
rect 37490 36318 37492 36370
rect 37324 36316 37492 36318
rect 37436 36306 37492 36316
rect 37660 36148 37716 36430
rect 37548 36092 37716 36148
rect 38332 36484 38388 36494
rect 37324 35924 37380 35934
rect 37324 35830 37380 35868
rect 37436 35810 37492 35822
rect 37436 35758 37438 35810
rect 37490 35758 37492 35810
rect 37436 35700 37492 35758
rect 37212 34972 37380 35028
rect 36988 34750 36990 34802
rect 37042 34750 37044 34802
rect 36652 33954 36708 33964
rect 36988 33908 37044 34750
rect 37212 34692 37268 34702
rect 37324 34692 37380 34972
rect 37436 34916 37492 35644
rect 37548 35138 37604 36092
rect 38332 35924 38388 36428
rect 38332 35830 38388 35868
rect 37548 35086 37550 35138
rect 37602 35086 37604 35138
rect 37548 35074 37604 35086
rect 37660 35698 37716 35710
rect 37660 35646 37662 35698
rect 37714 35646 37716 35698
rect 37436 34860 37604 34916
rect 37436 34692 37492 34702
rect 37324 34690 37492 34692
rect 37324 34638 37438 34690
rect 37490 34638 37492 34690
rect 37324 34636 37492 34638
rect 37100 34132 37156 34142
rect 37100 34038 37156 34076
rect 36988 33852 37156 33908
rect 36316 32398 36318 32450
rect 36370 32398 36372 32450
rect 36316 32386 36372 32398
rect 36988 33346 37044 33358
rect 36988 33294 36990 33346
rect 37042 33294 37044 33346
rect 36988 32004 37044 33294
rect 37100 32452 37156 33852
rect 37212 32788 37268 34636
rect 37436 34626 37492 34636
rect 37548 33572 37604 34860
rect 37660 34692 37716 35646
rect 37996 35700 38052 35710
rect 37884 35026 37940 35038
rect 37884 34974 37886 35026
rect 37938 34974 37940 35026
rect 37884 34916 37940 34974
rect 37884 34850 37940 34860
rect 37660 34626 37716 34636
rect 37884 34690 37940 34702
rect 37884 34638 37886 34690
rect 37938 34638 37940 34690
rect 37660 34020 37716 34030
rect 37660 33926 37716 33964
rect 37548 33478 37604 33516
rect 37212 32732 37380 32788
rect 37212 32564 37268 32602
rect 37212 32498 37268 32508
rect 37100 32386 37156 32396
rect 37212 32340 37268 32350
rect 37324 32340 37380 32732
rect 37660 32452 37716 32462
rect 37660 32358 37716 32396
rect 37268 32284 37380 32340
rect 37212 32274 37268 32284
rect 37884 32004 37940 34638
rect 37996 32564 38052 35644
rect 38108 35588 38164 35598
rect 38108 35138 38164 35532
rect 38220 35586 38276 35598
rect 38220 35534 38222 35586
rect 38274 35534 38276 35586
rect 38220 35476 38276 35534
rect 38220 35410 38276 35420
rect 38108 35086 38110 35138
rect 38162 35086 38164 35138
rect 38108 35074 38164 35086
rect 38108 33572 38164 33582
rect 38444 33572 38500 38612
rect 38780 38164 38836 38174
rect 38668 37940 38724 37950
rect 38668 35924 38724 37884
rect 38780 37380 38836 38108
rect 39004 37940 39060 37950
rect 38780 37044 38836 37324
rect 38892 37938 39060 37940
rect 38892 37886 39006 37938
rect 39058 37886 39060 37938
rect 38892 37884 39060 37886
rect 38892 37268 38948 37884
rect 39004 37874 39060 37884
rect 39228 37716 39284 38670
rect 39004 37660 39284 37716
rect 39004 37490 39060 37660
rect 39004 37438 39006 37490
rect 39058 37438 39060 37490
rect 39004 37426 39060 37438
rect 39228 37268 39284 37278
rect 38892 37266 39284 37268
rect 38892 37214 39230 37266
rect 39282 37214 39284 37266
rect 38892 37212 39284 37214
rect 39228 37156 39284 37212
rect 39228 37090 39284 37100
rect 38892 37044 38948 37054
rect 38780 37042 38948 37044
rect 38780 36990 38894 37042
rect 38946 36990 38948 37042
rect 38780 36988 38948 36990
rect 38892 36978 38948 36988
rect 38780 35924 38836 35934
rect 38668 35922 38836 35924
rect 38668 35870 38782 35922
rect 38834 35870 38836 35922
rect 38668 35868 38836 35870
rect 38780 35858 38836 35868
rect 39004 35924 39060 35934
rect 39004 35830 39060 35868
rect 39116 35700 39172 35710
rect 39116 35606 39172 35644
rect 38108 33458 38164 33516
rect 38108 33406 38110 33458
rect 38162 33406 38164 33458
rect 38108 33394 38164 33406
rect 38220 33516 38500 33572
rect 38556 35588 38612 35598
rect 38556 33572 38612 35532
rect 38780 35028 38836 35038
rect 38668 34692 38724 34702
rect 38668 34598 38724 34636
rect 38780 34018 38836 34972
rect 39340 35028 39396 38892
rect 39452 38946 39508 42364
rect 41132 41972 41188 41982
rect 41020 41970 41188 41972
rect 41020 41918 41134 41970
rect 41186 41918 41188 41970
rect 41020 41916 41188 41918
rect 40348 41858 40404 41870
rect 40348 41806 40350 41858
rect 40402 41806 40404 41858
rect 40348 41748 40404 41806
rect 40348 41682 40404 41692
rect 40124 41300 40180 41310
rect 40124 41298 40292 41300
rect 40124 41246 40126 41298
rect 40178 41246 40292 41298
rect 40124 41244 40292 41246
rect 40124 41234 40180 41244
rect 40236 40514 40292 41244
rect 40236 40462 40238 40514
rect 40290 40462 40292 40514
rect 40236 40404 40292 40462
rect 40348 41188 40404 41198
rect 40348 40516 40404 41132
rect 41020 40516 41076 41916
rect 41132 41906 41188 41916
rect 41356 41972 41412 41982
rect 41356 41970 41524 41972
rect 41356 41918 41358 41970
rect 41410 41918 41524 41970
rect 41356 41916 41524 41918
rect 41356 41906 41412 41916
rect 41244 41858 41300 41870
rect 41244 41806 41246 41858
rect 41298 41806 41300 41858
rect 41132 41076 41188 41086
rect 41132 40626 41188 41020
rect 41132 40574 41134 40626
rect 41186 40574 41188 40626
rect 41132 40562 41188 40574
rect 41244 40628 41300 41806
rect 41244 40572 41412 40628
rect 40348 40514 41076 40516
rect 40348 40462 40350 40514
rect 40402 40462 41076 40514
rect 40348 40460 41076 40462
rect 40348 40450 40404 40460
rect 40236 40338 40292 40348
rect 40796 40402 40852 40460
rect 40796 40350 40798 40402
rect 40850 40350 40852 40402
rect 40796 40338 40852 40350
rect 41244 40404 41300 40414
rect 41244 40310 41300 40348
rect 41356 40402 41412 40572
rect 41356 40350 41358 40402
rect 41410 40350 41412 40402
rect 41356 40338 41412 40350
rect 41468 40404 41524 41916
rect 41580 40404 41636 42476
rect 41692 41970 41748 41982
rect 41692 41918 41694 41970
rect 41746 41918 41748 41970
rect 41692 41748 41748 41918
rect 41748 41692 41860 41748
rect 41692 41682 41748 41692
rect 41692 40404 41748 40414
rect 41580 40348 41692 40404
rect 41468 40338 41524 40348
rect 40236 40178 40292 40190
rect 40236 40126 40238 40178
rect 40290 40126 40292 40178
rect 39452 38894 39454 38946
rect 39506 38894 39508 38946
rect 39452 38882 39508 38894
rect 39788 39508 39844 39518
rect 39676 38834 39732 38846
rect 39676 38782 39678 38834
rect 39730 38782 39732 38834
rect 39676 38612 39732 38782
rect 39676 38546 39732 38556
rect 39564 37380 39620 37390
rect 39564 37286 39620 37324
rect 39676 37378 39732 37390
rect 39676 37326 39678 37378
rect 39730 37326 39732 37378
rect 39676 37156 39732 37326
rect 39676 37090 39732 37100
rect 39340 34962 39396 34972
rect 38780 33966 38782 34018
rect 38834 33966 38836 34018
rect 38780 33954 38836 33966
rect 39116 34804 39172 34814
rect 38556 33516 38724 33572
rect 37996 32470 38052 32508
rect 38220 32116 38276 33516
rect 38444 33348 38500 33358
rect 36988 31938 37044 31948
rect 37772 31948 37940 32004
rect 38108 32060 38276 32116
rect 38332 33346 38500 33348
rect 38332 33294 38446 33346
rect 38498 33294 38500 33346
rect 38332 33292 38500 33294
rect 36204 31490 36260 31500
rect 37100 31890 37156 31902
rect 37100 31838 37102 31890
rect 37154 31838 37156 31890
rect 37100 31556 37156 31838
rect 37772 31892 37828 31948
rect 37772 31826 37828 31836
rect 37436 31780 37492 31790
rect 37436 31686 37492 31724
rect 37884 31780 37940 31790
rect 37884 31686 37940 31724
rect 37100 31490 37156 31500
rect 35756 30212 35812 30222
rect 35084 30146 35140 30156
rect 35308 30210 35812 30212
rect 35308 30158 35758 30210
rect 35810 30158 35812 30210
rect 35308 30156 35812 30158
rect 35308 29650 35364 30156
rect 35756 30146 35812 30156
rect 37100 30212 37156 30222
rect 37100 30118 37156 30156
rect 37772 30100 37828 30110
rect 37212 30098 37828 30100
rect 37212 30046 37774 30098
rect 37826 30046 37828 30098
rect 37212 30044 37828 30046
rect 35308 29598 35310 29650
rect 35362 29598 35364 29650
rect 35308 29586 35364 29598
rect 35532 29986 35588 29998
rect 35532 29934 35534 29986
rect 35586 29934 35588 29986
rect 35532 29428 35588 29934
rect 36540 29986 36596 29998
rect 36540 29934 36542 29986
rect 36594 29934 36596 29986
rect 35644 29428 35700 29438
rect 35532 29426 35700 29428
rect 35532 29374 35646 29426
rect 35698 29374 35700 29426
rect 35532 29372 35700 29374
rect 34972 28018 35028 28028
rect 35084 29204 35140 29214
rect 35084 28644 35140 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28082 35140 28588
rect 35308 28868 35364 28878
rect 35308 28644 35364 28812
rect 35644 28644 35700 29372
rect 35980 29314 36036 29326
rect 35980 29262 35982 29314
rect 36034 29262 36036 29314
rect 35980 28868 36036 29262
rect 36540 29316 36596 29934
rect 37212 29650 37268 30044
rect 37772 30034 37828 30044
rect 37212 29598 37214 29650
rect 37266 29598 37268 29650
rect 37212 29586 37268 29598
rect 37772 29876 37828 29886
rect 36876 29428 36932 29438
rect 36876 29334 36932 29372
rect 36988 29426 37044 29438
rect 36988 29374 36990 29426
rect 37042 29374 37044 29426
rect 36540 29092 36596 29260
rect 36988 29092 37044 29374
rect 36540 29036 37044 29092
rect 37436 29426 37492 29438
rect 37436 29374 37438 29426
rect 37490 29374 37492 29426
rect 35980 28802 36036 28812
rect 35868 28644 35924 28654
rect 35308 28642 35588 28644
rect 35308 28590 35310 28642
rect 35362 28590 35588 28642
rect 35308 28588 35588 28590
rect 35644 28642 35924 28644
rect 35644 28590 35870 28642
rect 35922 28590 35924 28642
rect 35644 28588 35924 28590
rect 35308 28578 35364 28588
rect 35532 28532 35588 28588
rect 35532 28476 35812 28532
rect 35084 28030 35086 28082
rect 35138 28030 35140 28082
rect 35084 28018 35140 28030
rect 35756 28082 35812 28476
rect 35756 28030 35758 28082
rect 35810 28030 35812 28082
rect 35756 28018 35812 28030
rect 34860 27570 34916 27580
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 33852 27134 33854 27186
rect 33906 27134 33908 27186
rect 33852 27122 33908 27134
rect 35868 26908 35924 28588
rect 36092 28644 36148 28654
rect 36092 28530 36148 28588
rect 36092 28478 36094 28530
rect 36146 28478 36148 28530
rect 36092 28466 36148 28478
rect 35756 26852 35924 26908
rect 35420 26628 35476 26638
rect 35476 26572 35588 26628
rect 35420 26562 35476 26572
rect 34412 26516 34468 26526
rect 33964 26460 34412 26516
rect 33964 26402 34020 26460
rect 34412 26422 34468 26460
rect 33964 26350 33966 26402
rect 34018 26350 34020 26402
rect 33964 26338 34020 26350
rect 33852 26066 33908 26078
rect 33852 26014 33854 26066
rect 33906 26014 33908 26066
rect 33852 25844 33908 26014
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 33852 25788 34356 25844
rect 35196 25834 35460 25844
rect 33852 25620 33908 25630
rect 34188 25620 34244 25630
rect 33852 25618 34188 25620
rect 33852 25566 33854 25618
rect 33906 25566 34188 25618
rect 33852 25564 34188 25566
rect 33852 25554 33908 25564
rect 34188 25526 34244 25564
rect 33740 25508 33796 25518
rect 33516 24994 33572 25004
rect 33628 25452 33740 25508
rect 33628 24722 33684 25452
rect 33740 25442 33796 25452
rect 33628 24670 33630 24722
rect 33682 24670 33684 24722
rect 33628 24658 33684 24670
rect 33740 25284 33796 25294
rect 33740 23938 33796 25228
rect 34076 25284 34132 25294
rect 34076 25190 34132 25228
rect 34188 24836 34244 24846
rect 34188 24722 34244 24780
rect 34188 24670 34190 24722
rect 34242 24670 34244 24722
rect 34188 24658 34244 24670
rect 33740 23886 33742 23938
rect 33794 23886 33796 23938
rect 33740 23874 33796 23886
rect 33516 23714 33572 23726
rect 33516 23662 33518 23714
rect 33570 23662 33572 23714
rect 33516 22820 33572 23662
rect 33628 23156 33684 23166
rect 33628 23062 33684 23100
rect 34076 23156 34132 23166
rect 34300 23156 34356 25788
rect 34972 25620 35028 25630
rect 34636 25508 34692 25518
rect 34636 25394 34692 25452
rect 34972 25506 35028 25564
rect 34972 25454 34974 25506
rect 35026 25454 35028 25506
rect 34972 25442 35028 25454
rect 34636 25342 34638 25394
rect 34690 25342 34692 25394
rect 34636 25330 34692 25342
rect 35308 25396 35364 25406
rect 35308 24612 35364 25340
rect 35420 25396 35476 25406
rect 35532 25396 35588 26572
rect 35420 25394 35588 25396
rect 35420 25342 35422 25394
rect 35474 25342 35588 25394
rect 35420 25340 35588 25342
rect 35756 25506 35812 26852
rect 36764 26178 36820 26190
rect 36764 26126 36766 26178
rect 36818 26126 36820 26178
rect 36204 25620 36260 25630
rect 36204 25526 36260 25564
rect 35756 25454 35758 25506
rect 35810 25454 35812 25506
rect 35420 25330 35476 25340
rect 35420 24724 35476 24734
rect 35420 24630 35476 24668
rect 35308 24546 35364 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35756 23938 35812 25454
rect 36764 25396 36820 26126
rect 36764 25330 36820 25340
rect 36092 25284 36148 25294
rect 36092 24834 36148 25228
rect 36092 24782 36094 24834
rect 36146 24782 36148 24834
rect 36092 24770 36148 24782
rect 36540 25172 36596 25182
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35756 23874 35812 23886
rect 35980 24612 36036 24622
rect 35980 23826 36036 24556
rect 35980 23774 35982 23826
rect 36034 23774 36036 23826
rect 35980 23762 36036 23774
rect 34132 23100 34356 23156
rect 34076 23062 34132 23100
rect 33516 22754 33572 22764
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22596 35588 22606
rect 33516 22484 33572 22494
rect 33516 22370 33572 22428
rect 33516 22318 33518 22370
rect 33570 22318 33572 22370
rect 33516 22306 33572 22318
rect 34300 22260 34356 22270
rect 34300 22258 34468 22260
rect 34300 22206 34302 22258
rect 34354 22206 34468 22258
rect 34300 22204 34468 22206
rect 34300 22194 34356 22204
rect 33180 17108 33236 17118
rect 33180 17014 33236 17052
rect 33068 16828 33236 16884
rect 33068 15874 33124 15886
rect 33068 15822 33070 15874
rect 33122 15822 33124 15874
rect 33068 15764 33124 15822
rect 33068 15698 33124 15708
rect 32620 14578 32676 14588
rect 32732 15092 33012 15148
rect 32732 13860 32788 15092
rect 32172 13010 32228 13020
rect 32284 13804 32788 13860
rect 32284 12292 32340 13804
rect 33068 13748 33124 13786
rect 33068 13682 33124 13692
rect 32396 13634 32452 13646
rect 32396 13582 32398 13634
rect 32450 13582 32452 13634
rect 32396 13074 32452 13582
rect 32396 13022 32398 13074
rect 32450 13022 32452 13074
rect 32396 12852 32452 13022
rect 32396 12786 32452 12796
rect 32508 13522 32564 13534
rect 33068 13524 33124 13534
rect 32508 13470 32510 13522
rect 32562 13470 32564 13522
rect 32508 12404 32564 13470
rect 32508 12338 32564 12348
rect 32732 13522 33124 13524
rect 32732 13470 33070 13522
rect 33122 13470 33124 13522
rect 32732 13468 33124 13470
rect 31612 11342 31614 11394
rect 31666 11342 31668 11394
rect 31612 11330 31668 11342
rect 31724 11676 31892 11732
rect 31948 12236 32340 12292
rect 31500 11118 31502 11170
rect 31554 11118 31556 11170
rect 31500 11106 31556 11118
rect 31164 10724 31220 10734
rect 31164 10630 31220 10668
rect 31724 10724 31780 11676
rect 31836 11508 31892 11518
rect 31836 11172 31892 11452
rect 31836 11106 31892 11116
rect 31724 10630 31780 10668
rect 31276 10612 31332 10622
rect 31276 10610 31556 10612
rect 31276 10558 31278 10610
rect 31330 10558 31556 10610
rect 31276 10556 31556 10558
rect 31276 10546 31332 10556
rect 31052 9986 31108 9996
rect 31164 9940 31220 9950
rect 31164 9826 31220 9884
rect 31164 9774 31166 9826
rect 31218 9774 31220 9826
rect 31164 9762 31220 9774
rect 31388 9828 31444 9838
rect 30716 9662 30718 9714
rect 30770 9662 30772 9714
rect 30716 9650 30772 9662
rect 30380 9602 30436 9614
rect 30380 9550 30382 9602
rect 30434 9550 30436 9602
rect 30380 8596 30436 9550
rect 30604 9604 30660 9614
rect 30604 9510 30660 9548
rect 31388 9266 31444 9772
rect 31388 9214 31390 9266
rect 31442 9214 31444 9266
rect 31388 9202 31444 9214
rect 31500 9714 31556 10556
rect 31836 9828 31892 9838
rect 31948 9828 32004 12236
rect 32732 12180 32788 13468
rect 33068 13458 33124 13468
rect 33180 13300 33236 16828
rect 33404 15148 33460 22092
rect 33628 21812 33684 21822
rect 33628 21718 33684 21756
rect 34412 21810 34468 22204
rect 34412 21758 34414 21810
rect 34466 21758 34468 21810
rect 34412 21746 34468 21758
rect 35532 21810 35588 22540
rect 36428 22596 36484 22606
rect 36428 22482 36484 22540
rect 36428 22430 36430 22482
rect 36482 22430 36484 22482
rect 36428 22418 36484 22430
rect 35532 21758 35534 21810
rect 35586 21758 35588 21810
rect 35532 21746 35588 21758
rect 36316 21812 36372 21822
rect 33964 21698 34020 21710
rect 33964 21646 33966 21698
rect 34018 21646 34020 21698
rect 33964 21588 34020 21646
rect 34524 21700 34580 21710
rect 34300 21588 34356 21598
rect 33964 21586 34356 21588
rect 33964 21534 34302 21586
rect 34354 21534 34356 21586
rect 33964 21532 34356 21534
rect 33516 20914 33572 20926
rect 33516 20862 33518 20914
rect 33570 20862 33572 20914
rect 33516 18452 33572 20862
rect 33964 20804 34020 20814
rect 33964 20710 34020 20748
rect 33740 20468 33796 20478
rect 33740 19236 33796 20412
rect 34300 19460 34356 21532
rect 34524 21586 34580 21644
rect 35756 21700 35812 21710
rect 36092 21700 36148 21710
rect 35756 21698 36260 21700
rect 35756 21646 35758 21698
rect 35810 21646 36094 21698
rect 36146 21646 36260 21698
rect 35756 21644 36260 21646
rect 35756 21634 35812 21644
rect 36092 21634 36148 21644
rect 34524 21534 34526 21586
rect 34578 21534 34580 21586
rect 34524 21522 34580 21534
rect 34860 21588 34916 21598
rect 34860 21494 34916 21532
rect 35084 21586 35140 21598
rect 35084 21534 35086 21586
rect 35138 21534 35140 21586
rect 34300 19394 34356 19404
rect 34188 19348 34244 19358
rect 34636 19348 34692 19358
rect 34188 19254 34244 19292
rect 34524 19292 34636 19348
rect 34076 19236 34132 19246
rect 33740 19234 34076 19236
rect 33740 19182 33742 19234
rect 33794 19182 34076 19234
rect 33740 19180 34076 19182
rect 33740 19170 33796 19180
rect 33852 18676 33908 18686
rect 33852 18582 33908 18620
rect 33516 18228 33572 18396
rect 33628 18564 33684 18574
rect 33628 18450 33684 18508
rect 33628 18398 33630 18450
rect 33682 18398 33684 18450
rect 33628 18386 33684 18398
rect 34076 18452 34132 19180
rect 34188 18452 34244 18462
rect 34076 18450 34244 18452
rect 34076 18398 34190 18450
rect 34242 18398 34244 18450
rect 34076 18396 34244 18398
rect 34188 18386 34244 18396
rect 33516 18172 33908 18228
rect 33628 16100 33684 16110
rect 33516 16044 33628 16100
rect 33852 16100 33908 18172
rect 34524 17444 34580 19292
rect 34636 19282 34692 19292
rect 34636 19010 34692 19022
rect 34636 18958 34638 19010
rect 34690 18958 34692 19010
rect 34636 18564 34692 18958
rect 34972 19012 35028 19022
rect 34972 18918 35028 18956
rect 35084 18676 35140 21534
rect 35644 21588 35700 21598
rect 35644 21494 35700 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35420 19236 35476 19246
rect 35420 19142 35476 19180
rect 35980 19012 36036 19022
rect 35980 19010 36148 19012
rect 35980 18958 35982 19010
rect 36034 18958 36148 19010
rect 35980 18956 36148 18958
rect 35980 18946 36036 18956
rect 35084 18610 35140 18620
rect 34636 18498 34692 18508
rect 35980 18564 36036 18574
rect 34748 18450 34804 18462
rect 34748 18398 34750 18450
rect 34802 18398 34804 18450
rect 34748 17668 34804 18398
rect 35308 18450 35364 18462
rect 35308 18398 35310 18450
rect 35362 18398 35364 18450
rect 35308 18340 35364 18398
rect 35308 18274 35364 18284
rect 35532 18452 35588 18462
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17778 35588 18396
rect 35980 18450 36036 18508
rect 35980 18398 35982 18450
rect 36034 18398 36036 18450
rect 35980 18386 36036 18398
rect 35532 17726 35534 17778
rect 35586 17726 35588 17778
rect 35084 17668 35140 17678
rect 34748 17666 35140 17668
rect 34748 17614 35086 17666
rect 35138 17614 35140 17666
rect 34748 17612 35140 17614
rect 35084 17444 35140 17612
rect 34524 17388 34916 17444
rect 33964 16100 34020 16110
rect 33852 16098 34020 16100
rect 33852 16046 33966 16098
rect 34018 16046 34020 16098
rect 33852 16044 34020 16046
rect 33516 15538 33572 16044
rect 33628 16006 33684 16044
rect 33964 16034 34020 16044
rect 34300 15988 34356 15998
rect 34300 15894 34356 15932
rect 33516 15486 33518 15538
rect 33570 15486 33572 15538
rect 33516 15474 33572 15486
rect 33852 15876 33908 15886
rect 33740 15204 33796 15214
rect 33404 15092 33572 15148
rect 32284 12124 32788 12180
rect 32844 13244 33236 13300
rect 33404 13522 33460 13534
rect 33404 13470 33406 13522
rect 33458 13470 33460 13522
rect 32060 11620 32116 11630
rect 32060 11526 32116 11564
rect 32284 11394 32340 12124
rect 32844 12068 32900 13244
rect 33068 13076 33124 13086
rect 33068 12402 33124 13020
rect 33404 13076 33460 13470
rect 33404 13010 33460 13020
rect 33068 12350 33070 12402
rect 33122 12350 33124 12402
rect 33068 12338 33124 12350
rect 33292 12962 33348 12974
rect 33292 12910 33294 12962
rect 33346 12910 33348 12962
rect 33292 12852 33348 12910
rect 33292 12178 33348 12796
rect 33292 12126 33294 12178
rect 33346 12126 33348 12178
rect 32284 11342 32286 11394
rect 32338 11342 32340 11394
rect 32284 11330 32340 11342
rect 32508 12012 32900 12068
rect 33180 12066 33236 12078
rect 33180 12014 33182 12066
rect 33234 12014 33236 12066
rect 32284 9940 32340 9950
rect 32284 9846 32340 9884
rect 31892 9772 32004 9828
rect 31836 9734 31892 9772
rect 31500 9662 31502 9714
rect 31554 9662 31556 9714
rect 31052 9154 31108 9166
rect 31052 9102 31054 9154
rect 31106 9102 31108 9154
rect 31052 8596 31108 9102
rect 30380 8540 31108 8596
rect 30604 8146 30660 8540
rect 30604 8094 30606 8146
rect 30658 8094 30660 8146
rect 30268 7756 30548 7812
rect 29820 7534 29822 7586
rect 29874 7534 29876 7586
rect 29820 7522 29876 7534
rect 27580 6690 28084 6692
rect 27580 6638 27582 6690
rect 27634 6638 28030 6690
rect 28082 6638 28084 6690
rect 27580 6636 28084 6638
rect 27580 6626 27636 6636
rect 28028 6626 28084 6636
rect 28140 7476 28196 7486
rect 27244 6526 27246 6578
rect 27298 6526 27300 6578
rect 27244 6514 27300 6526
rect 26012 6290 26068 6300
rect 28140 6244 28196 7420
rect 30492 7474 30548 7756
rect 30492 7422 30494 7474
rect 30546 7422 30548 7474
rect 30156 6692 30212 6702
rect 30268 6692 30324 6702
rect 30156 6690 30324 6692
rect 30156 6638 30158 6690
rect 30210 6638 30270 6690
rect 30322 6638 30324 6690
rect 30156 6636 30324 6638
rect 30156 6626 30212 6636
rect 30268 6580 30324 6636
rect 30268 6514 30324 6524
rect 30492 6692 30548 7422
rect 27580 6132 27636 6142
rect 27580 5794 27636 6076
rect 27580 5742 27582 5794
rect 27634 5742 27636 5794
rect 27580 5730 27636 5742
rect 25900 5182 25902 5234
rect 25954 5182 25956 5234
rect 25900 5170 25956 5182
rect 26012 4898 26068 4910
rect 26012 4846 26014 4898
rect 26066 4846 26068 4898
rect 26012 4450 26068 4846
rect 26012 4398 26014 4450
rect 26066 4398 26068 4450
rect 26012 4386 26068 4398
rect 25340 4340 25396 4350
rect 25340 4246 25396 4284
rect 24444 4174 24446 4226
rect 24498 4174 24500 4226
rect 24444 4162 24500 4174
rect 28140 4226 28196 6188
rect 30492 5906 30548 6636
rect 30492 5854 30494 5906
rect 30546 5854 30548 5906
rect 29708 5794 29764 5806
rect 29708 5742 29710 5794
rect 29762 5742 29764 5794
rect 29372 5460 29428 5470
rect 28588 4564 28644 4574
rect 28588 4470 28644 4508
rect 28140 4174 28142 4226
rect 28194 4174 28196 4226
rect 28140 4162 28196 4174
rect 29372 4226 29428 5404
rect 29708 5236 29764 5742
rect 29708 5170 29764 5180
rect 30492 4564 30548 5854
rect 30604 5796 30660 8094
rect 30940 8372 30996 8382
rect 30940 8258 30996 8316
rect 30940 8206 30942 8258
rect 30994 8206 30996 8258
rect 30716 8036 30772 8046
rect 30716 7942 30772 7980
rect 30940 7700 30996 8206
rect 31500 8258 31556 9662
rect 32508 8596 32564 12012
rect 33180 11956 33236 12014
rect 32620 11900 33236 11956
rect 32620 11394 32676 11900
rect 33068 11618 33124 11630
rect 33068 11566 33070 11618
rect 33122 11566 33124 11618
rect 33068 11506 33124 11566
rect 33068 11454 33070 11506
rect 33122 11454 33124 11506
rect 33068 11442 33124 11454
rect 32620 11342 32622 11394
rect 32674 11342 32676 11394
rect 32620 11330 32676 11342
rect 33292 11284 33348 12126
rect 33404 12740 33460 12750
rect 33404 12180 33460 12684
rect 33404 11618 33460 12124
rect 33404 11566 33406 11618
rect 33458 11566 33460 11618
rect 33404 11554 33460 11566
rect 33516 11396 33572 15092
rect 33740 14532 33796 15148
rect 33852 15148 33908 15820
rect 33964 15874 34020 15886
rect 33964 15822 33966 15874
rect 34018 15822 34020 15874
rect 33964 15540 34020 15822
rect 33964 15484 34692 15540
rect 33852 15092 34356 15148
rect 33740 14476 33908 14532
rect 33740 14306 33796 14318
rect 33740 14254 33742 14306
rect 33794 14254 33796 14306
rect 33740 13748 33796 14254
rect 33740 13682 33796 13692
rect 33852 13746 33908 14476
rect 34076 14196 34132 14206
rect 33852 13694 33854 13746
rect 33906 13694 33908 13746
rect 33628 12962 33684 12974
rect 33628 12910 33630 12962
rect 33682 12910 33684 12962
rect 33628 12180 33684 12910
rect 33852 12292 33908 13694
rect 33964 14140 34076 14196
rect 33964 13300 34020 14140
rect 34076 14130 34132 14140
rect 34300 13858 34356 15092
rect 34636 14642 34692 15484
rect 34636 14590 34638 14642
rect 34690 14590 34692 14642
rect 34636 14578 34692 14590
rect 34860 14196 34916 17388
rect 35084 17378 35140 17388
rect 35532 16996 35588 17726
rect 35532 16930 35588 16940
rect 35980 17444 36036 17454
rect 36092 17444 36148 18956
rect 36204 18788 36260 21644
rect 36316 21586 36372 21756
rect 36316 21534 36318 21586
rect 36370 21534 36372 21586
rect 36316 21522 36372 21534
rect 36316 18788 36372 18798
rect 36204 18732 36316 18788
rect 36316 18722 36372 18732
rect 36036 17388 36148 17444
rect 35980 16996 36036 17388
rect 36540 17332 36596 25116
rect 36764 21812 36820 21822
rect 36764 21718 36820 21756
rect 36876 18452 36932 29036
rect 37324 28644 37380 28654
rect 37324 28550 37380 28588
rect 37324 28420 37380 28430
rect 37212 28364 37324 28420
rect 37100 27300 37156 27310
rect 36988 26964 37044 26974
rect 36988 25506 37044 26908
rect 37100 26516 37156 27244
rect 37100 26450 37156 26460
rect 36988 25454 36990 25506
rect 37042 25454 37044 25506
rect 36988 25442 37044 25454
rect 37100 25284 37156 25294
rect 37100 25190 37156 25228
rect 37212 22258 37268 28364
rect 37324 28354 37380 28364
rect 37436 28196 37492 29374
rect 37772 28530 37828 29820
rect 37884 29428 37940 29438
rect 37884 28754 37940 29372
rect 37884 28702 37886 28754
rect 37938 28702 37940 28754
rect 37884 28690 37940 28702
rect 37772 28478 37774 28530
rect 37826 28478 37828 28530
rect 37772 28466 37828 28478
rect 37996 28530 38052 28542
rect 37996 28478 37998 28530
rect 38050 28478 38052 28530
rect 37436 28130 37492 28140
rect 37772 27746 37828 27758
rect 37772 27694 37774 27746
rect 37826 27694 37828 27746
rect 37772 27636 37828 27694
rect 37772 27570 37828 27580
rect 37996 27074 38052 28478
rect 38108 28420 38164 32060
rect 38220 31892 38276 31902
rect 38220 31778 38276 31836
rect 38220 31726 38222 31778
rect 38274 31726 38276 31778
rect 38220 31714 38276 31726
rect 38108 28354 38164 28364
rect 37996 27022 37998 27074
rect 38050 27022 38052 27074
rect 37660 26628 37716 26638
rect 37660 26516 37716 26572
rect 37436 26514 37716 26516
rect 37436 26462 37662 26514
rect 37714 26462 37716 26514
rect 37436 26460 37716 26462
rect 37324 25732 37380 25742
rect 37324 25396 37380 25676
rect 37324 25302 37380 25340
rect 37436 25284 37492 26460
rect 37660 26450 37716 26460
rect 37996 26516 38052 27022
rect 38108 28196 38164 28206
rect 38108 27970 38164 28140
rect 38108 27918 38110 27970
rect 38162 27918 38164 27970
rect 38108 27748 38164 27918
rect 38108 26964 38164 27692
rect 38220 27970 38276 27982
rect 38220 27918 38222 27970
rect 38274 27918 38276 27970
rect 38220 27300 38276 27918
rect 38220 27234 38276 27244
rect 38220 26964 38276 26974
rect 38164 26962 38276 26964
rect 38164 26910 38222 26962
rect 38274 26910 38276 26962
rect 38164 26908 38276 26910
rect 38108 26898 38164 26908
rect 38220 26898 38276 26908
rect 37996 26450 38052 26460
rect 38332 25732 38388 33292
rect 38444 33282 38500 33292
rect 38668 32788 38724 33516
rect 38892 33348 38948 33358
rect 38892 33254 38948 33292
rect 39116 33234 39172 34748
rect 39340 34692 39396 34702
rect 39228 34132 39284 34142
rect 39340 34132 39396 34636
rect 39284 34076 39396 34132
rect 39676 34132 39732 34142
rect 39228 34038 39284 34076
rect 39676 34038 39732 34076
rect 39788 33572 39844 39452
rect 40012 38834 40068 38846
rect 40012 38782 40014 38834
rect 40066 38782 40068 38834
rect 39900 37492 39956 37502
rect 40012 37492 40068 38782
rect 40236 38612 40292 40126
rect 41692 39618 41748 40348
rect 41692 39566 41694 39618
rect 41746 39566 41748 39618
rect 41692 39508 41748 39566
rect 41692 39442 41748 39452
rect 40236 38050 40292 38556
rect 40236 37998 40238 38050
rect 40290 37998 40292 38050
rect 40236 37986 40292 37998
rect 41580 38050 41636 38062
rect 41580 37998 41582 38050
rect 41634 37998 41636 38050
rect 39900 37490 40068 37492
rect 39900 37438 39902 37490
rect 39954 37438 40068 37490
rect 39900 37436 40068 37438
rect 40796 37826 40852 37838
rect 40796 37774 40798 37826
rect 40850 37774 40852 37826
rect 39900 37426 39956 37436
rect 40796 36708 40852 37774
rect 40908 37156 40964 37166
rect 40908 37062 40964 37100
rect 41244 37156 41300 37166
rect 40908 36708 40964 36718
rect 40796 36706 40964 36708
rect 40796 36654 40910 36706
rect 40962 36654 40964 36706
rect 40796 36652 40964 36654
rect 40908 36642 40964 36652
rect 41244 36706 41300 37100
rect 41244 36654 41246 36706
rect 41298 36654 41300 36706
rect 41244 36642 41300 36654
rect 41132 36260 41188 36270
rect 41580 36260 41636 37998
rect 41804 37268 41860 41692
rect 41804 37202 41860 37212
rect 41692 36260 41748 36270
rect 41132 36258 41748 36260
rect 41132 36206 41134 36258
rect 41186 36206 41694 36258
rect 41746 36206 41748 36258
rect 41132 36204 41748 36206
rect 40124 35252 40180 35262
rect 40124 34244 40180 35196
rect 40796 35028 40852 35038
rect 40796 34934 40852 34972
rect 40124 34130 40180 34188
rect 40124 34078 40126 34130
rect 40178 34078 40180 34130
rect 40124 34066 40180 34078
rect 40236 34468 40292 34478
rect 39116 33182 39118 33234
rect 39170 33182 39172 33234
rect 39116 33170 39172 33182
rect 39452 33516 39844 33572
rect 39004 32788 39060 32798
rect 38668 32786 39060 32788
rect 38668 32734 39006 32786
rect 39058 32734 39060 32786
rect 38668 32732 39060 32734
rect 39004 32722 39060 32732
rect 38444 32562 38500 32574
rect 38444 32510 38446 32562
rect 38498 32510 38500 32562
rect 38444 31780 38500 32510
rect 38780 31780 38836 31790
rect 38444 31714 38500 31724
rect 38668 31778 38836 31780
rect 38668 31726 38782 31778
rect 38834 31726 38836 31778
rect 38668 31724 38836 31726
rect 38668 29988 38724 31724
rect 38780 31714 38836 31724
rect 39452 31668 39508 33516
rect 39788 33346 39844 33358
rect 39788 33294 39790 33346
rect 39842 33294 39844 33346
rect 39564 32340 39620 32350
rect 39564 31890 39620 32284
rect 39564 31838 39566 31890
rect 39618 31838 39620 31890
rect 39564 31826 39620 31838
rect 39452 31612 39620 31668
rect 38668 28642 38724 29932
rect 39116 29204 39172 29214
rect 38668 28590 38670 28642
rect 38722 28590 38724 28642
rect 38668 28578 38724 28590
rect 38892 29148 39116 29204
rect 38780 28084 38836 28094
rect 38444 27972 38500 27982
rect 38444 27878 38500 27916
rect 38668 27858 38724 27870
rect 38668 27806 38670 27858
rect 38722 27806 38724 27858
rect 38668 27748 38724 27806
rect 38668 27682 38724 27692
rect 38668 27300 38724 27310
rect 38668 27186 38724 27244
rect 38668 27134 38670 27186
rect 38722 27134 38724 27186
rect 38668 27122 38724 27134
rect 38780 27188 38836 28028
rect 38892 28082 38948 29148
rect 39116 29138 39172 29148
rect 39340 28532 39396 28542
rect 39340 28530 39508 28532
rect 39340 28478 39342 28530
rect 39394 28478 39508 28530
rect 39340 28476 39508 28478
rect 39340 28466 39396 28476
rect 38892 28030 38894 28082
rect 38946 28030 38948 28082
rect 38892 28018 38948 28030
rect 39004 27972 39060 27982
rect 39004 27878 39060 27916
rect 39116 27970 39172 27982
rect 39116 27918 39118 27970
rect 39170 27918 39172 27970
rect 39116 27636 39172 27918
rect 39452 27746 39508 28476
rect 39452 27694 39454 27746
rect 39506 27694 39508 27746
rect 39452 27682 39508 27694
rect 39116 27570 39172 27580
rect 38892 27188 38948 27198
rect 38780 27132 38892 27188
rect 38220 25676 38388 25732
rect 38444 26516 38500 26526
rect 37548 25396 37604 25406
rect 37548 25302 37604 25340
rect 37436 25218 37492 25228
rect 37996 25284 38052 25294
rect 37996 25190 38052 25228
rect 38220 25282 38276 25676
rect 38444 25506 38500 26460
rect 38444 25454 38446 25506
rect 38498 25454 38500 25506
rect 38444 25442 38500 25454
rect 38332 25396 38388 25406
rect 38332 25302 38388 25340
rect 38220 25230 38222 25282
rect 38274 25230 38276 25282
rect 38220 24610 38276 25230
rect 38220 24558 38222 24610
rect 38274 24558 38276 24610
rect 38220 24546 38276 24558
rect 38444 24724 38500 24734
rect 38892 24724 38948 27132
rect 39228 26516 39284 26526
rect 39452 26516 39508 26526
rect 39228 26422 39284 26460
rect 39340 26460 39452 26516
rect 39116 26068 39172 26078
rect 39116 25974 39172 26012
rect 39004 25620 39060 25630
rect 39340 25620 39396 26460
rect 39452 26450 39508 26460
rect 39452 26292 39508 26302
rect 39452 26198 39508 26236
rect 39004 25618 39396 25620
rect 39004 25566 39006 25618
rect 39058 25566 39342 25618
rect 39394 25566 39396 25618
rect 39004 25564 39396 25566
rect 39004 25554 39060 25564
rect 39340 25554 39396 25564
rect 39228 25396 39284 25406
rect 39228 24946 39284 25340
rect 39564 25172 39620 31612
rect 39788 30324 39844 33294
rect 40236 33346 40292 34412
rect 41132 34356 41188 36204
rect 41692 36194 41748 36204
rect 40796 34300 41188 34356
rect 41244 35028 41300 35038
rect 41244 34354 41300 34972
rect 41244 34302 41246 34354
rect 41298 34302 41300 34354
rect 40236 33294 40238 33346
rect 40290 33294 40292 33346
rect 40236 33282 40292 33294
rect 40460 34132 40516 34142
rect 40460 32676 40516 34076
rect 40460 32582 40516 32620
rect 39900 30324 39956 30334
rect 39788 30322 39956 30324
rect 39788 30270 39902 30322
rect 39954 30270 39956 30322
rect 39788 30268 39956 30270
rect 39788 29876 39844 30268
rect 39900 30258 39956 30268
rect 40348 29988 40404 29998
rect 40348 29894 40404 29932
rect 39788 29810 39844 29820
rect 40236 29316 40292 29326
rect 40236 29222 40292 29260
rect 40124 29204 40180 29214
rect 40124 29110 40180 29148
rect 40012 27188 40068 27198
rect 40012 27094 40068 27132
rect 40796 26908 40852 34300
rect 41244 34290 41300 34302
rect 41468 34356 41524 34366
rect 41468 34262 41524 34300
rect 41244 34132 41300 34142
rect 41244 33348 41300 34076
rect 41692 34132 41748 34142
rect 41692 34130 41860 34132
rect 41692 34078 41694 34130
rect 41746 34078 41860 34130
rect 41692 34076 41860 34078
rect 41692 34066 41748 34076
rect 41580 34018 41636 34030
rect 41580 33966 41582 34018
rect 41634 33966 41636 34018
rect 41580 33348 41636 33966
rect 41692 33348 41748 33358
rect 41244 33346 41524 33348
rect 41244 33294 41246 33346
rect 41298 33294 41524 33346
rect 41244 33292 41524 33294
rect 41580 33346 41748 33348
rect 41580 33294 41694 33346
rect 41746 33294 41748 33346
rect 41580 33292 41748 33294
rect 41244 33282 41300 33292
rect 41468 33124 41524 33292
rect 41692 33282 41748 33292
rect 41804 33236 41860 34076
rect 41804 33170 41860 33180
rect 41468 33068 41748 33124
rect 40908 32564 40964 32574
rect 40908 32470 40964 32508
rect 41468 32562 41524 32574
rect 41468 32510 41470 32562
rect 41522 32510 41524 32562
rect 41468 31892 41524 32510
rect 41468 31826 41524 31836
rect 41692 31890 41748 33068
rect 41804 32676 41860 32686
rect 41804 32582 41860 32620
rect 41916 32564 41972 45276
rect 42140 44324 42196 45950
rect 42140 43708 42196 44268
rect 42140 43652 42532 43708
rect 42252 43428 42308 43438
rect 42252 42980 42308 43372
rect 42476 43428 42532 43652
rect 42476 43334 42532 43372
rect 42028 42644 42084 42654
rect 42028 42550 42084 42588
rect 42252 42642 42308 42924
rect 42252 42590 42254 42642
rect 42306 42590 42308 42642
rect 42252 42578 42308 42590
rect 42140 41858 42196 41870
rect 42140 41806 42142 41858
rect 42194 41806 42196 41858
rect 42140 40404 42196 41806
rect 42252 41076 42308 41086
rect 42252 40982 42308 41020
rect 42588 41076 42644 41086
rect 42140 40338 42196 40348
rect 42252 39394 42308 39406
rect 42252 39342 42254 39394
rect 42306 39342 42308 39394
rect 42252 39284 42308 39342
rect 42140 39228 42252 39284
rect 42140 38050 42196 39228
rect 42252 39218 42308 39228
rect 42140 37998 42142 38050
rect 42194 37998 42196 38050
rect 42140 37986 42196 37998
rect 42476 35700 42532 35710
rect 42364 34916 42420 34926
rect 42364 34356 42420 34860
rect 42140 34300 42364 34356
rect 42028 34132 42084 34142
rect 42028 34038 42084 34076
rect 42028 33348 42084 33358
rect 42140 33348 42196 34300
rect 42364 34262 42420 34300
rect 42028 33346 42196 33348
rect 42028 33294 42030 33346
rect 42082 33294 42196 33346
rect 42028 33292 42196 33294
rect 42364 33346 42420 33358
rect 42364 33294 42366 33346
rect 42418 33294 42420 33346
rect 42028 33282 42084 33292
rect 42364 33236 42420 33294
rect 42364 33170 42420 33180
rect 41916 32498 41972 32508
rect 42028 33122 42084 33134
rect 42028 33070 42030 33122
rect 42082 33070 42084 33122
rect 42028 32340 42084 33070
rect 42028 32274 42084 32284
rect 42252 32564 42308 32574
rect 42252 32450 42308 32508
rect 42252 32398 42254 32450
rect 42306 32398 42308 32450
rect 42252 32340 42308 32398
rect 42252 32274 42308 32284
rect 41692 31838 41694 31890
rect 41746 31838 41748 31890
rect 41692 31826 41748 31838
rect 42140 31892 42196 31902
rect 42476 31892 42532 35644
rect 42588 35252 42644 41020
rect 42700 36932 42756 47852
rect 42924 47572 42980 50372
rect 43148 48916 43204 48926
rect 43260 48916 43316 51324
rect 43372 49700 43428 51886
rect 43708 51604 43764 51614
rect 43708 51378 43764 51548
rect 43708 51326 43710 51378
rect 43762 51326 43764 51378
rect 43708 51314 43764 51326
rect 44156 50596 44212 51996
rect 44380 51268 44436 51278
rect 45276 51268 45332 51278
rect 44380 51266 44996 51268
rect 44380 51214 44382 51266
rect 44434 51214 44996 51266
rect 44380 51212 44996 51214
rect 44380 51202 44436 51212
rect 44940 50706 44996 51212
rect 44940 50654 44942 50706
rect 44994 50654 44996 50706
rect 44940 50642 44996 50654
rect 44156 50530 44212 50540
rect 44828 50596 44884 50606
rect 44828 50502 44884 50540
rect 45052 50372 45108 50382
rect 43372 49634 43428 49644
rect 44940 50370 45108 50372
rect 44940 50318 45054 50370
rect 45106 50318 45108 50370
rect 44940 50316 45108 50318
rect 43148 48914 43316 48916
rect 43148 48862 43150 48914
rect 43202 48862 43316 48914
rect 43148 48860 43316 48862
rect 43148 48850 43204 48860
rect 43036 48802 43092 48814
rect 43036 48750 43038 48802
rect 43090 48750 43092 48802
rect 43036 48244 43092 48750
rect 43036 48178 43092 48188
rect 43260 48242 43316 48860
rect 43372 48356 43428 48366
rect 43372 48262 43428 48300
rect 43260 48190 43262 48242
rect 43314 48190 43316 48242
rect 42924 47506 42980 47516
rect 43260 46788 43316 48190
rect 43484 48244 43540 48254
rect 43484 47236 43540 48188
rect 43932 48242 43988 48254
rect 43932 48190 43934 48242
rect 43986 48190 43988 48242
rect 43484 47170 43540 47180
rect 43596 47572 43652 47582
rect 43260 46722 43316 46732
rect 43596 45108 43652 47516
rect 43932 47012 43988 48190
rect 44268 47572 44324 47582
rect 44268 47478 44324 47516
rect 44828 47572 44884 47582
rect 44828 47458 44884 47516
rect 44828 47406 44830 47458
rect 44882 47406 44884 47458
rect 44828 47394 44884 47406
rect 43932 46946 43988 46956
rect 44828 47236 44884 47246
rect 44492 46676 44548 46686
rect 44492 46582 44548 46620
rect 44828 46674 44884 47180
rect 44828 46622 44830 46674
rect 44882 46622 44884 46674
rect 44828 46610 44884 46622
rect 43820 45108 43876 45118
rect 43596 45106 43876 45108
rect 43596 45054 43822 45106
rect 43874 45054 43876 45106
rect 43596 45052 43876 45054
rect 43820 45042 43876 45052
rect 44940 44884 44996 50316
rect 45052 50306 45108 50316
rect 45276 48244 45332 51212
rect 45500 50594 45556 52220
rect 45500 50542 45502 50594
rect 45554 50542 45556 50594
rect 45500 50530 45556 50542
rect 45836 50596 45892 50606
rect 45836 50502 45892 50540
rect 46060 50596 46116 54462
rect 46396 54516 46452 54526
rect 46396 54422 46452 54460
rect 46620 54514 46676 54526
rect 46620 54462 46622 54514
rect 46674 54462 46676 54514
rect 46620 53172 46676 54462
rect 46956 54516 47012 55132
rect 46956 54450 47012 54460
rect 46844 54404 46900 54414
rect 46844 54310 46900 54348
rect 47180 54404 47236 54414
rect 47740 54404 47796 55356
rect 47180 54402 47796 54404
rect 47180 54350 47182 54402
rect 47234 54350 47796 54402
rect 47180 54348 47796 54350
rect 47852 54404 47908 55918
rect 47180 54338 47236 54348
rect 47852 53844 47908 54348
rect 47516 53284 47572 53294
rect 46172 53170 46676 53172
rect 46172 53118 46622 53170
rect 46674 53118 46676 53170
rect 46172 53116 46676 53118
rect 46172 52722 46228 53116
rect 46620 53106 46676 53116
rect 46844 53172 46900 53182
rect 46900 53116 47012 53172
rect 46844 53078 46900 53116
rect 46396 52948 46452 52958
rect 46396 52854 46452 52892
rect 46732 52948 46788 52958
rect 46508 52836 46564 52846
rect 46732 52836 46788 52892
rect 46508 52742 46564 52780
rect 46620 52780 46788 52836
rect 46172 52670 46174 52722
rect 46226 52670 46228 52722
rect 46172 52658 46228 52670
rect 46620 52162 46676 52780
rect 46732 52276 46788 52314
rect 46732 52210 46788 52220
rect 46620 52110 46622 52162
rect 46674 52110 46676 52162
rect 46620 52098 46676 52110
rect 46956 52164 47012 53116
rect 47516 53170 47572 53228
rect 47516 53118 47518 53170
rect 47570 53118 47572 53170
rect 47068 52948 47124 52958
rect 47516 52948 47572 53118
rect 47068 52946 47348 52948
rect 47068 52894 47070 52946
rect 47122 52894 47348 52946
rect 47068 52892 47348 52894
rect 47068 52882 47124 52892
rect 47180 52724 47236 52734
rect 46956 52108 47124 52164
rect 47068 52050 47124 52108
rect 47068 51998 47070 52050
rect 47122 51998 47124 52050
rect 47068 51986 47124 51998
rect 46844 51938 46900 51950
rect 46844 51886 46846 51938
rect 46898 51886 46900 51938
rect 46844 51380 46900 51886
rect 47180 51602 47236 52668
rect 47292 52722 47348 52892
rect 47292 52670 47294 52722
rect 47346 52670 47348 52722
rect 47292 52658 47348 52670
rect 47292 52052 47348 52062
rect 47292 52050 47460 52052
rect 47292 51998 47294 52050
rect 47346 51998 47460 52050
rect 47292 51996 47460 51998
rect 47292 51986 47348 51996
rect 47180 51550 47182 51602
rect 47234 51550 47236 51602
rect 47180 51538 47236 51550
rect 46956 51380 47012 51390
rect 46508 51378 47012 51380
rect 46508 51326 46958 51378
rect 47010 51326 47012 51378
rect 46508 51324 47012 51326
rect 46508 51266 46564 51324
rect 46956 51314 47012 51324
rect 47292 51380 47348 51390
rect 47292 51286 47348 51324
rect 46508 51214 46510 51266
rect 46562 51214 46564 51266
rect 46508 51202 46564 51214
rect 47404 50932 47460 51996
rect 47180 50876 47460 50932
rect 46060 50530 46116 50540
rect 46732 50596 46788 50606
rect 47180 50596 47236 50876
rect 46732 50502 46788 50540
rect 46844 50594 47236 50596
rect 46844 50542 47182 50594
rect 47234 50542 47236 50594
rect 46844 50540 47236 50542
rect 46732 49140 46788 49150
rect 46844 49140 46900 50540
rect 47180 50530 47236 50540
rect 47404 50596 47460 50606
rect 47516 50596 47572 52892
rect 47628 52722 47684 52734
rect 47628 52670 47630 52722
rect 47682 52670 47684 52722
rect 47628 52276 47684 52670
rect 47628 52274 47796 52276
rect 47628 52222 47630 52274
rect 47682 52222 47796 52274
rect 47628 52220 47796 52222
rect 47628 52210 47684 52220
rect 47404 50594 47572 50596
rect 47404 50542 47406 50594
rect 47458 50542 47572 50594
rect 47404 50540 47572 50542
rect 47404 50530 47460 50540
rect 47516 50428 47572 50540
rect 47628 51378 47684 51390
rect 47628 51326 47630 51378
rect 47682 51326 47684 51378
rect 47628 50596 47684 51326
rect 47740 51044 47796 52220
rect 47852 51266 47908 53788
rect 47964 53284 48020 56252
rect 48076 56082 48132 57372
rect 48188 57362 48244 57372
rect 49196 56756 49252 56766
rect 48860 56754 49252 56756
rect 48860 56702 49198 56754
rect 49250 56702 49252 56754
rect 48860 56700 49252 56702
rect 48188 56308 48244 56318
rect 48188 56306 48804 56308
rect 48188 56254 48190 56306
rect 48242 56254 48804 56306
rect 48188 56252 48804 56254
rect 48188 56242 48244 56252
rect 48748 56194 48804 56252
rect 48860 56306 48916 56700
rect 49196 56690 49252 56700
rect 48860 56254 48862 56306
rect 48914 56254 48916 56306
rect 48860 56242 48916 56254
rect 48748 56142 48750 56194
rect 48802 56142 48804 56194
rect 48748 56130 48804 56142
rect 48076 56030 48078 56082
rect 48130 56030 48132 56082
rect 48076 56018 48132 56030
rect 49308 55188 49364 59166
rect 49420 59218 49476 59230
rect 49420 59166 49422 59218
rect 49474 59166 49476 59218
rect 49420 57428 49476 59166
rect 49644 59106 49700 59948
rect 49868 59220 49924 60062
rect 50204 59890 50260 60844
rect 50988 60676 51044 60686
rect 50988 60002 51044 60620
rect 50988 59950 50990 60002
rect 51042 59950 51044 60002
rect 50988 59938 51044 59950
rect 51100 60004 51156 63086
rect 51212 63138 51268 63982
rect 51324 63924 51380 63934
rect 51324 63830 51380 63868
rect 51212 63086 51214 63138
rect 51266 63086 51268 63138
rect 51212 63074 51268 63086
rect 51436 63250 51492 63262
rect 51436 63198 51438 63250
rect 51490 63198 51492 63250
rect 51436 61012 51492 63198
rect 51660 63250 51716 64542
rect 51660 63198 51662 63250
rect 51714 63198 51716 63250
rect 51660 63186 51716 63198
rect 51772 63140 51828 63150
rect 51996 63140 52052 65326
rect 51772 63138 52052 63140
rect 51772 63086 51774 63138
rect 51826 63086 52052 63138
rect 51772 63084 52052 63086
rect 52108 64484 52164 64494
rect 51660 62244 51716 62254
rect 51660 62150 51716 62188
rect 51436 60946 51492 60956
rect 51212 60786 51268 60798
rect 51660 60788 51716 60798
rect 51212 60734 51214 60786
rect 51266 60734 51268 60786
rect 51212 60228 51268 60734
rect 51212 60162 51268 60172
rect 51548 60732 51660 60788
rect 51212 60004 51268 60014
rect 51100 60002 51268 60004
rect 51100 59950 51214 60002
rect 51266 59950 51268 60002
rect 51100 59948 51268 59950
rect 50204 59838 50206 59890
rect 50258 59838 50260 59890
rect 50204 59826 50260 59838
rect 50540 59780 50596 59790
rect 50540 59778 50932 59780
rect 50540 59726 50542 59778
rect 50594 59726 50932 59778
rect 50540 59724 50932 59726
rect 50540 59714 50596 59724
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50876 59556 50932 59724
rect 51100 59778 51156 59790
rect 51100 59726 51102 59778
rect 51154 59726 51156 59778
rect 51100 59556 51156 59726
rect 50876 59500 51156 59556
rect 50428 59444 50484 59454
rect 49980 59220 50036 59230
rect 49868 59218 50036 59220
rect 49868 59166 49982 59218
rect 50034 59166 50036 59218
rect 49868 59164 50036 59166
rect 49980 59154 50036 59164
rect 49644 59054 49646 59106
rect 49698 59054 49700 59106
rect 49644 59042 49700 59054
rect 49420 57362 49476 57372
rect 49868 58884 49924 58894
rect 49308 55122 49364 55132
rect 49196 55074 49252 55086
rect 49196 55022 49198 55074
rect 49250 55022 49252 55074
rect 49196 54628 49252 55022
rect 49532 55076 49588 55086
rect 49532 54982 49588 55020
rect 49196 54562 49252 54572
rect 47964 53170 48020 53228
rect 47964 53118 47966 53170
rect 48018 53118 48020 53170
rect 47964 53106 48020 53118
rect 49756 52052 49812 52062
rect 48860 52050 49812 52052
rect 48860 51998 49758 52050
rect 49810 51998 49812 52050
rect 48860 51996 49812 51998
rect 48300 51604 48356 51614
rect 48300 51602 48804 51604
rect 48300 51550 48302 51602
rect 48354 51550 48804 51602
rect 48300 51548 48804 51550
rect 48300 51538 48356 51548
rect 48748 51490 48804 51548
rect 48860 51602 48916 51996
rect 49756 51986 49812 51996
rect 48860 51550 48862 51602
rect 48914 51550 48916 51602
rect 48860 51538 48916 51550
rect 48748 51438 48750 51490
rect 48802 51438 48804 51490
rect 48748 51426 48804 51438
rect 47852 51214 47854 51266
rect 47906 51214 47908 51266
rect 47852 51202 47908 51214
rect 48188 51266 48244 51278
rect 48188 51214 48190 51266
rect 48242 51214 48244 51266
rect 48188 51044 48244 51214
rect 47740 50988 48244 51044
rect 47628 50530 47684 50540
rect 47852 50482 47908 50494
rect 47852 50430 47854 50482
rect 47906 50430 47908 50482
rect 47852 50428 47908 50430
rect 46732 49138 46900 49140
rect 46732 49086 46734 49138
rect 46786 49086 46900 49138
rect 46732 49084 46900 49086
rect 46956 50370 47012 50382
rect 46956 50318 46958 50370
rect 47010 50318 47012 50370
rect 46732 49074 46788 49084
rect 45276 48178 45332 48188
rect 45612 47346 45668 47358
rect 45612 47294 45614 47346
rect 45666 47294 45668 47346
rect 45276 47012 45332 47022
rect 45052 46564 45108 46574
rect 45052 45890 45108 46508
rect 45052 45838 45054 45890
rect 45106 45838 45108 45890
rect 45052 45826 45108 45838
rect 45276 45890 45332 46956
rect 45276 45838 45278 45890
rect 45330 45838 45332 45890
rect 45276 45444 45332 45838
rect 45388 46676 45444 46686
rect 45388 45892 45444 46620
rect 45500 45892 45556 45902
rect 45388 45890 45556 45892
rect 45388 45838 45502 45890
rect 45554 45838 45556 45890
rect 45388 45836 45556 45838
rect 45500 45826 45556 45836
rect 45388 45668 45444 45678
rect 45612 45668 45668 47294
rect 45948 47012 46004 47022
rect 45948 46898 46004 46956
rect 45948 46846 45950 46898
rect 46002 46846 46004 46898
rect 45948 46834 46004 46846
rect 46172 46786 46228 46798
rect 46172 46734 46174 46786
rect 46226 46734 46228 46786
rect 45724 46676 45780 46686
rect 45724 46582 45780 46620
rect 45836 46564 45892 46574
rect 45836 46470 45892 46508
rect 45388 45666 45668 45668
rect 45388 45614 45390 45666
rect 45442 45614 45668 45666
rect 45388 45612 45668 45614
rect 45948 45668 46004 45678
rect 46172 45668 46228 46734
rect 45948 45666 46228 45668
rect 45948 45614 45950 45666
rect 46002 45614 46228 45666
rect 45948 45612 46228 45614
rect 45388 45602 45444 45612
rect 45276 45388 45444 45444
rect 44940 44818 44996 44828
rect 45388 44546 45444 45388
rect 45388 44494 45390 44546
rect 45442 44494 45444 44546
rect 45388 44482 45444 44494
rect 43596 44436 43652 44446
rect 43596 44434 44100 44436
rect 43596 44382 43598 44434
rect 43650 44382 44100 44434
rect 43596 44380 44100 44382
rect 43596 44370 43652 44380
rect 43932 44210 43988 44222
rect 43932 44158 43934 44210
rect 43986 44158 43988 44210
rect 43372 44100 43428 44110
rect 43036 43428 43092 43438
rect 43036 41300 43092 43372
rect 43372 41636 43428 44044
rect 43932 43708 43988 44158
rect 43708 43652 43988 43708
rect 44044 44210 44100 44380
rect 45500 44434 45556 44446
rect 45500 44382 45502 44434
rect 45554 44382 45556 44434
rect 44268 44324 44324 44334
rect 44716 44324 44772 44334
rect 44268 44322 44772 44324
rect 44268 44270 44270 44322
rect 44322 44270 44718 44322
rect 44770 44270 44772 44322
rect 44268 44268 44772 44270
rect 44268 44258 44324 44268
rect 44716 44258 44772 44268
rect 44044 44158 44046 44210
rect 44098 44158 44100 44210
rect 43484 42980 43540 42990
rect 43708 42980 43764 43652
rect 44044 43092 44100 44158
rect 45276 43538 45332 43550
rect 45276 43486 45278 43538
rect 45330 43486 45332 43538
rect 44940 43428 44996 43438
rect 45276 43428 45332 43486
rect 44996 43372 45332 43428
rect 44940 43334 44996 43372
rect 43540 42924 43764 42980
rect 43932 43036 44100 43092
rect 43484 41858 43540 42924
rect 43932 42644 43988 43036
rect 44156 42980 44212 42990
rect 44156 42866 44212 42924
rect 44156 42814 44158 42866
rect 44210 42814 44212 42866
rect 44156 42802 44212 42814
rect 43820 42642 43988 42644
rect 43820 42590 43934 42642
rect 43986 42590 43988 42642
rect 43820 42588 43988 42590
rect 43820 41970 43876 42588
rect 43932 42578 43988 42588
rect 45164 42532 45220 42542
rect 45276 42532 45332 42542
rect 45164 42530 45276 42532
rect 45164 42478 45166 42530
rect 45218 42478 45276 42530
rect 45164 42476 45276 42478
rect 45164 42466 45220 42476
rect 43820 41918 43822 41970
rect 43874 41918 43876 41970
rect 43820 41906 43876 41918
rect 43932 42420 43988 42430
rect 43484 41806 43486 41858
rect 43538 41806 43540 41858
rect 43484 41794 43540 41806
rect 43820 41748 43876 41758
rect 43932 41748 43988 42364
rect 43820 41746 43988 41748
rect 43820 41694 43822 41746
rect 43874 41694 43988 41746
rect 43820 41692 43988 41694
rect 44492 41972 44548 41982
rect 44492 41858 44548 41916
rect 44492 41806 44494 41858
rect 44546 41806 44548 41858
rect 43820 41682 43876 41692
rect 44492 41636 44548 41806
rect 43372 41580 43652 41636
rect 43484 41300 43540 41310
rect 43036 41298 43540 41300
rect 43036 41246 43486 41298
rect 43538 41246 43540 41298
rect 43036 41244 43540 41246
rect 43036 41186 43092 41244
rect 43036 41134 43038 41186
rect 43090 41134 43092 41186
rect 43036 41122 43092 41134
rect 43484 40740 43540 41244
rect 43484 40674 43540 40684
rect 43484 40516 43540 40526
rect 43596 40516 43652 41580
rect 44044 41580 44548 41636
rect 44044 40964 44100 41580
rect 44156 41412 44212 41422
rect 45164 41412 45220 41422
rect 44156 41410 45220 41412
rect 44156 41358 44158 41410
rect 44210 41358 45166 41410
rect 45218 41358 45220 41410
rect 44156 41356 45220 41358
rect 44156 41346 44212 41356
rect 45164 41346 45220 41356
rect 44268 41074 44324 41086
rect 44268 41022 44270 41074
rect 44322 41022 44324 41074
rect 44156 40964 44212 40974
rect 44044 40962 44212 40964
rect 44044 40910 44158 40962
rect 44210 40910 44212 40962
rect 44044 40908 44212 40910
rect 43484 40514 43652 40516
rect 43484 40462 43486 40514
rect 43538 40462 43652 40514
rect 43484 40460 43652 40462
rect 43484 40450 43540 40460
rect 43820 40402 43876 40414
rect 43820 40350 43822 40402
rect 43874 40350 43876 40402
rect 43708 40290 43764 40302
rect 43708 40238 43710 40290
rect 43762 40238 43764 40290
rect 43372 39620 43428 39630
rect 43708 39620 43764 40238
rect 43820 40180 43876 40350
rect 43876 40124 43988 40180
rect 43820 40114 43876 40124
rect 43428 39564 43764 39620
rect 43820 39620 43876 39630
rect 43932 39620 43988 40124
rect 43820 39618 43988 39620
rect 43820 39566 43822 39618
rect 43874 39566 43988 39618
rect 43820 39564 43988 39566
rect 43372 39526 43428 39564
rect 43820 39554 43876 39564
rect 44156 39396 44212 40908
rect 44268 40404 44324 41022
rect 45164 41076 45220 41086
rect 45276 41076 45332 42476
rect 45500 42420 45556 44382
rect 45612 44322 45668 44334
rect 45612 44270 45614 44322
rect 45666 44270 45668 44322
rect 45612 42980 45668 44270
rect 45612 42886 45668 42924
rect 45612 42756 45668 42766
rect 45612 42642 45668 42700
rect 45612 42590 45614 42642
rect 45666 42590 45668 42642
rect 45612 42578 45668 42590
rect 45724 42642 45780 42654
rect 45724 42590 45726 42642
rect 45778 42590 45780 42642
rect 45500 42354 45556 42364
rect 45724 41860 45780 42590
rect 45948 42532 46004 45612
rect 46956 44548 47012 50318
rect 47068 50370 47124 50382
rect 47516 50372 47908 50428
rect 47068 50318 47070 50370
rect 47122 50318 47124 50370
rect 47068 50036 47124 50318
rect 47068 49980 47348 50036
rect 47292 49922 47348 49980
rect 49868 49924 49924 58828
rect 50428 56980 50484 59388
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50316 56978 50484 56980
rect 50316 56926 50430 56978
rect 50482 56926 50484 56978
rect 50316 56924 50484 56926
rect 49980 56868 50036 56878
rect 50316 56868 50372 56924
rect 50428 56914 50484 56924
rect 49980 56866 50372 56868
rect 49980 56814 49982 56866
rect 50034 56814 50372 56866
rect 49980 56812 50372 56814
rect 49980 56802 50036 56812
rect 49980 56308 50036 56318
rect 49980 56214 50036 56252
rect 50316 56308 50372 56812
rect 50988 56756 51044 59500
rect 50316 56242 50372 56252
rect 50428 56700 51044 56756
rect 51100 57540 51156 57550
rect 50316 56084 50372 56094
rect 50316 55990 50372 56028
rect 49980 55188 50036 55198
rect 49980 55094 50036 55132
rect 50316 55074 50372 55086
rect 50316 55022 50318 55074
rect 50370 55022 50372 55074
rect 50316 54516 50372 55022
rect 50316 54450 50372 54460
rect 50428 55076 50484 56700
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50876 56308 50932 56318
rect 50876 56082 50932 56252
rect 50876 56030 50878 56082
rect 50930 56030 50932 56082
rect 50876 55468 50932 56030
rect 50876 55412 51044 55468
rect 50428 51940 50484 55020
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50876 54516 50932 54526
rect 50876 54422 50932 54460
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50988 53060 51044 55412
rect 50764 53004 50988 53060
rect 51100 53060 51156 57484
rect 51212 54626 51268 59948
rect 51436 59444 51492 59454
rect 51436 59218 51492 59388
rect 51436 59166 51438 59218
rect 51490 59166 51492 59218
rect 51436 59154 51492 59166
rect 51548 57876 51604 60732
rect 51660 60722 51716 60732
rect 51660 60004 51716 60014
rect 51772 60004 51828 63084
rect 52108 62580 52164 64428
rect 52332 64146 52388 65436
rect 54124 65380 54180 65390
rect 54124 65286 54180 65324
rect 52780 64484 52836 64494
rect 52780 64390 52836 64428
rect 54012 64484 54068 64494
rect 54012 64390 54068 64428
rect 54348 64482 54404 64494
rect 54348 64430 54350 64482
rect 54402 64430 54404 64482
rect 52332 64094 52334 64146
rect 52386 64094 52388 64146
rect 52332 64082 52388 64094
rect 54124 63924 54180 63934
rect 53564 63922 54180 63924
rect 53564 63870 54126 63922
rect 54178 63870 54180 63922
rect 53564 63868 54180 63870
rect 53564 63362 53620 63868
rect 54124 63858 54180 63868
rect 53564 63310 53566 63362
rect 53618 63310 53620 63362
rect 53564 63298 53620 63310
rect 53004 63252 53060 63262
rect 53900 63252 53956 63262
rect 53060 63196 53172 63252
rect 53004 63158 53060 63196
rect 52108 62486 52164 62524
rect 52444 62468 52500 62478
rect 52444 62374 52500 62412
rect 52892 62244 52948 62254
rect 52780 61684 52836 61694
rect 52892 61684 52948 62188
rect 52780 61682 52948 61684
rect 52780 61630 52782 61682
rect 52834 61630 52948 61682
rect 52780 61628 52948 61630
rect 52780 60676 52836 61628
rect 53116 61570 53172 63196
rect 53900 63158 53956 63196
rect 53228 63138 53284 63150
rect 53228 63086 53230 63138
rect 53282 63086 53284 63138
rect 53228 62468 53284 63086
rect 53228 62402 53284 62412
rect 54124 63138 54180 63150
rect 54124 63086 54126 63138
rect 54178 63086 54180 63138
rect 53116 61518 53118 61570
rect 53170 61518 53172 61570
rect 53116 61506 53172 61518
rect 53452 62354 53508 62366
rect 53452 62302 53454 62354
rect 53506 62302 53508 62354
rect 53004 60788 53060 60798
rect 53004 60694 53060 60732
rect 53340 60788 53396 60798
rect 53452 60788 53508 62302
rect 54124 62244 54180 63086
rect 54124 62178 54180 62188
rect 54348 61570 54404 64430
rect 54460 63588 54516 66220
rect 55020 66210 55076 66220
rect 54908 65490 54964 65502
rect 54908 65438 54910 65490
rect 54962 65438 54964 65490
rect 54908 65380 54964 65438
rect 54908 65314 54964 65324
rect 55020 65492 55076 65502
rect 54572 64706 54628 64718
rect 54572 64654 54574 64706
rect 54626 64654 54628 64706
rect 54572 64148 54628 64654
rect 54572 64054 54628 64092
rect 54908 64484 54964 64494
rect 54796 63922 54852 63934
rect 54796 63870 54798 63922
rect 54850 63870 54852 63922
rect 54684 63812 54740 63822
rect 54684 63718 54740 63756
rect 54460 63522 54516 63532
rect 54460 63364 54516 63374
rect 54796 63364 54852 63870
rect 54460 63362 54852 63364
rect 54460 63310 54462 63362
rect 54514 63310 54852 63362
rect 54460 63308 54852 63310
rect 54460 63298 54516 63308
rect 54348 61518 54350 61570
rect 54402 61518 54404 61570
rect 54348 61506 54404 61518
rect 54908 63250 54964 64428
rect 55020 64036 55076 65436
rect 55020 63970 55076 63980
rect 55132 63812 55188 69200
rect 56028 66500 56084 66510
rect 56028 66406 56084 66444
rect 57148 65492 57204 69200
rect 58156 66164 58212 66174
rect 57820 65602 57876 65614
rect 57820 65550 57822 65602
rect 57874 65550 57876 65602
rect 57148 65426 57204 65436
rect 57596 65492 57652 65502
rect 57596 65398 57652 65436
rect 55356 65380 55412 65390
rect 55244 64932 55300 64942
rect 55244 64818 55300 64876
rect 55244 64766 55246 64818
rect 55298 64766 55300 64818
rect 55244 64754 55300 64766
rect 55356 64484 55412 65324
rect 55468 65378 55524 65390
rect 55468 65326 55470 65378
rect 55522 65326 55524 65378
rect 55468 65268 55524 65326
rect 55468 65202 55524 65212
rect 57372 64596 57428 64606
rect 57372 64594 57540 64596
rect 57372 64542 57374 64594
rect 57426 64542 57540 64594
rect 57372 64540 57540 64542
rect 57372 64530 57428 64540
rect 55356 64418 55412 64428
rect 55244 64036 55300 64046
rect 56028 64036 56084 64046
rect 56812 64036 56868 64046
rect 55300 63980 55412 64036
rect 55244 63970 55300 63980
rect 55132 63746 55188 63756
rect 54908 63198 54910 63250
rect 54962 63198 54964 63250
rect 54460 61124 54516 61134
rect 54460 60898 54516 61068
rect 54460 60846 54462 60898
rect 54514 60846 54516 60898
rect 54460 60834 54516 60846
rect 53396 60732 53508 60788
rect 54684 60788 54740 60798
rect 53340 60694 53396 60732
rect 54684 60694 54740 60732
rect 52780 60610 52836 60620
rect 51660 60002 51828 60004
rect 51660 59950 51662 60002
rect 51714 59950 51828 60002
rect 51660 59948 51828 59950
rect 51884 60228 51940 60238
rect 51884 60002 51940 60172
rect 54908 60114 54964 63198
rect 55020 63700 55076 63710
rect 55020 61682 55076 63644
rect 55244 63252 55300 63262
rect 55244 63158 55300 63196
rect 55356 62242 55412 63980
rect 55916 64034 56868 64036
rect 55916 63982 56030 64034
rect 56082 63982 56814 64034
rect 56866 63982 56868 64034
rect 55916 63980 56868 63982
rect 55356 62190 55358 62242
rect 55410 62190 55412 62242
rect 55356 62178 55412 62190
rect 55804 63588 55860 63598
rect 55020 61630 55022 61682
rect 55074 61630 55076 61682
rect 55020 61618 55076 61630
rect 55468 61572 55524 61582
rect 55468 61478 55524 61516
rect 54908 60062 54910 60114
rect 54962 60062 54964 60114
rect 51884 59950 51886 60002
rect 51938 59950 51940 60002
rect 51660 59938 51716 59948
rect 51660 57876 51716 57886
rect 51548 57874 51716 57876
rect 51548 57822 51662 57874
rect 51714 57822 51716 57874
rect 51548 57820 51716 57822
rect 51660 57810 51716 57820
rect 51436 57652 51492 57662
rect 51436 57558 51492 57596
rect 51548 57538 51604 57550
rect 51548 57486 51550 57538
rect 51602 57486 51604 57538
rect 51548 56196 51604 57486
rect 51660 56196 51716 56206
rect 51548 56194 51716 56196
rect 51548 56142 51662 56194
rect 51714 56142 51716 56194
rect 51548 56140 51716 56142
rect 51660 56130 51716 56140
rect 51436 56084 51492 56094
rect 51212 54574 51214 54626
rect 51266 54574 51268 54626
rect 51212 53396 51268 54574
rect 51324 54740 51380 54750
rect 51324 53508 51380 54684
rect 51436 53732 51492 56028
rect 51884 56084 51940 59950
rect 52108 60004 52164 60014
rect 52108 59910 52164 59948
rect 53340 60004 53396 60014
rect 51996 59778 52052 59790
rect 51996 59726 51998 59778
rect 52050 59726 52052 59778
rect 51996 58546 52052 59726
rect 52108 59106 52164 59118
rect 52108 59054 52110 59106
rect 52162 59054 52164 59106
rect 52108 58658 52164 59054
rect 52108 58606 52110 58658
rect 52162 58606 52164 58658
rect 52108 58594 52164 58606
rect 51996 58494 51998 58546
rect 52050 58494 52052 58546
rect 51996 58482 52052 58494
rect 53004 58434 53060 58446
rect 53004 58382 53006 58434
rect 53058 58382 53060 58434
rect 52556 58324 52612 58334
rect 52556 57874 52612 58268
rect 53004 58324 53060 58382
rect 53004 58258 53060 58268
rect 52556 57822 52558 57874
rect 52610 57822 52612 57874
rect 52556 57810 52612 57822
rect 51996 57650 52052 57662
rect 51996 57598 51998 57650
rect 52050 57598 52052 57650
rect 51996 56532 52052 57598
rect 51996 56466 52052 56476
rect 52780 56532 52836 56542
rect 51884 56018 51940 56028
rect 52780 55410 52836 56476
rect 52780 55358 52782 55410
rect 52834 55358 52836 55410
rect 52780 55346 52836 55358
rect 53340 55298 53396 59948
rect 54236 60004 54292 60014
rect 54908 60004 54964 60062
rect 55244 61124 55300 61134
rect 55244 60114 55300 61068
rect 55804 60898 55860 63532
rect 55804 60846 55806 60898
rect 55858 60846 55860 60898
rect 55804 60834 55860 60846
rect 55244 60062 55246 60114
rect 55298 60062 55300 60114
rect 55244 60050 55300 60062
rect 54236 59106 54292 59948
rect 54236 59054 54238 59106
rect 54290 59054 54292 59106
rect 54236 59042 54292 59054
rect 54684 59948 54908 60004
rect 54684 59444 54740 59948
rect 54908 59938 54964 59948
rect 55916 59444 55972 63980
rect 56028 63970 56084 63980
rect 56812 63970 56868 63980
rect 56364 63812 56420 63822
rect 56364 61794 56420 63756
rect 56588 63700 56644 63710
rect 56588 63606 56644 63644
rect 56924 63700 56980 63710
rect 56924 63698 57428 63700
rect 56924 63646 56926 63698
rect 56978 63646 57428 63698
rect 56924 63644 57428 63646
rect 56924 63634 56980 63644
rect 56700 63588 56756 63598
rect 56700 62354 56756 63532
rect 57372 63250 57428 63644
rect 57372 63198 57374 63250
rect 57426 63198 57428 63250
rect 57372 63186 57428 63198
rect 57484 62804 57540 64540
rect 57036 62748 57540 62804
rect 56700 62302 56702 62354
rect 56754 62302 56756 62354
rect 56700 62290 56756 62302
rect 56924 62466 56980 62478
rect 56924 62414 56926 62466
rect 56978 62414 56980 62466
rect 56364 61742 56366 61794
rect 56418 61742 56420 61794
rect 56364 61730 56420 61742
rect 56924 60900 56980 62414
rect 57036 61010 57092 62748
rect 57372 62466 57428 62478
rect 57372 62414 57374 62466
rect 57426 62414 57428 62466
rect 57036 60958 57038 61010
rect 57090 60958 57092 61010
rect 57036 60946 57092 60958
rect 57148 62354 57204 62366
rect 57148 62302 57150 62354
rect 57202 62302 57204 62354
rect 56924 60834 56980 60844
rect 57148 60898 57204 62302
rect 57372 61124 57428 62414
rect 57372 61058 57428 61068
rect 57484 62354 57540 62366
rect 57484 62302 57486 62354
rect 57538 62302 57540 62354
rect 57148 60846 57150 60898
rect 57202 60846 57204 60898
rect 57148 60834 57204 60846
rect 57372 60900 57428 60910
rect 57372 60806 57428 60844
rect 56700 60786 56756 60798
rect 56700 60734 56702 60786
rect 56754 60734 56756 60786
rect 56028 60676 56084 60686
rect 56028 60674 56532 60676
rect 56028 60622 56030 60674
rect 56082 60622 56532 60674
rect 56028 60620 56532 60622
rect 56028 60610 56084 60620
rect 56028 59444 56084 59454
rect 55916 59388 56028 59444
rect 54684 58548 54740 59388
rect 56028 59350 56084 59388
rect 56476 59220 56532 60620
rect 56588 59220 56644 59230
rect 56476 59218 56644 59220
rect 56476 59166 56590 59218
rect 56642 59166 56644 59218
rect 56476 59164 56644 59166
rect 56588 59154 56644 59164
rect 55580 59106 55636 59118
rect 55580 59054 55582 59106
rect 55634 59054 55636 59106
rect 55580 58994 55636 59054
rect 55580 58942 55582 58994
rect 55634 58942 55636 58994
rect 55580 58930 55636 58942
rect 56140 58994 56196 59006
rect 56140 58942 56142 58994
rect 56194 58942 56196 58994
rect 54236 58546 54740 58548
rect 54236 58494 54686 58546
rect 54738 58494 54740 58546
rect 54236 58492 54740 58494
rect 56140 58548 56196 58942
rect 56700 58548 56756 60734
rect 57484 60788 57540 62302
rect 57708 60788 57764 60798
rect 57484 60732 57708 60788
rect 57820 60788 57876 65550
rect 58156 65492 58212 66108
rect 58156 65398 58212 65436
rect 58044 64706 58100 64718
rect 58044 64654 58046 64706
rect 58098 64654 58100 64706
rect 58044 64484 58100 64654
rect 58044 63138 58100 64428
rect 58044 63086 58046 63138
rect 58098 63086 58100 63138
rect 58044 63074 58100 63086
rect 57932 61124 57988 61134
rect 57932 61010 57988 61068
rect 57932 60958 57934 61010
rect 57986 60958 57988 61010
rect 57932 60946 57988 60958
rect 57820 60732 57988 60788
rect 57708 60694 57764 60732
rect 56924 60564 56980 60574
rect 56924 60470 56980 60508
rect 57372 59892 57428 59902
rect 56812 59890 57428 59892
rect 56812 59838 57374 59890
rect 57426 59838 57428 59890
rect 56812 59836 57428 59838
rect 56812 59442 56868 59836
rect 57372 59826 57428 59836
rect 56812 59390 56814 59442
rect 56866 59390 56868 59442
rect 56812 59378 56868 59390
rect 56924 59444 56980 59454
rect 56924 59330 56980 59388
rect 56924 59278 56926 59330
rect 56978 59278 56980 59330
rect 56924 59266 56980 59278
rect 57708 59108 57764 59118
rect 57708 59106 57876 59108
rect 57708 59054 57710 59106
rect 57762 59054 57876 59106
rect 57708 59052 57876 59054
rect 57708 59042 57764 59052
rect 56140 58492 56756 58548
rect 54236 56308 54292 58492
rect 54684 58482 54740 58492
rect 55356 56980 55412 56990
rect 53900 56306 54292 56308
rect 53900 56254 54238 56306
rect 54290 56254 54292 56306
rect 53900 56252 54292 56254
rect 53340 55246 53342 55298
rect 53394 55246 53396 55298
rect 53340 55234 53396 55246
rect 53788 55970 53844 55982
rect 53788 55918 53790 55970
rect 53842 55918 53844 55970
rect 52780 55074 52836 55086
rect 52780 55022 52782 55074
rect 52834 55022 52836 55074
rect 51884 54740 51940 54750
rect 51884 54646 51940 54684
rect 51660 54516 51716 54526
rect 51660 53956 51716 54460
rect 51660 53890 51716 53900
rect 52668 53956 52724 53966
rect 52668 53862 52724 53900
rect 52780 53844 52836 55022
rect 52892 55076 52948 55086
rect 52892 54982 52948 55020
rect 53116 55074 53172 55086
rect 53116 55022 53118 55074
rect 53170 55022 53172 55074
rect 53116 54740 53172 55022
rect 53116 54674 53172 54684
rect 53788 55076 53844 55918
rect 53004 53844 53060 53854
rect 52780 53778 52836 53788
rect 52892 53788 53004 53844
rect 51436 53730 51940 53732
rect 51436 53678 51438 53730
rect 51490 53678 51940 53730
rect 51436 53676 51940 53678
rect 51436 53666 51492 53676
rect 51660 53508 51716 53518
rect 51324 53452 51604 53508
rect 51212 53340 51380 53396
rect 51100 53004 51268 53060
rect 50764 52948 50820 53004
rect 50988 52966 51044 53004
rect 50540 52946 50820 52948
rect 50540 52894 50766 52946
rect 50818 52894 50820 52946
rect 50540 52892 50820 52894
rect 50540 52162 50596 52892
rect 50764 52882 50820 52892
rect 51212 52274 51268 53004
rect 51324 52724 51380 53340
rect 51548 53172 51604 53452
rect 51660 53414 51716 53452
rect 51548 53058 51604 53116
rect 51548 53006 51550 53058
rect 51602 53006 51604 53058
rect 51548 52994 51604 53006
rect 51660 53060 51716 53070
rect 51716 53004 51828 53060
rect 51660 52994 51716 53004
rect 51324 52658 51380 52668
rect 51212 52222 51214 52274
rect 51266 52222 51268 52274
rect 50540 52110 50542 52162
rect 50594 52110 50596 52162
rect 50540 52098 50596 52110
rect 50988 52162 51044 52174
rect 50988 52110 50990 52162
rect 51042 52110 51044 52162
rect 50988 51940 51044 52110
rect 50428 51884 51044 51940
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 47292 49870 47294 49922
rect 47346 49870 47348 49922
rect 47292 49858 47348 49870
rect 48972 49868 49924 49924
rect 50428 50316 50932 50372
rect 47404 49588 47460 49598
rect 47404 49494 47460 49532
rect 48860 49588 48916 49598
rect 48860 49138 48916 49532
rect 48860 49086 48862 49138
rect 48914 49086 48916 49138
rect 48860 49074 48916 49086
rect 47964 48132 48020 48142
rect 47740 47570 47796 47582
rect 47740 47518 47742 47570
rect 47794 47518 47796 47570
rect 47740 47236 47796 47518
rect 47740 47170 47796 47180
rect 47628 46900 47684 46910
rect 47628 46674 47684 46844
rect 47628 46622 47630 46674
rect 47682 46622 47684 46674
rect 47628 46564 47684 46622
rect 47628 46498 47684 46508
rect 47852 46452 47908 46462
rect 46508 44492 47124 44548
rect 46508 44322 46564 44492
rect 46508 44270 46510 44322
rect 46562 44270 46564 44322
rect 46508 44258 46564 44270
rect 46732 44380 47012 44436
rect 46620 44098 46676 44110
rect 46620 44046 46622 44098
rect 46674 44046 46676 44098
rect 46620 43708 46676 44046
rect 46060 43652 46676 43708
rect 46060 43650 46116 43652
rect 46060 43598 46062 43650
rect 46114 43598 46116 43650
rect 46060 43586 46116 43598
rect 46620 43428 46676 43438
rect 46620 42756 46676 43372
rect 46732 42866 46788 44380
rect 46956 44322 47012 44380
rect 46956 44270 46958 44322
rect 47010 44270 47012 44322
rect 46956 44258 47012 44270
rect 46844 44210 46900 44222
rect 46844 44158 46846 44210
rect 46898 44158 46900 44210
rect 46844 43428 46900 44158
rect 47068 44100 47124 44492
rect 46844 43362 46900 43372
rect 46956 44044 47124 44100
rect 46732 42814 46734 42866
rect 46786 42814 46788 42866
rect 46732 42802 46788 42814
rect 46620 42662 46676 42700
rect 45948 42466 46004 42476
rect 46396 42532 46452 42542
rect 46396 42438 46452 42476
rect 46844 42532 46900 42542
rect 46956 42532 47012 44044
rect 46844 42530 47012 42532
rect 46844 42478 46846 42530
rect 46898 42478 47012 42530
rect 46844 42476 47012 42478
rect 45724 41794 45780 41804
rect 46844 41860 46900 42476
rect 46844 41794 46900 41804
rect 45500 41300 45556 41310
rect 45500 41298 46004 41300
rect 45500 41246 45502 41298
rect 45554 41246 46004 41298
rect 45500 41244 46004 41246
rect 45500 41234 45556 41244
rect 45220 41020 45332 41076
rect 45164 41010 45220 41020
rect 45388 40964 45444 40974
rect 45276 40962 45444 40964
rect 45276 40910 45390 40962
rect 45442 40910 45444 40962
rect 45276 40908 45444 40910
rect 45164 40740 45220 40750
rect 44716 40404 44772 40414
rect 45164 40404 45220 40684
rect 44268 40402 44772 40404
rect 44268 40350 44718 40402
rect 44770 40350 44772 40402
rect 44268 40348 44772 40350
rect 44716 39844 44772 40348
rect 44716 39778 44772 39788
rect 44828 40402 45220 40404
rect 44828 40350 45166 40402
rect 45218 40350 45220 40402
rect 44828 40348 45220 40350
rect 44268 39508 44324 39518
rect 44268 39414 44324 39452
rect 43708 39340 44212 39396
rect 43036 37156 43092 37166
rect 43036 37062 43092 37100
rect 42700 36866 42756 36876
rect 42588 35186 42644 35196
rect 42700 35586 42756 35598
rect 42700 35534 42702 35586
rect 42754 35534 42756 35586
rect 42700 34468 42756 35534
rect 43708 35252 43764 39340
rect 44828 39060 44884 40348
rect 45164 40338 45220 40348
rect 45276 39730 45332 40908
rect 45388 40898 45444 40908
rect 45948 40514 46004 41244
rect 45948 40462 45950 40514
rect 46002 40462 46004 40514
rect 45948 40450 46004 40462
rect 47740 40292 47796 40302
rect 47516 40236 47740 40292
rect 47404 40180 47460 40190
rect 45836 39844 45892 39854
rect 45836 39750 45892 39788
rect 47404 39842 47460 40124
rect 47404 39790 47406 39842
rect 47458 39790 47460 39842
rect 47404 39778 47460 39790
rect 45276 39678 45278 39730
rect 45330 39678 45332 39730
rect 45276 39666 45332 39678
rect 47516 39730 47572 40236
rect 47740 40226 47796 40236
rect 47516 39678 47518 39730
rect 47570 39678 47572 39730
rect 47516 39666 47572 39678
rect 45388 39618 45444 39630
rect 45388 39566 45390 39618
rect 45442 39566 45444 39618
rect 45052 39508 45108 39518
rect 45052 39414 45108 39452
rect 45388 39284 45444 39566
rect 45724 39508 45780 39518
rect 45724 39414 45780 39452
rect 45836 39394 45892 39406
rect 45836 39342 45838 39394
rect 45890 39342 45892 39394
rect 45836 39284 45892 39342
rect 45388 39228 45892 39284
rect 44268 39058 44884 39060
rect 44268 39006 44830 39058
rect 44882 39006 44884 39058
rect 44268 39004 44884 39006
rect 44268 37492 44324 39004
rect 44828 38994 44884 39004
rect 45836 38948 45892 39228
rect 45836 38892 46340 38948
rect 45948 38724 46004 38734
rect 45724 38722 46004 38724
rect 45724 38670 45950 38722
rect 46002 38670 46004 38722
rect 45724 38668 46004 38670
rect 45724 38164 45780 38668
rect 45948 38658 46004 38668
rect 46172 38724 46228 38734
rect 46172 38630 46228 38668
rect 46284 38668 46340 38892
rect 46284 38612 46564 38668
rect 46508 38610 46676 38612
rect 46508 38558 46510 38610
rect 46562 38558 46676 38610
rect 46508 38556 46676 38558
rect 46508 38546 46564 38556
rect 45388 38052 45444 38062
rect 43820 37490 44324 37492
rect 43820 37438 44270 37490
rect 44322 37438 44324 37490
rect 43820 37436 44324 37438
rect 43820 37266 43876 37436
rect 44268 37426 44324 37436
rect 45276 38050 45444 38052
rect 45276 37998 45390 38050
rect 45442 37998 45444 38050
rect 45276 37996 45444 37998
rect 45724 38052 45780 38108
rect 46396 38164 46452 38174
rect 46396 38070 46452 38108
rect 45836 38052 45892 38062
rect 45724 38050 45892 38052
rect 45724 37998 45838 38050
rect 45890 37998 45892 38050
rect 45724 37996 45892 37998
rect 45276 37826 45332 37996
rect 45388 37986 45444 37996
rect 45836 37986 45892 37996
rect 46060 38052 46116 38062
rect 46060 37938 46116 37996
rect 46060 37886 46062 37938
rect 46114 37886 46116 37938
rect 46060 37874 46116 37886
rect 46508 37940 46564 37950
rect 45276 37774 45278 37826
rect 45330 37774 45332 37826
rect 43820 37214 43822 37266
rect 43874 37214 43876 37266
rect 43820 37202 43876 37214
rect 44044 36372 44100 36382
rect 44044 36370 44996 36372
rect 44044 36318 44046 36370
rect 44098 36318 44996 36370
rect 44044 36316 44996 36318
rect 44044 36306 44100 36316
rect 43820 36258 43876 36270
rect 43820 36206 43822 36258
rect 43874 36206 43876 36258
rect 43820 35476 43876 36206
rect 43932 36258 43988 36270
rect 43932 36206 43934 36258
rect 43986 36206 43988 36258
rect 43932 35924 43988 36206
rect 43932 35868 44884 35924
rect 44828 35810 44884 35868
rect 44828 35758 44830 35810
rect 44882 35758 44884 35810
rect 44828 35746 44884 35758
rect 43820 35420 44100 35476
rect 43708 35186 43764 35196
rect 44044 35026 44100 35420
rect 44716 35252 44772 35262
rect 44772 35196 44884 35252
rect 44716 35186 44772 35196
rect 44044 34974 44046 35026
rect 44098 34974 44100 35026
rect 44044 34962 44100 34974
rect 43932 34916 43988 34954
rect 43932 34850 43988 34860
rect 44268 34916 44324 34926
rect 42700 34402 42756 34412
rect 43596 34802 43652 34814
rect 44156 34804 44212 34814
rect 43596 34750 43598 34802
rect 43650 34750 43652 34802
rect 43596 34468 43652 34750
rect 43596 34402 43652 34412
rect 44044 34802 44212 34804
rect 44044 34750 44158 34802
rect 44210 34750 44212 34802
rect 44044 34748 44212 34750
rect 44044 34356 44100 34748
rect 44156 34738 44212 34748
rect 43708 34300 44100 34356
rect 44268 34354 44324 34860
rect 44828 34804 44884 35196
rect 44940 35138 44996 36316
rect 44940 35086 44942 35138
rect 44994 35086 44996 35138
rect 44940 35074 44996 35086
rect 44940 34804 44996 34814
rect 44828 34802 44996 34804
rect 44828 34750 44942 34802
rect 44994 34750 44996 34802
rect 44828 34748 44996 34750
rect 44940 34738 44996 34748
rect 45052 34802 45108 34814
rect 45052 34750 45054 34802
rect 45106 34750 45108 34802
rect 44268 34302 44270 34354
rect 44322 34302 44324 34354
rect 43372 33236 43428 33246
rect 43708 33236 43764 34300
rect 44268 34290 44324 34302
rect 44492 34468 44548 34478
rect 44492 34354 44548 34412
rect 44492 34302 44494 34354
rect 44546 34302 44548 34354
rect 44492 34290 44548 34302
rect 43932 34130 43988 34142
rect 43932 34078 43934 34130
rect 43986 34078 43988 34130
rect 43932 33348 43988 34078
rect 44604 34132 44660 34142
rect 44604 34038 44660 34076
rect 45052 34132 45108 34750
rect 45052 34066 45108 34076
rect 43428 33234 43764 33236
rect 43428 33182 43710 33234
rect 43762 33182 43764 33234
rect 43428 33180 43764 33182
rect 43372 32786 43428 33180
rect 43708 33170 43764 33180
rect 43820 33346 43988 33348
rect 43820 33294 43934 33346
rect 43986 33294 43988 33346
rect 43820 33292 43988 33294
rect 43372 32734 43374 32786
rect 43426 32734 43428 32786
rect 43372 32722 43428 32734
rect 43596 32452 43652 32462
rect 43596 32358 43652 32396
rect 42140 31890 42532 31892
rect 42140 31838 42142 31890
rect 42194 31838 42532 31890
rect 42140 31836 42532 31838
rect 42588 32340 42644 32350
rect 43260 32340 43316 32350
rect 42140 31826 42196 31836
rect 42364 30994 42420 31836
rect 42364 30942 42366 30994
rect 42418 30942 42420 30994
rect 41692 30884 41748 30894
rect 41468 29316 41524 29326
rect 41468 28754 41524 29260
rect 41468 28702 41470 28754
rect 41522 28702 41524 28754
rect 41468 28690 41524 28702
rect 40908 28532 40964 28542
rect 40908 27188 40964 28476
rect 41132 27860 41188 27870
rect 41132 27766 41188 27804
rect 40908 27074 40964 27132
rect 40908 27022 40910 27074
rect 40962 27022 40964 27074
rect 40908 27010 40964 27022
rect 40460 26852 40852 26908
rect 41692 26908 41748 30828
rect 42364 30212 42420 30942
rect 41916 30156 42364 30212
rect 41916 29988 41972 30156
rect 42364 30146 42420 30156
rect 42588 29988 42644 32284
rect 43036 32338 43316 32340
rect 43036 32286 43262 32338
rect 43314 32286 43316 32338
rect 43036 32284 43316 32286
rect 43036 31106 43092 32284
rect 43260 32274 43316 32284
rect 43708 32004 43764 32014
rect 43820 32004 43876 33292
rect 43932 33282 43988 33292
rect 43708 32002 43876 32004
rect 43708 31950 43710 32002
rect 43762 31950 43876 32002
rect 43708 31948 43876 31950
rect 43932 32562 43988 32574
rect 43932 32510 43934 32562
rect 43986 32510 43988 32562
rect 43932 32004 43988 32510
rect 44156 32562 44212 32574
rect 44156 32510 44158 32562
rect 44210 32510 44212 32562
rect 44044 32452 44100 32462
rect 44044 32358 44100 32396
rect 44044 32004 44100 32014
rect 43932 32002 44100 32004
rect 43932 31950 44046 32002
rect 44098 31950 44100 32002
rect 43932 31948 44100 31950
rect 43708 31938 43764 31948
rect 43036 31054 43038 31106
rect 43090 31054 43092 31106
rect 43036 31042 43092 31054
rect 43932 30772 43988 31948
rect 44044 31938 44100 31948
rect 44156 31780 44212 32510
rect 44492 32564 44548 32574
rect 44940 32564 44996 32574
rect 45276 32564 45332 37774
rect 45948 37826 46004 37838
rect 45948 37774 45950 37826
rect 46002 37774 46004 37826
rect 45948 37492 46004 37774
rect 45948 37436 46452 37492
rect 46396 37378 46452 37436
rect 46508 37490 46564 37884
rect 46508 37438 46510 37490
rect 46562 37438 46564 37490
rect 46508 37426 46564 37438
rect 46620 37490 46676 38556
rect 46620 37438 46622 37490
rect 46674 37438 46676 37490
rect 46620 37426 46676 37438
rect 46396 37326 46398 37378
rect 46450 37326 46452 37378
rect 46396 37314 46452 37326
rect 46172 37268 46228 37278
rect 45836 37044 45892 37054
rect 45500 35700 45556 35710
rect 45500 35606 45556 35644
rect 45500 35252 45556 35262
rect 45500 35026 45556 35196
rect 45500 34974 45502 35026
rect 45554 34974 45556 35026
rect 45500 34962 45556 34974
rect 45724 34132 45780 34142
rect 45724 34038 45780 34076
rect 44492 32562 45332 32564
rect 44492 32510 44494 32562
rect 44546 32510 44942 32562
rect 44994 32510 45332 32562
rect 44492 32508 45332 32510
rect 44268 31780 44324 31790
rect 44156 31724 44268 31780
rect 44268 31686 44324 31724
rect 41804 29204 41860 29214
rect 41804 27970 41860 29148
rect 41804 27918 41806 27970
rect 41858 27918 41860 27970
rect 41804 27906 41860 27918
rect 41916 28754 41972 29932
rect 41916 28702 41918 28754
rect 41970 28702 41972 28754
rect 41916 27860 41972 28702
rect 41916 27188 41972 27804
rect 41916 27094 41972 27132
rect 42364 29932 42644 29988
rect 43484 30716 43988 30772
rect 41692 26852 41972 26908
rect 40124 26516 40180 26526
rect 40124 26422 40180 26460
rect 39788 26404 39844 26414
rect 39676 26402 39956 26404
rect 39676 26350 39790 26402
rect 39842 26350 39956 26402
rect 39676 26348 39956 26350
rect 39676 26180 39732 26348
rect 39788 26338 39844 26348
rect 39676 26114 39732 26124
rect 39788 26068 39844 26078
rect 39788 25730 39844 26012
rect 39788 25678 39790 25730
rect 39842 25678 39844 25730
rect 39788 25666 39844 25678
rect 39900 25730 39956 26348
rect 39900 25678 39902 25730
rect 39954 25678 39956 25730
rect 39900 25666 39956 25678
rect 40348 25732 40404 25742
rect 40124 25508 40180 25518
rect 40124 25414 40180 25452
rect 39564 25106 39620 25116
rect 40236 25394 40292 25406
rect 40236 25342 40238 25394
rect 40290 25342 40292 25394
rect 39228 24894 39230 24946
rect 39282 24894 39284 24946
rect 39228 24882 39284 24894
rect 38892 24668 39060 24724
rect 38444 24050 38500 24668
rect 38444 23998 38446 24050
rect 38498 23998 38500 24050
rect 38108 23268 38164 23278
rect 37884 23156 37940 23166
rect 37884 22370 37940 23100
rect 38108 23156 38164 23212
rect 38444 23156 38500 23998
rect 38668 24610 38724 24622
rect 38668 24558 38670 24610
rect 38722 24558 38724 24610
rect 38108 23154 38276 23156
rect 38108 23102 38110 23154
rect 38162 23102 38276 23154
rect 38108 23100 38276 23102
rect 38108 23090 38164 23100
rect 37884 22318 37886 22370
rect 37938 22318 37940 22370
rect 37884 22306 37940 22318
rect 37212 22206 37214 22258
rect 37266 22206 37268 22258
rect 37212 22036 37268 22206
rect 37324 22260 37380 22270
rect 37324 22166 37380 22204
rect 37436 22260 37492 22270
rect 37436 22258 37828 22260
rect 37436 22206 37438 22258
rect 37490 22206 37828 22258
rect 37436 22204 37828 22206
rect 37436 22194 37492 22204
rect 37212 21980 37716 22036
rect 37100 21698 37156 21710
rect 37100 21646 37102 21698
rect 37154 21646 37156 21698
rect 36988 19460 37044 19470
rect 36988 19234 37044 19404
rect 36988 19182 36990 19234
rect 37042 19182 37044 19234
rect 36988 19170 37044 19182
rect 37100 19236 37156 21646
rect 37660 21588 37716 21980
rect 37772 21812 37828 22204
rect 37772 21756 38164 21812
rect 38108 21698 38164 21756
rect 38108 21646 38110 21698
rect 38162 21646 38164 21698
rect 38108 21634 38164 21646
rect 37772 21588 37828 21598
rect 37660 21586 37828 21588
rect 37660 21534 37774 21586
rect 37826 21534 37828 21586
rect 37660 21532 37828 21534
rect 37772 21522 37828 21532
rect 37100 19170 37156 19180
rect 37212 20244 37268 20254
rect 37212 19234 37268 20188
rect 37772 20244 37828 20254
rect 37772 20150 37828 20188
rect 37212 19182 37214 19234
rect 37266 19182 37268 19234
rect 37100 19010 37156 19022
rect 37100 18958 37102 19010
rect 37154 18958 37156 19010
rect 37100 18564 37156 18958
rect 37100 18498 37156 18508
rect 36876 18386 36932 18396
rect 37212 17780 37268 19182
rect 37548 19236 37604 19246
rect 37996 19236 38052 19246
rect 37548 19234 38052 19236
rect 37548 19182 37550 19234
rect 37602 19182 37998 19234
rect 38050 19182 38052 19234
rect 37548 19180 38052 19182
rect 37548 19170 37604 19180
rect 37996 19170 38052 19180
rect 37884 19010 37940 19022
rect 37884 18958 37886 19010
rect 37938 18958 37940 19010
rect 37884 18788 37940 18958
rect 37884 18722 37940 18732
rect 38108 19010 38164 19022
rect 38108 18958 38110 19010
rect 38162 18958 38164 19010
rect 37212 17714 37268 17724
rect 37884 18340 37940 18350
rect 35980 16930 36036 16940
rect 36092 17276 36596 17332
rect 37884 17666 37940 18284
rect 37884 17614 37886 17666
rect 37938 17614 37940 17666
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34972 16324 35028 16334
rect 34972 15314 35028 16268
rect 35644 16210 35700 16222
rect 35644 16158 35646 16210
rect 35698 16158 35700 16210
rect 35532 16100 35588 16110
rect 34972 15262 34974 15314
rect 35026 15262 35028 15314
rect 34972 15148 35028 15262
rect 35308 15986 35364 15998
rect 35308 15934 35310 15986
rect 35362 15934 35364 15986
rect 35308 15148 35364 15934
rect 35532 15986 35588 16044
rect 35532 15934 35534 15986
rect 35586 15934 35588 15986
rect 35532 15922 35588 15934
rect 35644 15426 35700 16158
rect 36092 16210 36148 17276
rect 37884 16324 37940 17614
rect 38108 18338 38164 18958
rect 38108 18286 38110 18338
rect 38162 18286 38164 18338
rect 38108 16660 38164 18286
rect 38108 16594 38164 16604
rect 38220 16436 38276 23100
rect 38444 23090 38500 23100
rect 38556 23154 38612 23166
rect 38556 23102 38558 23154
rect 38610 23102 38612 23154
rect 38332 23042 38388 23054
rect 38332 22990 38334 23042
rect 38386 22990 38388 23042
rect 38332 21586 38388 22990
rect 38556 22596 38612 23102
rect 38556 22530 38612 22540
rect 38556 22370 38612 22382
rect 38556 22318 38558 22370
rect 38610 22318 38612 22370
rect 38444 22260 38500 22270
rect 38556 22260 38612 22318
rect 38500 22204 38612 22260
rect 38444 22194 38500 22204
rect 38668 21924 38724 24558
rect 38780 23154 38836 23166
rect 38780 23102 38782 23154
rect 38834 23102 38836 23154
rect 38780 22484 38836 23102
rect 38780 22418 38836 22428
rect 38332 21534 38334 21586
rect 38386 21534 38388 21586
rect 38332 21522 38388 21534
rect 38556 21868 38724 21924
rect 38556 20244 38612 21868
rect 39004 21812 39060 24668
rect 40236 24052 40292 25342
rect 40236 23986 40292 23996
rect 40012 23716 40068 23726
rect 39228 23268 39284 23278
rect 39228 23174 39284 23212
rect 38556 20178 38612 20188
rect 38668 21756 39060 21812
rect 38332 19012 38388 19022
rect 38556 19012 38612 19022
rect 38332 18918 38388 18956
rect 38444 18956 38556 19012
rect 38668 19012 38724 21756
rect 39004 21586 39060 21598
rect 39004 21534 39006 21586
rect 39058 21534 39060 21586
rect 38780 19572 38836 19582
rect 38780 19234 38836 19516
rect 38780 19182 38782 19234
rect 38834 19182 38836 19234
rect 38780 19170 38836 19182
rect 38892 19012 38948 19022
rect 38668 18956 38836 19012
rect 38444 17780 38500 18956
rect 38556 18946 38612 18956
rect 38556 18340 38612 18350
rect 38556 18246 38612 18284
rect 38556 17780 38612 17790
rect 38444 17778 38612 17780
rect 38444 17726 38558 17778
rect 38610 17726 38612 17778
rect 38444 17724 38612 17726
rect 38556 17714 38612 17724
rect 37884 16258 37940 16268
rect 38108 16380 38276 16436
rect 36092 16158 36094 16210
rect 36146 16158 36148 16210
rect 36092 16100 36148 16158
rect 36092 16034 36148 16044
rect 37772 15988 37828 15998
rect 35644 15374 35646 15426
rect 35698 15374 35700 15426
rect 35644 15362 35700 15374
rect 37548 15764 37604 15774
rect 34972 15092 35140 15148
rect 35308 15092 35588 15148
rect 34860 14130 34916 14140
rect 34972 14530 35028 14542
rect 34972 14478 34974 14530
rect 35026 14478 35028 14530
rect 34300 13806 34302 13858
rect 34354 13806 34356 13858
rect 34300 13794 34356 13806
rect 34524 13916 34916 13972
rect 34524 13858 34580 13916
rect 34524 13806 34526 13858
rect 34578 13806 34580 13858
rect 34524 13794 34580 13806
rect 34748 13746 34804 13758
rect 34748 13694 34750 13746
rect 34802 13694 34804 13746
rect 34076 13634 34132 13646
rect 34748 13636 34804 13694
rect 34076 13582 34078 13634
rect 34130 13582 34132 13634
rect 34076 13524 34132 13582
rect 34188 13580 34804 13636
rect 34188 13524 34244 13580
rect 34076 13468 34244 13524
rect 34636 13412 34692 13580
rect 34860 13412 34916 13916
rect 34524 13356 34692 13412
rect 34748 13356 34916 13412
rect 34972 13634 35028 14478
rect 35084 14084 35140 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14644 35588 15092
rect 35420 14588 35588 14644
rect 37100 14644 37156 14654
rect 35420 14530 35476 14588
rect 35420 14478 35422 14530
rect 35474 14478 35476 14530
rect 35420 14466 35476 14478
rect 35084 14028 35588 14084
rect 35308 13858 35364 13870
rect 35308 13806 35310 13858
rect 35362 13806 35364 13858
rect 34972 13582 34974 13634
rect 35026 13582 35028 13634
rect 33964 13244 34244 13300
rect 33964 13076 34020 13086
rect 33964 12738 34020 13020
rect 33964 12686 33966 12738
rect 34018 12686 34020 12738
rect 33964 12674 34020 12686
rect 33852 12236 34132 12292
rect 33740 12180 33796 12190
rect 33628 12178 33908 12180
rect 33628 12126 33742 12178
rect 33794 12126 33908 12178
rect 33628 12124 33908 12126
rect 33740 12114 33796 12124
rect 33292 11218 33348 11228
rect 33404 11340 33572 11396
rect 32620 10836 32676 10846
rect 32620 9716 32676 10780
rect 33404 10276 33460 11340
rect 33516 11172 33572 11182
rect 33516 10948 33572 11116
rect 33516 10882 33572 10892
rect 33292 10220 33460 10276
rect 32732 10052 32788 10062
rect 32732 10050 33124 10052
rect 32732 9998 32734 10050
rect 32786 9998 33124 10050
rect 32732 9996 33124 9998
rect 32732 9986 32788 9996
rect 32732 9716 32788 9726
rect 32620 9660 32732 9716
rect 32732 9622 32788 9660
rect 32844 9714 32900 9726
rect 32844 9662 32846 9714
rect 32898 9662 32900 9714
rect 32844 9268 32900 9662
rect 32844 9202 32900 9212
rect 32508 8540 32676 8596
rect 32508 8372 32564 8382
rect 31500 8206 31502 8258
rect 31554 8206 31556 8258
rect 31164 8148 31220 8158
rect 31164 8054 31220 8092
rect 31500 7924 31556 8206
rect 32172 8316 32508 8372
rect 32172 8258 32228 8316
rect 32172 8206 32174 8258
rect 32226 8206 32228 8258
rect 32172 8194 32228 8206
rect 31612 8148 31668 8158
rect 31612 8054 31668 8092
rect 30940 7634 30996 7644
rect 31276 7868 31556 7924
rect 31724 8034 31780 8046
rect 31724 7982 31726 8034
rect 31778 7982 31780 8034
rect 31276 6692 31332 7868
rect 31500 7700 31556 7710
rect 31500 7606 31556 7644
rect 31724 7364 31780 7982
rect 31724 7298 31780 7308
rect 31836 7362 31892 7374
rect 31836 7310 31838 7362
rect 31890 7310 31892 7362
rect 31836 6692 31892 7310
rect 32284 6804 32340 8316
rect 32508 8278 32564 8316
rect 31164 6690 31332 6692
rect 31164 6638 31278 6690
rect 31330 6638 31332 6690
rect 31164 6636 31332 6638
rect 30940 6580 30996 6590
rect 31164 6580 31220 6636
rect 31276 6626 31332 6636
rect 31612 6636 31836 6692
rect 30940 6578 31220 6580
rect 30940 6526 30942 6578
rect 30994 6526 31220 6578
rect 30940 6524 31220 6526
rect 30940 6514 30996 6524
rect 30716 6466 30772 6478
rect 30716 6414 30718 6466
rect 30770 6414 30772 6466
rect 30716 6132 30772 6414
rect 30716 6066 30772 6076
rect 30828 6466 30884 6478
rect 30828 6414 30830 6466
rect 30882 6414 30884 6466
rect 30828 6020 30884 6414
rect 31388 6466 31444 6478
rect 31388 6414 31390 6466
rect 31442 6414 31444 6466
rect 31276 6244 31332 6254
rect 30828 5954 30884 5964
rect 31164 6130 31220 6142
rect 31164 6078 31166 6130
rect 31218 6078 31220 6130
rect 30940 5908 30996 5918
rect 30940 5906 31108 5908
rect 30940 5854 30942 5906
rect 30994 5854 31108 5906
rect 30940 5852 31108 5854
rect 30940 5796 30996 5852
rect 30604 5740 30996 5796
rect 30828 5572 30884 5582
rect 30716 5516 30828 5572
rect 30716 5122 30772 5516
rect 30828 5506 30884 5516
rect 31052 5348 31108 5852
rect 31164 5460 31220 6078
rect 31276 6018 31332 6188
rect 31276 5966 31278 6018
rect 31330 5966 31332 6018
rect 31276 5954 31332 5966
rect 31388 5906 31444 6414
rect 31388 5854 31390 5906
rect 31442 5854 31444 5906
rect 31388 5842 31444 5854
rect 31500 6466 31556 6478
rect 31500 6414 31502 6466
rect 31554 6414 31556 6466
rect 31500 5460 31556 6414
rect 31164 5404 31444 5460
rect 31052 5292 31220 5348
rect 30940 5236 30996 5246
rect 30996 5180 31108 5236
rect 30940 5170 30996 5180
rect 30716 5070 30718 5122
rect 30770 5070 30772 5122
rect 30716 5058 30772 5070
rect 30828 5124 30884 5134
rect 30828 5030 30884 5068
rect 31052 5122 31108 5180
rect 31052 5070 31054 5122
rect 31106 5070 31108 5122
rect 31052 5058 31108 5070
rect 31164 5122 31220 5292
rect 31164 5070 31166 5122
rect 31218 5070 31220 5122
rect 31164 5058 31220 5070
rect 30492 4498 30548 4508
rect 31388 4452 31444 5404
rect 31500 5394 31556 5404
rect 31612 5234 31668 6636
rect 31836 6626 31892 6636
rect 31948 6802 32340 6804
rect 31948 6750 32286 6802
rect 32338 6750 32340 6802
rect 31948 6748 32340 6750
rect 31948 6690 32004 6748
rect 32284 6738 32340 6748
rect 31948 6638 31950 6690
rect 32002 6638 32004 6690
rect 31948 6580 32004 6638
rect 32396 6692 32452 6702
rect 32284 6580 32340 6590
rect 31948 6514 32004 6524
rect 32172 6524 32284 6580
rect 32060 6244 32116 6254
rect 32060 6130 32116 6188
rect 32060 6078 32062 6130
rect 32114 6078 32116 6130
rect 32060 6066 32116 6078
rect 32172 5684 32228 6524
rect 32284 6514 32340 6524
rect 31612 5182 31614 5234
rect 31666 5182 31668 5234
rect 31612 5170 31668 5182
rect 32060 5236 32116 5246
rect 32172 5236 32228 5628
rect 32060 5234 32228 5236
rect 32060 5182 32062 5234
rect 32114 5182 32228 5234
rect 32060 5180 32228 5182
rect 32396 6132 32452 6636
rect 32620 6580 32676 8540
rect 33068 8484 33124 9996
rect 33292 9940 33348 10220
rect 33292 9874 33348 9884
rect 33404 10052 33460 10062
rect 33180 9828 33236 9838
rect 33180 9734 33236 9772
rect 33404 9826 33460 9996
rect 33404 9774 33406 9826
rect 33458 9774 33460 9826
rect 33404 9762 33460 9774
rect 33740 9940 33796 9950
rect 33740 9826 33796 9884
rect 33740 9774 33742 9826
rect 33794 9774 33796 9826
rect 33740 9762 33796 9774
rect 33292 9716 33348 9726
rect 33292 9380 33348 9660
rect 33292 9266 33348 9324
rect 33292 9214 33294 9266
rect 33346 9214 33348 9266
rect 33292 9202 33348 9214
rect 33404 9602 33460 9614
rect 33404 9550 33406 9602
rect 33458 9550 33460 9602
rect 33404 9156 33460 9550
rect 33852 9268 33908 12124
rect 33964 11620 34020 11630
rect 33964 11506 34020 11564
rect 33964 11454 33966 11506
rect 34018 11454 34020 11506
rect 33964 11442 34020 11454
rect 34076 9828 34132 12236
rect 34076 9714 34132 9772
rect 34076 9662 34078 9714
rect 34130 9662 34132 9714
rect 34076 9650 34132 9662
rect 33852 9174 33908 9212
rect 33516 9156 33572 9166
rect 33404 9154 33572 9156
rect 33404 9102 33518 9154
rect 33570 9102 33572 9154
rect 33404 9100 33572 9102
rect 33068 8428 33460 8484
rect 33404 7476 33460 8428
rect 33516 8372 33572 9100
rect 33628 9156 33684 9166
rect 33628 9154 33796 9156
rect 33628 9102 33630 9154
rect 33682 9102 33796 9154
rect 33628 9100 33796 9102
rect 33628 9090 33684 9100
rect 33628 8372 33684 8382
rect 33516 8370 33684 8372
rect 33516 8318 33630 8370
rect 33682 8318 33684 8370
rect 33516 8316 33684 8318
rect 33628 8306 33684 8316
rect 33740 8260 33796 9100
rect 34188 8484 34244 13244
rect 34524 13186 34580 13356
rect 34524 13134 34526 13186
rect 34578 13134 34580 13186
rect 34524 13122 34580 13134
rect 34636 13076 34692 13086
rect 34636 12982 34692 13020
rect 34524 12404 34580 12414
rect 34524 12310 34580 12348
rect 34300 12178 34356 12190
rect 34300 12126 34302 12178
rect 34354 12126 34356 12178
rect 34300 12068 34356 12126
rect 34300 12002 34356 12012
rect 34636 12180 34692 12190
rect 34748 12180 34804 13356
rect 34972 13188 35028 13582
rect 34972 13122 35028 13132
rect 35084 13746 35140 13758
rect 35084 13694 35086 13746
rect 35138 13694 35140 13746
rect 35084 13076 35140 13694
rect 35308 13524 35364 13806
rect 35308 13458 35364 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13010 35140 13020
rect 34860 12964 34916 12974
rect 34860 12870 34916 12908
rect 35196 12962 35252 12974
rect 35532 12964 35588 14028
rect 35868 13972 35924 13982
rect 35756 13634 35812 13646
rect 35756 13582 35758 13634
rect 35810 13582 35812 13634
rect 35756 13524 35812 13582
rect 35756 13458 35812 13468
rect 35868 13300 35924 13916
rect 35756 13244 35924 13300
rect 35196 12910 35198 12962
rect 35250 12910 35252 12962
rect 34972 12850 35028 12862
rect 34972 12798 34974 12850
rect 35026 12798 35028 12850
rect 34860 12292 34916 12302
rect 34972 12292 35028 12798
rect 35196 12404 35252 12910
rect 35196 12338 35252 12348
rect 35308 12908 35588 12964
rect 35644 13188 35700 13198
rect 35644 12962 35700 13132
rect 35644 12910 35646 12962
rect 35698 12910 35700 12962
rect 34860 12290 35028 12292
rect 34860 12238 34862 12290
rect 34914 12238 35028 12290
rect 34860 12236 35028 12238
rect 34860 12226 34916 12236
rect 34636 12178 34804 12180
rect 34636 12126 34638 12178
rect 34690 12126 34804 12178
rect 34636 12124 34804 12126
rect 35308 12180 35364 12908
rect 35644 12898 35700 12910
rect 35532 12738 35588 12750
rect 35532 12686 35534 12738
rect 35586 12686 35588 12738
rect 35532 12516 35588 12686
rect 35532 12450 35588 12460
rect 35308 12178 35588 12180
rect 35308 12126 35310 12178
rect 35362 12126 35588 12178
rect 35308 12124 35588 12126
rect 34636 11956 34692 12124
rect 35308 12114 35364 12124
rect 34636 11890 34692 11900
rect 35084 12068 35140 12078
rect 35084 11506 35140 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 11454 35086 11506
rect 35138 11454 35140 11506
rect 35084 11442 35140 11454
rect 35532 11508 35588 12124
rect 35532 11442 35588 11452
rect 35532 11284 35588 11294
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35420 9940 35476 9950
rect 35532 9940 35588 11228
rect 35420 9938 35588 9940
rect 35420 9886 35422 9938
rect 35474 9886 35588 9938
rect 35420 9884 35588 9886
rect 35420 9874 35476 9884
rect 34524 9828 34580 9838
rect 34412 9714 34468 9726
rect 34412 9662 34414 9714
rect 34466 9662 34468 9714
rect 34412 9156 34468 9662
rect 34412 9090 34468 9100
rect 34188 8418 34244 8428
rect 33964 8260 34020 8270
rect 33740 8258 34020 8260
rect 33740 8206 33966 8258
rect 34018 8206 34020 8258
rect 33740 8204 34020 8206
rect 33740 8034 33796 8046
rect 33740 7982 33742 8034
rect 33794 7982 33796 8034
rect 33516 7476 33572 7486
rect 33404 7474 33572 7476
rect 33404 7422 33518 7474
rect 33570 7422 33572 7474
rect 33404 7420 33572 7422
rect 33516 7410 33572 7420
rect 33628 7476 33684 7486
rect 33740 7476 33796 7982
rect 33964 8036 34020 8204
rect 33964 7970 34020 7980
rect 33628 7474 33796 7476
rect 33628 7422 33630 7474
rect 33682 7422 33796 7474
rect 33628 7420 33796 7422
rect 33852 7588 33908 7598
rect 33628 7410 33684 7420
rect 33852 7364 33908 7532
rect 34188 7476 34244 7486
rect 34188 7382 34244 7420
rect 34300 7474 34356 7486
rect 34300 7422 34302 7474
rect 34354 7422 34356 7474
rect 32620 6514 32676 6524
rect 33740 7308 33908 7364
rect 33628 6356 33684 6366
rect 33740 6356 33796 7308
rect 34300 6580 34356 7422
rect 33684 6300 33796 6356
rect 33852 6524 34356 6580
rect 34524 7474 34580 9772
rect 35644 9828 35700 9838
rect 35644 9734 35700 9772
rect 35756 9604 35812 13244
rect 35868 13076 35924 13086
rect 35868 12962 35924 13020
rect 37100 13076 37156 14588
rect 37548 14532 37604 15708
rect 37772 15202 37828 15932
rect 37884 15876 37940 15886
rect 37884 15782 37940 15820
rect 38108 15538 38164 16380
rect 38332 16324 38388 16334
rect 38220 16268 38332 16324
rect 38220 16210 38276 16268
rect 38332 16258 38388 16268
rect 38220 16158 38222 16210
rect 38274 16158 38276 16210
rect 38220 16146 38276 16158
rect 38108 15486 38110 15538
rect 38162 15486 38164 15538
rect 38108 15474 38164 15486
rect 38556 15876 38612 15886
rect 38444 15316 38500 15326
rect 38444 15222 38500 15260
rect 37772 15150 37774 15202
rect 37826 15150 37828 15202
rect 37548 14530 37716 14532
rect 37548 14478 37550 14530
rect 37602 14478 37716 14530
rect 37548 14476 37716 14478
rect 37548 14466 37604 14476
rect 37212 14306 37268 14318
rect 37212 14254 37214 14306
rect 37266 14254 37268 14306
rect 37212 13524 37268 14254
rect 37212 13458 37268 13468
rect 37548 13634 37604 13646
rect 37548 13582 37550 13634
rect 37602 13582 37604 13634
rect 37548 13524 37604 13582
rect 37548 13458 37604 13468
rect 37660 13522 37716 14476
rect 37660 13470 37662 13522
rect 37714 13470 37716 13522
rect 37660 13458 37716 13470
rect 37100 12982 37156 13020
rect 35868 12910 35870 12962
rect 35922 12910 35924 12962
rect 35868 12628 35924 12910
rect 36316 12964 36372 12974
rect 36316 12870 36372 12908
rect 35868 12562 35924 12572
rect 35980 12516 36036 12526
rect 35980 12290 36036 12460
rect 35980 12238 35982 12290
rect 36034 12238 36036 12290
rect 35980 12226 36036 12238
rect 37660 11956 37716 11966
rect 35308 9548 35812 9604
rect 35868 9826 35924 9838
rect 35868 9774 35870 9826
rect 35922 9774 35924 9826
rect 35084 9044 35140 9054
rect 34524 7422 34526 7474
rect 34578 7422 34580 7474
rect 33628 6290 33684 6300
rect 32396 6130 32788 6132
rect 32396 6078 32398 6130
rect 32450 6078 32788 6130
rect 32396 6076 32788 6078
rect 32060 5124 32116 5180
rect 32060 5058 32116 5068
rect 31500 4452 31556 4462
rect 31388 4450 31556 4452
rect 31388 4398 31502 4450
rect 31554 4398 31556 4450
rect 31388 4396 31556 4398
rect 31500 4386 31556 4396
rect 32284 4340 32340 4350
rect 32396 4340 32452 6076
rect 32732 5124 32788 6076
rect 33852 6018 33908 6524
rect 33852 5966 33854 6018
rect 33906 5966 33908 6018
rect 33852 5954 33908 5966
rect 33740 5684 33796 5694
rect 33516 5682 33796 5684
rect 33516 5630 33742 5682
rect 33794 5630 33796 5682
rect 33516 5628 33796 5630
rect 33516 5234 33572 5628
rect 33740 5618 33796 5628
rect 33516 5182 33518 5234
rect 33570 5182 33572 5234
rect 33516 5170 33572 5182
rect 34524 5236 34580 7422
rect 34972 8036 35028 8046
rect 34972 7252 35028 7980
rect 34972 7186 35028 7196
rect 35084 7474 35140 8988
rect 35308 9042 35364 9548
rect 35532 9156 35588 9166
rect 35532 9062 35588 9100
rect 35308 8990 35310 9042
rect 35362 8990 35364 9042
rect 35308 8978 35364 8990
rect 35868 9044 35924 9774
rect 36092 9828 36148 9838
rect 36092 9734 36148 9772
rect 37100 9828 37156 9838
rect 36540 9716 36596 9726
rect 36540 9622 36596 9660
rect 37100 9156 37156 9772
rect 37660 9826 37716 11900
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37660 9762 37716 9774
rect 37772 9714 37828 15150
rect 38556 15204 38612 15820
rect 38668 15204 38724 15214
rect 38556 15202 38724 15204
rect 38556 15150 38670 15202
rect 38722 15150 38724 15202
rect 38556 15148 38724 15150
rect 38332 14756 38388 14766
rect 38332 14642 38388 14700
rect 38332 14590 38334 14642
rect 38386 14590 38388 14642
rect 38332 14578 38388 14590
rect 37884 14306 37940 14318
rect 37884 14254 37886 14306
rect 37938 14254 37940 14306
rect 37884 13524 37940 14254
rect 37884 13458 37940 13468
rect 38108 13634 38164 13646
rect 38108 13582 38110 13634
rect 38162 13582 38164 13634
rect 38108 13522 38164 13582
rect 38108 13470 38110 13522
rect 38162 13470 38164 13522
rect 38108 13458 38164 13470
rect 38444 13634 38500 13646
rect 38444 13582 38446 13634
rect 38498 13582 38500 13634
rect 38444 13524 38500 13582
rect 38444 13458 38500 13468
rect 38108 12066 38164 12078
rect 38108 12014 38110 12066
rect 38162 12014 38164 12066
rect 38108 11956 38164 12014
rect 38108 11890 38164 11900
rect 38332 11508 38388 11518
rect 38332 11414 38388 11452
rect 37884 11284 37940 11294
rect 38556 11284 38612 15148
rect 38668 15138 38724 15148
rect 38780 12740 38836 18956
rect 38892 18918 38948 18956
rect 39004 15540 39060 21534
rect 39340 19348 39396 19358
rect 39116 19292 39340 19348
rect 39116 19234 39172 19292
rect 39340 19282 39396 19292
rect 39788 19348 39844 19358
rect 39788 19254 39844 19292
rect 39116 19182 39118 19234
rect 39170 19182 39172 19234
rect 39116 19170 39172 19182
rect 39340 19124 39396 19134
rect 39340 19122 39732 19124
rect 39340 19070 39342 19122
rect 39394 19070 39732 19122
rect 39340 19068 39732 19070
rect 39340 19058 39396 19068
rect 39564 18788 39620 18798
rect 39564 18674 39620 18732
rect 39564 18622 39566 18674
rect 39618 18622 39620 18674
rect 39564 18610 39620 18622
rect 39676 18674 39732 19068
rect 39676 18622 39678 18674
rect 39730 18622 39732 18674
rect 39676 18610 39732 18622
rect 39788 18562 39844 18574
rect 39788 18510 39790 18562
rect 39842 18510 39844 18562
rect 39788 17780 39844 18510
rect 39788 17714 39844 17724
rect 38892 15484 39060 15540
rect 39116 16660 39172 16670
rect 38892 15148 38948 15484
rect 39116 15426 39172 16604
rect 39116 15374 39118 15426
rect 39170 15374 39172 15426
rect 39116 15362 39172 15374
rect 39564 15876 39620 15886
rect 39564 15316 39620 15820
rect 39564 15222 39620 15260
rect 39900 15314 39956 15326
rect 39900 15262 39902 15314
rect 39954 15262 39956 15314
rect 39676 15202 39732 15214
rect 39676 15150 39678 15202
rect 39730 15150 39732 15202
rect 39676 15148 39732 15150
rect 38892 15092 39284 15148
rect 39676 15092 39844 15148
rect 39004 14418 39060 14430
rect 39004 14366 39006 14418
rect 39058 14366 39060 14418
rect 39004 13748 39060 14366
rect 39004 13682 39060 13692
rect 39228 14306 39284 15092
rect 39788 14532 39844 15092
rect 39676 14530 39844 14532
rect 39676 14478 39790 14530
rect 39842 14478 39844 14530
rect 39676 14476 39844 14478
rect 39564 14420 39620 14430
rect 39228 14254 39230 14306
rect 39282 14254 39284 14306
rect 39004 13524 39060 13534
rect 38780 12646 38836 12684
rect 38892 13522 39060 13524
rect 38892 13470 39006 13522
rect 39058 13470 39060 13522
rect 38892 13468 39060 13470
rect 38780 12178 38836 12190
rect 38780 12126 38782 12178
rect 38834 12126 38836 12178
rect 38780 11844 38836 12126
rect 38892 11956 38948 13468
rect 39004 13458 39060 13468
rect 39116 13522 39172 13534
rect 39116 13470 39118 13522
rect 39170 13470 39172 13522
rect 39116 13412 39172 13470
rect 39228 13524 39284 14254
rect 39340 14364 39564 14420
rect 39340 13746 39396 14364
rect 39564 14326 39620 14364
rect 39340 13694 39342 13746
rect 39394 13694 39396 13746
rect 39340 13682 39396 13694
rect 39564 13748 39620 13758
rect 39676 13748 39732 14476
rect 39788 14466 39844 14476
rect 39564 13746 39732 13748
rect 39564 13694 39566 13746
rect 39618 13694 39732 13746
rect 39564 13692 39732 13694
rect 39564 13682 39620 13692
rect 39228 13468 39844 13524
rect 39116 13346 39172 13356
rect 39228 13300 39284 13310
rect 39228 13188 39284 13244
rect 39116 13132 39284 13188
rect 39004 12404 39060 12414
rect 39004 12310 39060 12348
rect 39116 12290 39172 13132
rect 39676 12962 39732 12974
rect 39676 12910 39678 12962
rect 39730 12910 39732 12962
rect 39676 12740 39732 12910
rect 39676 12674 39732 12684
rect 39676 12516 39732 12526
rect 39340 12404 39396 12414
rect 39396 12348 39620 12404
rect 39340 12338 39396 12348
rect 39116 12238 39118 12290
rect 39170 12238 39172 12290
rect 39116 12226 39172 12238
rect 39228 12178 39284 12190
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 39228 11956 39284 12126
rect 39564 12178 39620 12348
rect 39564 12126 39566 12178
rect 39618 12126 39620 12178
rect 39564 12114 39620 12126
rect 38892 11900 39284 11956
rect 38780 11778 38836 11788
rect 39452 11508 39508 11518
rect 39452 11394 39508 11452
rect 39452 11342 39454 11394
rect 39506 11342 39508 11394
rect 38668 11284 38724 11294
rect 38556 11228 38668 11284
rect 37884 11190 37940 11228
rect 38668 11190 38724 11228
rect 39004 11170 39060 11182
rect 39004 11118 39006 11170
rect 39058 11118 39060 11170
rect 39004 10164 39060 11118
rect 39004 10098 39060 10108
rect 37772 9662 37774 9714
rect 37826 9662 37828 9714
rect 37772 9650 37828 9662
rect 37324 9492 37380 9502
rect 37100 9154 37268 9156
rect 37100 9102 37102 9154
rect 37154 9102 37268 9154
rect 37100 9100 37268 9102
rect 37100 9090 37156 9100
rect 35868 8978 35924 8988
rect 35420 8930 35476 8942
rect 35420 8878 35422 8930
rect 35474 8878 35476 8930
rect 35420 8820 35476 8878
rect 35420 8764 35588 8820
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35308 8484 35364 8494
rect 35532 8484 35588 8764
rect 35308 8482 35924 8484
rect 35308 8430 35310 8482
rect 35362 8430 35924 8482
rect 35308 8428 35924 8430
rect 35308 8418 35364 8428
rect 35532 8258 35588 8270
rect 35532 8206 35534 8258
rect 35586 8206 35588 8258
rect 35532 7700 35588 8206
rect 35868 8258 35924 8428
rect 35868 8206 35870 8258
rect 35922 8206 35924 8258
rect 35868 8194 35924 8206
rect 36316 8260 36372 8270
rect 36316 8146 36372 8204
rect 36316 8094 36318 8146
rect 36370 8094 36372 8146
rect 36316 8082 36372 8094
rect 36764 8148 36820 8158
rect 35532 7634 35588 7644
rect 35980 8034 36036 8046
rect 35980 7982 35982 8034
rect 36034 7982 36036 8034
rect 35644 7588 35700 7598
rect 35644 7494 35700 7532
rect 35084 7422 35086 7474
rect 35138 7422 35140 7474
rect 34524 5170 34580 5180
rect 32732 5122 33236 5124
rect 32732 5070 32734 5122
rect 32786 5070 33236 5122
rect 32732 5068 33236 5070
rect 32732 5058 32788 5068
rect 33180 4562 33236 5068
rect 33180 4510 33182 4562
rect 33234 4510 33236 4562
rect 33180 4498 33236 4510
rect 32284 4338 32452 4340
rect 32284 4286 32286 4338
rect 32338 4286 32452 4338
rect 32284 4284 32452 4286
rect 32284 4274 32340 4284
rect 29372 4174 29374 4226
rect 29426 4174 29428 4226
rect 29372 4162 29428 4174
rect 34300 4228 34356 4238
rect 35084 4228 35140 7422
rect 35308 7474 35364 7486
rect 35308 7422 35310 7474
rect 35362 7422 35364 7474
rect 35308 7252 35364 7422
rect 35420 7476 35476 7486
rect 35980 7476 36036 7982
rect 36092 8034 36148 8046
rect 36092 7982 36094 8034
rect 36146 7982 36148 8034
rect 36092 7700 36148 7982
rect 36764 7700 36820 8092
rect 36092 7634 36148 7644
rect 36540 7698 36820 7700
rect 36540 7646 36766 7698
rect 36818 7646 36820 7698
rect 36540 7644 36820 7646
rect 36428 7588 36484 7598
rect 36428 7494 36484 7532
rect 36092 7476 36148 7486
rect 35980 7474 36148 7476
rect 35980 7422 36094 7474
rect 36146 7422 36148 7474
rect 35980 7420 36148 7422
rect 35420 7382 35476 7420
rect 36092 7410 36148 7420
rect 36540 7364 36596 7644
rect 36764 7634 36820 7644
rect 36204 7308 36596 7364
rect 35980 7252 36036 7262
rect 35308 7196 35588 7252
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35420 6020 35476 6030
rect 35532 6020 35588 7196
rect 35980 7158 36036 7196
rect 36204 6802 36260 7308
rect 37212 7028 37268 9100
rect 37324 9154 37380 9436
rect 37324 9102 37326 9154
rect 37378 9102 37380 9154
rect 37324 9090 37380 9102
rect 37660 9156 37716 9166
rect 37660 9062 37716 9100
rect 39228 9156 39284 9166
rect 39228 9062 39284 9100
rect 37548 8930 37604 8942
rect 37548 8878 37550 8930
rect 37602 8878 37604 8930
rect 37436 7700 37492 7710
rect 37436 7252 37492 7644
rect 37548 7476 37604 8878
rect 39004 8036 39060 8046
rect 38444 7700 38500 7710
rect 37884 7698 38500 7700
rect 37884 7646 38446 7698
rect 38498 7646 38500 7698
rect 37884 7644 38500 7646
rect 37884 7476 37940 7644
rect 38444 7634 38500 7644
rect 38892 7700 38948 7710
rect 39004 7700 39060 7980
rect 38948 7644 39060 7700
rect 39340 8034 39396 8046
rect 39340 7982 39342 8034
rect 39394 7982 39396 8034
rect 38892 7634 38948 7644
rect 37548 7474 37940 7476
rect 37548 7422 37886 7474
rect 37938 7422 37940 7474
rect 37548 7420 37940 7422
rect 37884 7410 37940 7420
rect 38108 7476 38164 7486
rect 38108 7382 38164 7420
rect 38668 7476 38724 7486
rect 39116 7476 39172 7486
rect 38724 7420 39060 7476
rect 38668 7382 38724 7420
rect 38220 7364 38276 7374
rect 37548 7252 37604 7262
rect 37436 7250 37604 7252
rect 37436 7198 37550 7250
rect 37602 7198 37604 7250
rect 37436 7196 37604 7198
rect 37548 7140 37604 7196
rect 37548 7084 38052 7140
rect 37996 7028 38052 7084
rect 36204 6750 36206 6802
rect 36258 6750 36260 6802
rect 36204 6738 36260 6750
rect 36988 6972 37940 7028
rect 35420 6018 35588 6020
rect 35420 5966 35422 6018
rect 35474 5966 35588 6018
rect 35420 5964 35588 5966
rect 35420 5954 35476 5964
rect 35532 5684 35588 5694
rect 35532 5682 36484 5684
rect 35532 5630 35534 5682
rect 35586 5630 36484 5682
rect 35532 5628 36484 5630
rect 35532 5618 35588 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 5236 35700 5246
rect 35644 5142 35700 5180
rect 36428 4450 36484 5628
rect 36988 5234 37044 6972
rect 37884 6690 37940 6972
rect 37996 6962 38052 6972
rect 37884 6638 37886 6690
rect 37938 6638 37940 6690
rect 37884 6626 37940 6638
rect 38220 6690 38276 7308
rect 38556 7362 38612 7374
rect 38556 7310 38558 7362
rect 38610 7310 38612 7362
rect 38556 7252 38612 7310
rect 38556 7196 38948 7252
rect 38780 7028 38836 7038
rect 38780 6914 38836 6972
rect 38780 6862 38782 6914
rect 38834 6862 38836 6914
rect 38780 6850 38836 6862
rect 38892 6914 38948 7196
rect 38892 6862 38894 6914
rect 38946 6862 38948 6914
rect 38892 6850 38948 6862
rect 39004 6916 39060 7420
rect 39116 7382 39172 7420
rect 39004 6850 39060 6860
rect 39340 7364 39396 7982
rect 38220 6638 38222 6690
rect 38274 6638 38276 6690
rect 38220 6626 38276 6638
rect 39340 6692 39396 7308
rect 39340 6626 39396 6636
rect 38556 6580 38612 6590
rect 38556 6486 38612 6524
rect 38108 6466 38164 6478
rect 38108 6414 38110 6466
rect 38162 6414 38164 6466
rect 36988 5182 36990 5234
rect 37042 5182 37044 5234
rect 36988 5170 37044 5182
rect 37660 5348 37716 5358
rect 37660 4564 37716 5292
rect 36428 4398 36430 4450
rect 36482 4398 36484 4450
rect 36428 4386 36484 4398
rect 37212 4562 37716 4564
rect 37212 4510 37662 4562
rect 37714 4510 37716 4562
rect 37212 4508 37716 4510
rect 37212 4338 37268 4508
rect 37660 4498 37716 4508
rect 38108 4450 38164 6414
rect 39452 5348 39508 11342
rect 39676 10948 39732 12460
rect 39788 12180 39844 13468
rect 39900 13300 39956 15262
rect 40012 13970 40068 23660
rect 40348 21812 40404 25676
rect 40348 21718 40404 21756
rect 40348 20132 40404 20142
rect 40348 19236 40404 20076
rect 40348 19170 40404 19180
rect 40236 18900 40292 18910
rect 40236 18450 40292 18844
rect 40236 18398 40238 18450
rect 40290 18398 40292 18450
rect 40236 18340 40292 18398
rect 40236 18274 40292 18284
rect 40460 14644 40516 26852
rect 41916 26516 41972 26852
rect 41916 26422 41972 26460
rect 41468 26404 41524 26414
rect 41468 26310 41524 26348
rect 40684 26292 40740 26302
rect 40684 25732 40740 26236
rect 41132 26292 41188 26302
rect 41132 26198 41188 26236
rect 41020 26068 41076 26078
rect 41020 25974 41076 26012
rect 41356 26066 41412 26078
rect 41356 26014 41358 26066
rect 41410 26014 41412 26066
rect 40684 25730 40964 25732
rect 40684 25678 40686 25730
rect 40738 25678 40964 25730
rect 40684 25676 40964 25678
rect 40684 25666 40740 25676
rect 40684 25508 40740 25518
rect 40572 25396 40628 25406
rect 40572 25302 40628 25340
rect 40684 25394 40740 25452
rect 40684 25342 40686 25394
rect 40738 25342 40740 25394
rect 40684 25330 40740 25342
rect 40908 24834 40964 25676
rect 41356 25396 41412 26014
rect 41356 25330 41412 25340
rect 41916 25506 41972 25518
rect 41916 25454 41918 25506
rect 41970 25454 41972 25506
rect 41468 25284 41524 25294
rect 41468 25190 41524 25228
rect 41692 25282 41748 25294
rect 41692 25230 41694 25282
rect 41746 25230 41748 25282
rect 40908 24782 40910 24834
rect 40962 24782 40964 24834
rect 40908 24770 40964 24782
rect 41132 24836 41188 24846
rect 41132 24742 41188 24780
rect 41020 24612 41076 24622
rect 40460 14578 40516 14588
rect 40572 24610 41076 24612
rect 40572 24558 41022 24610
rect 41074 24558 41076 24610
rect 40572 24556 41076 24558
rect 40012 13918 40014 13970
rect 40066 13918 40068 13970
rect 40012 13412 40068 13918
rect 40572 13524 40628 24556
rect 41020 24546 41076 24556
rect 41244 23492 41300 23502
rect 41020 23156 41076 23166
rect 41244 23156 41300 23436
rect 41076 23100 41300 23156
rect 41020 23062 41076 23100
rect 40684 22484 40740 22494
rect 40684 22390 40740 22428
rect 41244 22370 41300 23100
rect 41244 22318 41246 22370
rect 41298 22318 41300 22370
rect 41244 22306 41300 22318
rect 41468 22260 41524 22270
rect 41468 21810 41524 22204
rect 41468 21758 41470 21810
rect 41522 21758 41524 21810
rect 41468 21746 41524 21758
rect 41580 21812 41636 21822
rect 41580 21698 41636 21756
rect 41580 21646 41582 21698
rect 41634 21646 41636 21698
rect 41580 21634 41636 21646
rect 41132 21588 41188 21598
rect 40908 21586 41188 21588
rect 40908 21534 41134 21586
rect 41186 21534 41188 21586
rect 40908 21532 41188 21534
rect 40908 20018 40964 21532
rect 41132 21522 41188 21532
rect 41580 20578 41636 20590
rect 41580 20526 41582 20578
rect 41634 20526 41636 20578
rect 41244 20132 41300 20142
rect 41244 20038 41300 20076
rect 40908 19966 40910 20018
rect 40962 19966 40964 20018
rect 40908 19572 40964 19966
rect 41468 20020 41524 20030
rect 41580 20020 41636 20526
rect 41692 20580 41748 25230
rect 41916 25284 41972 25454
rect 41916 25218 41972 25228
rect 42140 25060 42196 25070
rect 42140 24834 42196 25004
rect 42140 24782 42142 24834
rect 42194 24782 42196 24834
rect 42140 24770 42196 24782
rect 41804 24724 41860 24734
rect 41804 24630 41860 24668
rect 42140 23380 42196 23390
rect 41804 23378 42196 23380
rect 41804 23326 42142 23378
rect 42194 23326 42196 23378
rect 41804 23324 42196 23326
rect 42364 23380 42420 29932
rect 42924 29652 42980 29662
rect 43484 29652 43540 30716
rect 42924 29650 43540 29652
rect 42924 29598 42926 29650
rect 42978 29598 43486 29650
rect 43538 29598 43540 29650
rect 42924 29596 43540 29598
rect 42924 29586 42980 29596
rect 43484 29586 43540 29596
rect 44044 29314 44100 29326
rect 44044 29262 44046 29314
rect 44098 29262 44100 29314
rect 42812 29204 42868 29214
rect 42812 29110 42868 29148
rect 43148 29204 43204 29214
rect 43148 29202 43428 29204
rect 43148 29150 43150 29202
rect 43202 29150 43428 29202
rect 43148 29148 43428 29150
rect 43148 29138 43204 29148
rect 43372 28756 43428 29148
rect 43820 29202 43876 29214
rect 43820 29150 43822 29202
rect 43874 29150 43876 29202
rect 43484 28756 43540 28766
rect 43372 28754 43540 28756
rect 43372 28702 43486 28754
rect 43538 28702 43540 28754
rect 43372 28700 43540 28702
rect 43484 28690 43540 28700
rect 42700 28644 42756 28654
rect 43036 28644 43092 28654
rect 42700 28642 43092 28644
rect 42700 28590 42702 28642
rect 42754 28590 43038 28642
rect 43090 28590 43092 28642
rect 42700 28588 43092 28590
rect 42700 28578 42756 28588
rect 42588 27188 42644 27198
rect 42588 26290 42644 27132
rect 42588 26238 42590 26290
rect 42642 26238 42644 26290
rect 42476 25396 42532 25406
rect 42476 25302 42532 25340
rect 42588 25284 42644 26238
rect 42924 25284 42980 25294
rect 42588 25282 42980 25284
rect 42588 25230 42926 25282
rect 42978 25230 42980 25282
rect 42588 25228 42980 25230
rect 42700 24724 42756 24734
rect 42700 24630 42756 24668
rect 42924 23604 42980 25228
rect 43036 25060 43092 28588
rect 43372 28420 43428 28430
rect 43372 28326 43428 28364
rect 43596 28420 43652 28430
rect 43820 28420 43876 29150
rect 44044 28420 44100 29262
rect 43596 28418 43876 28420
rect 43596 28366 43598 28418
rect 43650 28366 43876 28418
rect 43596 28364 43876 28366
rect 43932 28364 44044 28420
rect 43596 27524 43652 28364
rect 43932 27746 43988 28364
rect 44044 28354 44100 28364
rect 44380 28756 44436 28766
rect 44380 28082 44436 28700
rect 44380 28030 44382 28082
rect 44434 28030 44436 28082
rect 44380 28018 44436 28030
rect 43932 27694 43934 27746
rect 43986 27694 43988 27746
rect 43932 27682 43988 27694
rect 43596 27468 44100 27524
rect 43932 26852 43988 26862
rect 43820 26796 43932 26852
rect 43708 26516 43764 26526
rect 43260 26178 43316 26190
rect 43260 26126 43262 26178
rect 43314 26126 43316 26178
rect 43260 25732 43316 26126
rect 43596 25732 43652 25742
rect 43260 25730 43652 25732
rect 43260 25678 43598 25730
rect 43650 25678 43652 25730
rect 43260 25676 43652 25678
rect 43596 25666 43652 25676
rect 43036 24994 43092 25004
rect 43708 25506 43764 26460
rect 43708 25454 43710 25506
rect 43762 25454 43764 25506
rect 43708 25396 43764 25454
rect 43148 24892 43540 24948
rect 43148 24722 43204 24892
rect 43148 24670 43150 24722
rect 43202 24670 43204 24722
rect 43148 24658 43204 24670
rect 43372 24724 43428 24734
rect 42924 23538 42980 23548
rect 43260 23828 43316 23838
rect 42476 23380 42532 23390
rect 43148 23380 43204 23390
rect 42364 23378 43204 23380
rect 42364 23326 42478 23378
rect 42530 23326 43150 23378
rect 43202 23326 43204 23378
rect 42364 23324 43204 23326
rect 41804 21698 41860 23324
rect 42140 23314 42196 23324
rect 42476 23314 42532 23324
rect 43148 23314 43204 23324
rect 42028 23154 42084 23166
rect 42028 23102 42030 23154
rect 42082 23102 42084 23154
rect 42028 22596 42084 23102
rect 42252 23156 42308 23166
rect 42252 23062 42308 23100
rect 42028 22540 42308 22596
rect 42028 22260 42084 22270
rect 42028 22166 42084 22204
rect 41804 21646 41806 21698
rect 41858 21646 41860 21698
rect 41804 21634 41860 21646
rect 41692 20524 41972 20580
rect 41804 20020 41860 20030
rect 41580 20018 41860 20020
rect 41580 19966 41806 20018
rect 41858 19966 41860 20018
rect 41580 19964 41860 19966
rect 41468 19926 41524 19964
rect 41020 19908 41076 19918
rect 41020 19814 41076 19852
rect 40908 18564 40964 19516
rect 41244 18788 41300 18798
rect 41244 18674 41300 18732
rect 41244 18622 41246 18674
rect 41298 18622 41300 18674
rect 41244 18610 41300 18622
rect 40908 18498 40964 18508
rect 41356 18452 41412 18462
rect 41356 18358 41412 18396
rect 41468 18450 41524 18462
rect 41468 18398 41470 18450
rect 41522 18398 41524 18450
rect 41468 17892 41524 18398
rect 41468 17826 41524 17836
rect 40684 17780 40740 17790
rect 40684 15316 40740 17724
rect 41468 17668 41524 17678
rect 41692 17668 41748 19964
rect 41804 19954 41860 19964
rect 41804 19010 41860 19022
rect 41804 18958 41806 19010
rect 41858 18958 41860 19010
rect 41804 18450 41860 18958
rect 41804 18398 41806 18450
rect 41858 18398 41860 18450
rect 41804 18340 41860 18398
rect 41804 18274 41860 18284
rect 41468 17666 41692 17668
rect 41468 17614 41470 17666
rect 41522 17614 41692 17666
rect 41468 17612 41692 17614
rect 41020 16772 41076 16782
rect 41468 16772 41524 17612
rect 41692 17574 41748 17612
rect 41020 16770 41524 16772
rect 41020 16718 41022 16770
rect 41074 16718 41470 16770
rect 41522 16718 41524 16770
rect 41020 16716 41524 16718
rect 41020 16324 41076 16716
rect 40908 15316 40964 15326
rect 40684 15314 40964 15316
rect 40684 15262 40910 15314
rect 40962 15262 40964 15314
rect 40684 15260 40964 15262
rect 40908 15250 40964 15260
rect 41020 15316 41076 16268
rect 41468 16210 41524 16716
rect 41468 16158 41470 16210
rect 41522 16158 41524 16210
rect 41468 16146 41524 16158
rect 40572 13458 40628 13468
rect 40908 14420 40964 14430
rect 40012 13346 40068 13356
rect 39900 13234 39956 13244
rect 39900 12404 39956 12414
rect 39900 12402 40180 12404
rect 39900 12350 39902 12402
rect 39954 12350 40180 12402
rect 39900 12348 40180 12350
rect 39900 12338 39956 12348
rect 39900 12180 39956 12190
rect 39788 12178 39956 12180
rect 39788 12126 39902 12178
rect 39954 12126 39956 12178
rect 39788 12124 39956 12126
rect 39900 12114 39956 12124
rect 40124 11508 40180 12348
rect 40908 12290 40964 14364
rect 40908 12238 40910 12290
rect 40962 12238 40964 12290
rect 40908 12226 40964 12238
rect 41020 13074 41076 15260
rect 41132 15876 41188 15886
rect 41132 15314 41188 15820
rect 41916 15764 41972 20524
rect 42140 20020 42196 20030
rect 42140 19346 42196 19964
rect 42140 19294 42142 19346
rect 42194 19294 42196 19346
rect 42140 19282 42196 19294
rect 42252 19460 42308 22540
rect 42588 19908 42644 19918
rect 42588 19814 42644 19852
rect 42252 19234 42308 19404
rect 42252 19182 42254 19234
rect 42306 19182 42308 19234
rect 42252 19170 42308 19182
rect 42028 19012 42084 19022
rect 42028 18918 42084 18956
rect 42364 18676 42420 18686
rect 42140 18564 42196 18574
rect 42140 18470 42196 18508
rect 42364 18450 42420 18620
rect 43148 18676 43204 18686
rect 42364 18398 42366 18450
rect 42418 18398 42420 18450
rect 42364 18386 42420 18398
rect 42588 18452 42644 18462
rect 42588 18358 42644 18396
rect 43148 18450 43204 18620
rect 43148 18398 43150 18450
rect 43202 18398 43204 18450
rect 43148 18386 43204 18398
rect 42252 18338 42308 18350
rect 42252 18286 42254 18338
rect 42306 18286 42308 18338
rect 42140 17780 42196 17790
rect 42252 17780 42308 18286
rect 42140 17778 42308 17780
rect 42140 17726 42142 17778
rect 42194 17726 42308 17778
rect 42140 17724 42308 17726
rect 43036 18228 43092 18238
rect 42140 17714 42196 17724
rect 41916 15698 41972 15708
rect 41132 15262 41134 15314
rect 41186 15262 41188 15314
rect 41132 15250 41188 15262
rect 41916 15316 41972 15326
rect 41916 15222 41972 15260
rect 42588 15202 42644 15214
rect 42588 15150 42590 15202
rect 42642 15150 42644 15202
rect 42588 15148 42644 15150
rect 43036 15148 43092 18172
rect 41468 15090 41524 15102
rect 41468 15038 41470 15090
rect 41522 15038 41524 15090
rect 41468 14644 41524 15038
rect 41468 14550 41524 14588
rect 41692 15092 41748 15102
rect 41692 14530 41748 15036
rect 42476 15092 42644 15148
rect 42812 15092 42868 15102
rect 41692 14478 41694 14530
rect 41746 14478 41748 14530
rect 41692 14466 41748 14478
rect 41916 14532 41972 14542
rect 41916 14438 41972 14476
rect 41468 14308 41524 14318
rect 41020 13022 41022 13074
rect 41074 13022 41076 13074
rect 40236 12178 40292 12190
rect 40236 12126 40238 12178
rect 40290 12126 40292 12178
rect 40236 12068 40292 12126
rect 40236 12002 40292 12012
rect 40236 11508 40292 11518
rect 40124 11506 40292 11508
rect 40124 11454 40238 11506
rect 40290 11454 40292 11506
rect 40124 11452 40292 11454
rect 40236 11442 40292 11452
rect 41020 11508 41076 13022
rect 41132 13860 41188 13870
rect 41132 12852 41188 13804
rect 41468 13858 41524 14252
rect 41468 13806 41470 13858
rect 41522 13806 41524 13858
rect 41468 13794 41524 13806
rect 41916 13972 41972 13982
rect 41132 12402 41188 12796
rect 41132 12350 41134 12402
rect 41186 12350 41188 12402
rect 41132 12338 41188 12350
rect 41692 13746 41748 13758
rect 41692 13694 41694 13746
rect 41746 13694 41748 13746
rect 41692 12292 41748 13694
rect 41916 13746 41972 13916
rect 42476 13970 42532 15092
rect 42588 14644 42644 14654
rect 42588 14530 42644 14588
rect 42588 14478 42590 14530
rect 42642 14478 42644 14530
rect 42588 14466 42644 14478
rect 42812 14530 42868 15036
rect 42812 14478 42814 14530
rect 42866 14478 42868 14530
rect 42700 14308 42756 14318
rect 42700 14214 42756 14252
rect 42476 13918 42478 13970
rect 42530 13918 42532 13970
rect 42476 13906 42532 13918
rect 42812 13858 42868 14478
rect 42812 13806 42814 13858
rect 42866 13806 42868 13858
rect 42812 13794 42868 13806
rect 42924 15092 43092 15148
rect 41916 13694 41918 13746
rect 41970 13694 41972 13746
rect 41916 13682 41972 13694
rect 42364 13748 42420 13758
rect 42700 13748 42756 13758
rect 42364 13746 42756 13748
rect 42364 13694 42366 13746
rect 42418 13694 42702 13746
rect 42754 13694 42756 13746
rect 42364 13692 42756 13694
rect 42364 13682 42420 13692
rect 42700 13682 42756 13692
rect 42140 13636 42196 13646
rect 42028 12852 42084 12862
rect 42028 12758 42084 12796
rect 42140 12516 42196 13580
rect 42476 13524 42532 13534
rect 42364 13300 42420 13310
rect 42140 12450 42196 12460
rect 42252 13244 42364 13300
rect 41244 12236 41748 12292
rect 41244 12066 41300 12236
rect 41244 12014 41246 12066
rect 41298 12014 41300 12066
rect 41244 12002 41300 12014
rect 41692 12066 41748 12078
rect 41692 12014 41694 12066
rect 41746 12014 41748 12066
rect 41692 11844 41748 12014
rect 41692 11778 41748 11788
rect 42140 12068 42196 12078
rect 41020 11442 41076 11452
rect 39676 10882 39732 10892
rect 41804 10610 41860 10622
rect 41804 10558 41806 10610
rect 41858 10558 41860 10610
rect 40236 10164 40292 10174
rect 39564 9714 39620 9726
rect 39564 9662 39566 9714
rect 39618 9662 39620 9714
rect 39564 9154 39620 9662
rect 40236 9266 40292 10108
rect 41804 10164 41860 10558
rect 42140 10388 42196 12012
rect 42252 11508 42308 13244
rect 42364 13234 42420 13244
rect 42364 12738 42420 12750
rect 42364 12686 42366 12738
rect 42418 12686 42420 12738
rect 42364 12404 42420 12686
rect 42364 12338 42420 12348
rect 42364 11508 42420 11518
rect 42252 11506 42420 11508
rect 42252 11454 42366 11506
rect 42418 11454 42420 11506
rect 42252 11452 42420 11454
rect 42364 11442 42420 11452
rect 42252 11060 42308 11070
rect 42252 10500 42308 11004
rect 42252 10406 42308 10444
rect 42140 10322 42196 10332
rect 41804 10098 41860 10108
rect 42252 9940 42308 9950
rect 41468 9826 41524 9838
rect 41468 9774 41470 9826
rect 41522 9774 41524 9826
rect 40348 9716 40404 9726
rect 40348 9622 40404 9660
rect 40236 9214 40238 9266
rect 40290 9214 40292 9266
rect 40236 9202 40292 9214
rect 39564 9102 39566 9154
rect 39618 9102 39620 9154
rect 39564 7812 39620 9102
rect 39788 9156 39844 9166
rect 39564 7746 39620 7756
rect 39676 8036 39732 8046
rect 39676 7252 39732 7980
rect 39788 7586 39844 9100
rect 39788 7534 39790 7586
rect 39842 7534 39844 7586
rect 39788 7522 39844 7534
rect 39900 9154 39956 9166
rect 39900 9102 39902 9154
rect 39954 9102 39956 9154
rect 39900 7476 39956 9102
rect 41468 7924 41524 9774
rect 42252 9380 42308 9884
rect 42476 9716 42532 13468
rect 42588 12852 42644 12862
rect 42588 12402 42644 12796
rect 42588 12350 42590 12402
rect 42642 12350 42644 12402
rect 42588 12338 42644 12350
rect 42812 12738 42868 12750
rect 42812 12686 42814 12738
rect 42866 12686 42868 12738
rect 42812 12404 42868 12686
rect 42812 12338 42868 12348
rect 42924 11788 42980 15092
rect 43036 14532 43092 14542
rect 43036 14418 43092 14476
rect 43036 14366 43038 14418
rect 43090 14366 43092 14418
rect 43036 14354 43092 14366
rect 43260 13972 43316 23772
rect 43260 13878 43316 13916
rect 43372 12964 43428 24668
rect 43372 12738 43428 12908
rect 43372 12686 43374 12738
rect 43426 12686 43428 12738
rect 43372 11788 43428 12686
rect 43484 24612 43540 24892
rect 43484 12404 43540 24556
rect 43596 24610 43652 24622
rect 43596 24558 43598 24610
rect 43650 24558 43652 24610
rect 43596 24500 43652 24558
rect 43596 23716 43652 24444
rect 43708 23828 43764 25340
rect 43708 23762 43764 23772
rect 43596 23650 43652 23660
rect 43708 23042 43764 23054
rect 43708 22990 43710 23042
rect 43762 22990 43764 23042
rect 43708 22260 43764 22990
rect 43708 22194 43764 22204
rect 43596 18338 43652 18350
rect 43596 18286 43598 18338
rect 43650 18286 43652 18338
rect 43596 18228 43652 18286
rect 43596 18162 43652 18172
rect 43708 14308 43764 14318
rect 43820 14308 43876 26796
rect 43932 26758 43988 26796
rect 44044 26852 44100 27468
rect 44268 26964 44324 27002
rect 44268 26898 44324 26908
rect 44156 26852 44212 26862
rect 44044 26850 44212 26852
rect 44044 26798 44158 26850
rect 44210 26798 44212 26850
rect 44044 26796 44212 26798
rect 43932 25732 43988 25742
rect 43932 25638 43988 25676
rect 44044 25730 44100 26796
rect 44156 26786 44212 26796
rect 44044 25678 44046 25730
rect 44098 25678 44100 25730
rect 44044 25666 44100 25678
rect 44380 24610 44436 24622
rect 44380 24558 44382 24610
rect 44434 24558 44436 24610
rect 44044 23828 44100 23838
rect 44380 23828 44436 24558
rect 44100 23772 44436 23828
rect 44044 23762 44100 23772
rect 44156 23380 44212 23390
rect 44156 23286 44212 23324
rect 44156 23156 44212 23166
rect 44156 22482 44212 23100
rect 44156 22430 44158 22482
rect 44210 22430 44212 22482
rect 44156 21924 44212 22430
rect 44156 21858 44212 21868
rect 43932 18450 43988 18462
rect 43932 18398 43934 18450
rect 43986 18398 43988 18450
rect 43932 18228 43988 18398
rect 44492 18452 44548 32508
rect 44940 32498 44996 32508
rect 45388 31892 45444 31902
rect 45388 31798 45444 31836
rect 45164 31780 45220 31790
rect 45164 30882 45220 31724
rect 45164 30830 45166 30882
rect 45218 30830 45220 30882
rect 45164 30818 45220 30830
rect 45612 30882 45668 30894
rect 45612 30830 45614 30882
rect 45666 30830 45668 30882
rect 45276 30212 45332 30222
rect 45276 28756 45332 30156
rect 45612 30212 45668 30830
rect 45612 30146 45668 30156
rect 45332 28700 45668 28756
rect 45276 28662 45332 28700
rect 45612 28642 45668 28700
rect 45612 28590 45614 28642
rect 45666 28590 45668 28642
rect 45612 28578 45668 28590
rect 45052 27074 45108 27086
rect 45052 27022 45054 27074
rect 45106 27022 45108 27074
rect 44828 26962 44884 26974
rect 44828 26910 44830 26962
rect 44882 26910 44884 26962
rect 44828 26852 44884 26910
rect 44828 26786 44884 26796
rect 44940 26850 44996 26862
rect 44940 26798 44942 26850
rect 44994 26798 44996 26850
rect 44940 25732 44996 26798
rect 44940 25666 44996 25676
rect 45052 25508 45108 27022
rect 45164 26964 45220 26974
rect 45164 25618 45220 26908
rect 45388 26962 45444 26974
rect 45388 26910 45390 26962
rect 45442 26910 45444 26962
rect 45388 26180 45444 26910
rect 45164 25566 45166 25618
rect 45218 25566 45220 25618
rect 45164 25554 45220 25566
rect 45276 26178 45444 26180
rect 45276 26126 45390 26178
rect 45442 26126 45444 26178
rect 45276 26124 45444 26126
rect 45052 25414 45108 25452
rect 44828 25394 44884 25406
rect 44828 25342 44830 25394
rect 44882 25342 44884 25394
rect 44828 25284 44884 25342
rect 45276 25394 45332 26124
rect 45388 26114 45444 26124
rect 45276 25342 45278 25394
rect 45330 25342 45332 25394
rect 45276 25330 45332 25342
rect 45724 25506 45780 25518
rect 45724 25454 45726 25506
rect 45778 25454 45780 25506
rect 44828 25218 44884 25228
rect 44828 24612 44884 24622
rect 44828 24518 44884 24556
rect 45276 24612 45332 24622
rect 45724 24612 45780 25454
rect 45836 25284 45892 36988
rect 46060 35026 46116 35038
rect 46060 34974 46062 35026
rect 46114 34974 46116 35026
rect 45948 34132 46004 34142
rect 46060 34132 46116 34974
rect 45948 34130 46116 34132
rect 45948 34078 45950 34130
rect 46002 34078 46116 34130
rect 45948 34076 46116 34078
rect 45948 33572 46004 34076
rect 45948 33506 46004 33516
rect 45948 25508 46004 25518
rect 45948 25414 46004 25452
rect 45836 24946 45892 25228
rect 45836 24894 45838 24946
rect 45890 24894 45892 24946
rect 45836 24882 45892 24894
rect 46172 24946 46228 37212
rect 47740 35252 47796 35262
rect 47292 34356 47348 34366
rect 47180 34242 47236 34254
rect 47180 34190 47182 34242
rect 47234 34190 47236 34242
rect 46620 34020 46676 34030
rect 46956 34020 47012 34030
rect 46620 34018 47012 34020
rect 46620 33966 46622 34018
rect 46674 33966 46958 34018
rect 47010 33966 47012 34018
rect 46620 33964 47012 33966
rect 46620 33954 46676 33964
rect 46956 33954 47012 33964
rect 47180 33796 47236 34190
rect 47292 34018 47348 34300
rect 47740 34020 47796 35196
rect 47292 33966 47294 34018
rect 47346 33966 47348 34018
rect 47292 33954 47348 33966
rect 47628 34018 47796 34020
rect 47628 33966 47742 34018
rect 47794 33966 47796 34018
rect 47628 33964 47796 33966
rect 47628 33796 47684 33964
rect 47740 33954 47796 33964
rect 47180 33740 47684 33796
rect 46732 32564 46788 32574
rect 46732 32470 46788 32508
rect 47404 32564 47460 32574
rect 47404 32470 47460 32508
rect 46508 32450 46564 32462
rect 46508 32398 46510 32450
rect 46562 32398 46564 32450
rect 46508 30434 46564 32398
rect 47516 31668 47572 31678
rect 47516 31574 47572 31612
rect 46508 30382 46510 30434
rect 46562 30382 46564 30434
rect 46508 30370 46564 30382
rect 46956 30324 47012 30334
rect 46620 30268 46956 30324
rect 46620 30210 46676 30268
rect 46956 30230 47012 30268
rect 46620 30158 46622 30210
rect 46674 30158 46676 30210
rect 46620 30146 46676 30158
rect 46508 29986 46564 29998
rect 46508 29934 46510 29986
rect 46562 29934 46564 29986
rect 46508 29316 46564 29934
rect 46508 29250 46564 29260
rect 46396 28530 46452 28542
rect 46396 28478 46398 28530
rect 46450 28478 46452 28530
rect 46396 26404 46452 28478
rect 46396 26338 46452 26348
rect 47628 26292 47684 33740
rect 47852 26516 47908 46396
rect 47964 28980 48020 48076
rect 48860 48132 48916 48142
rect 48860 48038 48916 48076
rect 48524 47234 48580 47246
rect 48524 47182 48526 47234
rect 48578 47182 48580 47234
rect 48076 46674 48132 46686
rect 48076 46622 48078 46674
rect 48130 46622 48132 46674
rect 48076 45668 48132 46622
rect 48412 45892 48468 45902
rect 48412 45798 48468 45836
rect 48132 45612 48356 45668
rect 48076 45574 48132 45612
rect 48300 45332 48356 45612
rect 48524 45332 48580 47182
rect 48748 46788 48804 46798
rect 48748 46694 48804 46732
rect 48748 45332 48804 45342
rect 48300 45330 48804 45332
rect 48300 45278 48302 45330
rect 48354 45278 48750 45330
rect 48802 45278 48804 45330
rect 48300 45276 48804 45278
rect 48300 45266 48356 45276
rect 48748 45266 48804 45276
rect 48972 43708 49028 49868
rect 49868 49700 49924 49710
rect 49644 49698 49924 49700
rect 49644 49646 49870 49698
rect 49922 49646 49924 49698
rect 49644 49644 49924 49646
rect 49644 49026 49700 49644
rect 49644 48974 49646 49026
rect 49698 48974 49700 49026
rect 49644 48962 49700 48974
rect 49196 48356 49252 48366
rect 49084 48244 49140 48254
rect 49084 47684 49140 48188
rect 49196 48242 49252 48300
rect 49196 48190 49198 48242
rect 49250 48190 49252 48242
rect 49196 48132 49252 48190
rect 49196 48066 49252 48076
rect 49644 48244 49700 48254
rect 49644 48130 49700 48188
rect 49644 48078 49646 48130
rect 49698 48078 49700 48130
rect 49644 48066 49700 48078
rect 49756 47908 49812 47918
rect 49084 47628 49252 47684
rect 49084 45220 49140 45230
rect 49084 45126 49140 45164
rect 49196 43708 49252 47628
rect 49756 47570 49812 47852
rect 49756 47518 49758 47570
rect 49810 47518 49812 47570
rect 49756 47506 49812 47518
rect 49868 47460 49924 49644
rect 50428 49698 50484 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50876 50034 50932 50316
rect 50876 49982 50878 50034
rect 50930 49982 50932 50034
rect 50876 49970 50932 49982
rect 50428 49646 50430 49698
rect 50482 49646 50484 49698
rect 49308 46676 49364 46686
rect 49756 46676 49812 46686
rect 49364 46620 49588 46676
rect 49308 46582 49364 46620
rect 48748 43652 49028 43708
rect 49084 43652 49252 43708
rect 49308 45890 49364 45902
rect 49308 45838 49310 45890
rect 49362 45838 49364 45890
rect 49308 45780 49364 45838
rect 49308 43708 49364 45724
rect 49532 45892 49588 46620
rect 49756 46582 49812 46620
rect 49532 45778 49588 45836
rect 49532 45726 49534 45778
rect 49586 45726 49588 45778
rect 49532 45714 49588 45726
rect 49868 45108 49924 47404
rect 49980 49028 50036 49038
rect 49980 47684 50036 48972
rect 50092 48244 50148 48254
rect 50428 48244 50484 49646
rect 50764 49924 50820 49934
rect 50764 49138 50820 49868
rect 50764 49086 50766 49138
rect 50818 49086 50820 49138
rect 50764 49074 50820 49086
rect 50876 49364 50932 49374
rect 50652 49028 50708 49038
rect 50652 48934 50708 48972
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50092 48242 50484 48244
rect 50092 48190 50094 48242
rect 50146 48190 50484 48242
rect 50092 48188 50484 48190
rect 50092 47908 50148 48188
rect 50876 48130 50932 49308
rect 50988 48802 51044 51884
rect 51100 51156 51156 51166
rect 51100 50034 51156 51100
rect 51212 50708 51268 52222
rect 51772 52274 51828 53004
rect 51772 52222 51774 52274
rect 51826 52222 51828 52274
rect 51772 52210 51828 52222
rect 51884 51602 51940 53676
rect 52780 53508 52836 53518
rect 52780 53414 52836 53452
rect 51884 51550 51886 51602
rect 51938 51550 51940 51602
rect 51884 51538 51940 51550
rect 52780 51604 52836 51614
rect 52892 51604 52948 53788
rect 53004 53750 53060 53788
rect 53676 53508 53732 53518
rect 53676 52834 53732 53452
rect 53788 52948 53844 55020
rect 53900 55524 53956 56252
rect 54236 56242 54292 56252
rect 55244 56978 55412 56980
rect 55244 56926 55358 56978
rect 55410 56926 55412 56978
rect 55244 56924 55412 56926
rect 54908 56084 54964 56094
rect 53900 53842 53956 55468
rect 54796 56082 54964 56084
rect 54796 56030 54910 56082
rect 54962 56030 54964 56082
rect 54796 56028 54964 56030
rect 54572 54292 54628 54302
rect 53900 53790 53902 53842
rect 53954 53790 53956 53842
rect 53900 53778 53956 53790
rect 54460 54290 54628 54292
rect 54460 54238 54574 54290
rect 54626 54238 54628 54290
rect 54460 54236 54628 54238
rect 54236 53618 54292 53630
rect 54236 53566 54238 53618
rect 54290 53566 54292 53618
rect 54124 52948 54180 52958
rect 53788 52946 54180 52948
rect 53788 52894 54126 52946
rect 54178 52894 54180 52946
rect 53788 52892 54180 52894
rect 54124 52882 54180 52892
rect 53676 52782 53678 52834
rect 53730 52782 53732 52834
rect 53340 52276 53396 52286
rect 52780 51602 52948 51604
rect 52780 51550 52782 51602
rect 52834 51550 52948 51602
rect 52780 51548 52948 51550
rect 53228 52164 53284 52174
rect 52780 51538 52836 51548
rect 53228 51490 53284 52108
rect 53228 51438 53230 51490
rect 53282 51438 53284 51490
rect 53228 51426 53284 51438
rect 52108 51380 52164 51390
rect 52444 51380 52500 51390
rect 52108 51378 52276 51380
rect 52108 51326 52110 51378
rect 52162 51326 52276 51378
rect 52108 51324 52276 51326
rect 52108 51314 52164 51324
rect 51772 51156 51828 51166
rect 51772 51062 51828 51100
rect 52220 51156 52276 51324
rect 52444 51286 52500 51324
rect 53116 51156 53172 51166
rect 52220 51154 53172 51156
rect 52220 51102 53118 51154
rect 53170 51102 53172 51154
rect 52220 51100 53172 51102
rect 51212 50642 51268 50652
rect 51100 49982 51102 50034
rect 51154 49982 51156 50034
rect 51100 49970 51156 49982
rect 52220 49922 52276 51100
rect 53116 51090 53172 51100
rect 53228 50820 53284 50830
rect 52220 49870 52222 49922
rect 52274 49870 52276 49922
rect 52220 49858 52276 49870
rect 52668 49924 52724 49934
rect 51996 49810 52052 49822
rect 51996 49758 51998 49810
rect 52050 49758 52052 49810
rect 51660 49700 51716 49710
rect 51996 49700 52052 49758
rect 52668 49810 52724 49868
rect 52668 49758 52670 49810
rect 52722 49758 52724 49810
rect 52668 49746 52724 49758
rect 51660 49698 52052 49700
rect 51660 49646 51662 49698
rect 51714 49646 52052 49698
rect 51660 49644 52052 49646
rect 52444 49698 52500 49710
rect 52444 49646 52446 49698
rect 52498 49646 52500 49698
rect 51660 49364 51716 49644
rect 52444 49364 52500 49646
rect 52444 49308 53060 49364
rect 51660 49298 51716 49308
rect 53004 49250 53060 49308
rect 53004 49198 53006 49250
rect 53058 49198 53060 49250
rect 53004 49186 53060 49198
rect 51548 49028 51604 49038
rect 51548 48934 51604 48972
rect 52780 49026 52836 49038
rect 52780 48974 52782 49026
rect 52834 48974 52836 49026
rect 50988 48750 50990 48802
rect 51042 48750 51044 48802
rect 50988 48738 51044 48750
rect 52108 48804 52164 48814
rect 52780 48804 52836 48974
rect 53228 49026 53284 50764
rect 53228 48974 53230 49026
rect 53282 48974 53284 49026
rect 53228 48962 53284 48974
rect 53116 48804 53172 48814
rect 52108 48802 52836 48804
rect 52108 48750 52110 48802
rect 52162 48750 52836 48802
rect 52108 48748 52836 48750
rect 53004 48802 53172 48804
rect 53004 48750 53118 48802
rect 53170 48750 53172 48802
rect 53004 48748 53172 48750
rect 50876 48078 50878 48130
rect 50930 48078 50932 48130
rect 50876 48066 50932 48078
rect 50092 47842 50148 47852
rect 50204 48018 50260 48030
rect 50204 47966 50206 48018
rect 50258 47966 50260 48018
rect 50204 47684 50260 47966
rect 49980 47628 50260 47684
rect 49980 45780 50036 47628
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50540 46676 50596 46686
rect 50540 46582 50596 46620
rect 50092 46562 50148 46574
rect 50092 46510 50094 46562
rect 50146 46510 50148 46562
rect 50092 46452 50148 46510
rect 51100 46564 51156 46574
rect 51100 46562 51380 46564
rect 51100 46510 51102 46562
rect 51154 46510 51380 46562
rect 51100 46508 51380 46510
rect 51100 46498 51156 46508
rect 50092 46386 50148 46396
rect 50652 46172 51044 46228
rect 50652 46002 50708 46172
rect 50652 45950 50654 46002
rect 50706 45950 50708 46002
rect 50652 45938 50708 45950
rect 50876 46002 50932 46014
rect 50876 45950 50878 46002
rect 50930 45950 50932 46002
rect 49980 45686 50036 45724
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50764 45220 50820 45230
rect 50876 45220 50932 45950
rect 50764 45218 50932 45220
rect 50764 45166 50766 45218
rect 50818 45166 50932 45218
rect 50764 45164 50932 45166
rect 50988 45666 51044 46172
rect 50988 45614 50990 45666
rect 51042 45614 51044 45666
rect 50988 45220 51044 45614
rect 50764 45154 50820 45164
rect 49980 45108 50036 45118
rect 49868 45052 49980 45108
rect 49980 45014 50036 45052
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 49308 43652 49476 43708
rect 48188 43428 48244 43438
rect 48188 43334 48244 43372
rect 48188 40628 48244 40638
rect 48076 40292 48132 40302
rect 48076 40198 48132 40236
rect 48188 38668 48244 40572
rect 48748 40402 48804 43652
rect 49084 41972 49140 43652
rect 49084 41906 49140 41916
rect 49196 41970 49252 41982
rect 49196 41918 49198 41970
rect 49250 41918 49252 41970
rect 48748 40350 48750 40402
rect 48802 40350 48804 40402
rect 48748 40338 48804 40350
rect 49196 40404 49252 41918
rect 49196 40338 49252 40348
rect 49308 40402 49364 40414
rect 49308 40350 49310 40402
rect 49362 40350 49364 40402
rect 49308 39844 49364 40350
rect 49084 39788 49364 39844
rect 48972 39396 49028 39406
rect 49084 39396 49140 39788
rect 48972 39394 49140 39396
rect 48972 39342 48974 39394
rect 49026 39342 49140 39394
rect 48972 39340 49140 39342
rect 49196 39618 49252 39630
rect 49196 39566 49198 39618
rect 49250 39566 49252 39618
rect 49196 39396 49252 39566
rect 49420 39396 49476 43652
rect 50092 42980 50148 42990
rect 50092 42978 50372 42980
rect 50092 42926 50094 42978
rect 50146 42926 50372 42978
rect 50092 42924 50372 42926
rect 50092 42914 50148 42924
rect 50204 42644 50260 42654
rect 50204 42550 50260 42588
rect 49644 42532 49700 42542
rect 50092 42532 50148 42542
rect 49644 42530 50148 42532
rect 49644 42478 49646 42530
rect 49698 42478 50094 42530
rect 50146 42478 50148 42530
rect 49644 42476 50148 42478
rect 49644 41972 49700 42476
rect 50092 42466 50148 42476
rect 49644 41906 49700 41916
rect 49868 41858 49924 41870
rect 49868 41806 49870 41858
rect 49922 41806 49924 41858
rect 49868 41412 49924 41806
rect 49868 41346 49924 41356
rect 50316 41410 50372 42924
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50316 41358 50318 41410
rect 50370 41358 50372 41410
rect 50316 41346 50372 41358
rect 50540 41412 50596 41422
rect 50540 41298 50596 41356
rect 50540 41246 50542 41298
rect 50594 41246 50596 41298
rect 50540 41234 50596 41246
rect 50540 40964 50596 40974
rect 50876 40964 50932 40974
rect 50540 40962 50876 40964
rect 50540 40910 50542 40962
rect 50594 40910 50876 40962
rect 50540 40908 50876 40910
rect 50540 40898 50596 40908
rect 50876 40898 50932 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50988 40516 51044 45164
rect 51212 45778 51268 45790
rect 51212 45726 51214 45778
rect 51266 45726 51268 45778
rect 51212 44546 51268 45726
rect 51212 44494 51214 44546
rect 51266 44494 51268 44546
rect 51212 44482 51268 44494
rect 51324 43708 51380 46508
rect 52108 46452 52164 48748
rect 53004 48354 53060 48748
rect 53116 48738 53172 48748
rect 53004 48302 53006 48354
rect 53058 48302 53060 48354
rect 53004 48290 53060 48302
rect 53340 48020 53396 52220
rect 53676 52164 53732 52782
rect 53676 52098 53732 52108
rect 54012 52722 54068 52734
rect 54012 52670 54014 52722
rect 54066 52670 54068 52722
rect 54012 50820 54068 52670
rect 54124 52164 54180 52174
rect 54124 52070 54180 52108
rect 54012 50754 54068 50764
rect 54236 50260 54292 53566
rect 54460 52946 54516 54236
rect 54572 54226 54628 54236
rect 54796 54180 54852 56028
rect 54908 56018 54964 56028
rect 55132 55970 55188 55982
rect 55132 55918 55134 55970
rect 55186 55918 55188 55970
rect 54908 55524 54964 55534
rect 54908 55300 54964 55468
rect 55132 55524 55188 55918
rect 55132 55458 55188 55468
rect 55244 55468 55300 56924
rect 55356 56914 55412 56924
rect 55580 56754 55636 56766
rect 55580 56702 55582 56754
rect 55634 56702 55636 56754
rect 55356 56642 55412 56654
rect 55356 56590 55358 56642
rect 55410 56590 55412 56642
rect 55356 55748 55412 56590
rect 55580 55858 55636 56702
rect 55580 55806 55582 55858
rect 55634 55806 55636 55858
rect 55580 55794 55636 55806
rect 55356 55692 55524 55748
rect 55468 55636 55524 55692
rect 55468 55580 55748 55636
rect 55692 55468 55748 55580
rect 56588 55468 56644 58492
rect 55244 55412 55412 55468
rect 55580 55412 55636 55422
rect 55692 55412 55860 55468
rect 55356 55410 55636 55412
rect 55356 55358 55582 55410
rect 55634 55358 55636 55410
rect 55356 55356 55636 55358
rect 55580 55346 55636 55356
rect 55020 55300 55076 55310
rect 54908 55298 55020 55300
rect 54908 55246 54910 55298
rect 54962 55246 55020 55298
rect 54908 55244 55020 55246
rect 54908 55206 54964 55244
rect 54796 53618 54852 54124
rect 54908 54292 54964 54302
rect 54908 53730 54964 54236
rect 54908 53678 54910 53730
rect 54962 53678 54964 53730
rect 54908 53666 54964 53678
rect 54796 53566 54798 53618
rect 54850 53566 54852 53618
rect 54796 53554 54852 53566
rect 55020 53172 55076 55244
rect 55132 54628 55188 54638
rect 55132 54402 55188 54572
rect 55132 54350 55134 54402
rect 55186 54350 55188 54402
rect 55132 54180 55188 54350
rect 55132 54114 55188 54124
rect 55804 54626 55860 55412
rect 55804 54574 55806 54626
rect 55858 54574 55860 54626
rect 55804 53844 55860 54574
rect 56476 55412 56532 55422
rect 56588 55412 56980 55468
rect 56476 54516 56532 55356
rect 56364 54514 56532 54516
rect 56364 54462 56478 54514
rect 56530 54462 56532 54514
rect 56364 54460 56532 54462
rect 55916 54402 55972 54414
rect 56140 54404 56196 54414
rect 55916 54350 55918 54402
rect 55970 54350 55972 54402
rect 55916 53844 55972 54350
rect 56028 54348 56140 54404
rect 56028 54290 56084 54348
rect 56140 54338 56196 54348
rect 56028 54238 56030 54290
rect 56082 54238 56084 54290
rect 56028 54226 56084 54238
rect 56028 53844 56084 53854
rect 55916 53842 56084 53844
rect 55916 53790 56030 53842
rect 56082 53790 56084 53842
rect 55916 53788 56084 53790
rect 55244 53730 55300 53742
rect 55244 53678 55246 53730
rect 55298 53678 55300 53730
rect 55244 53172 55300 53678
rect 55020 53170 55300 53172
rect 55020 53118 55022 53170
rect 55074 53118 55300 53170
rect 55020 53116 55300 53118
rect 55020 53106 55076 53116
rect 54460 52894 54462 52946
rect 54514 52894 54516 52946
rect 54460 52882 54516 52894
rect 54348 52722 54404 52734
rect 54348 52670 54350 52722
rect 54402 52670 54404 52722
rect 54348 51940 54404 52670
rect 55804 52388 55860 53788
rect 56028 53778 56084 53788
rect 56364 53284 56420 54460
rect 56476 54450 56532 54460
rect 56812 54628 56868 54638
rect 56812 54514 56868 54572
rect 56812 54462 56814 54514
rect 56866 54462 56868 54514
rect 56812 54450 56868 54462
rect 56700 54404 56756 54414
rect 56700 54310 56756 54348
rect 56252 53228 56420 53284
rect 55916 52388 55972 52398
rect 55804 52386 55972 52388
rect 55804 52334 55918 52386
rect 55970 52334 55972 52386
rect 55804 52332 55972 52334
rect 55916 52322 55972 52332
rect 56140 52388 56196 52398
rect 56140 52294 56196 52332
rect 56252 52386 56308 53228
rect 56252 52334 56254 52386
rect 56306 52334 56308 52386
rect 55132 52164 55188 52174
rect 56252 52164 56308 52334
rect 56588 52388 56644 52398
rect 56644 52332 56756 52388
rect 56588 52322 56644 52332
rect 54460 51940 54516 51950
rect 54348 51938 54516 51940
rect 54348 51886 54462 51938
rect 54514 51886 54516 51938
rect 54348 51884 54516 51886
rect 54460 51492 54516 51884
rect 54684 51492 54740 51502
rect 54460 51436 54684 51492
rect 54236 50204 54516 50260
rect 54460 49924 54516 50204
rect 54124 49026 54180 49038
rect 54124 48974 54126 49026
rect 54178 48974 54180 49026
rect 53900 48804 53956 48814
rect 54124 48804 54180 48974
rect 54460 49026 54516 49868
rect 54460 48974 54462 49026
rect 54514 48974 54516 49026
rect 54460 48962 54516 48974
rect 53900 48802 54180 48804
rect 53900 48750 53902 48802
rect 53954 48750 54180 48802
rect 53900 48748 54180 48750
rect 54684 48802 54740 51436
rect 55132 51378 55188 52108
rect 55916 52108 56308 52164
rect 55468 51604 55524 51614
rect 55468 51490 55524 51548
rect 55916 51602 55972 52108
rect 56252 51940 56308 51950
rect 55916 51550 55918 51602
rect 55970 51550 55972 51602
rect 55916 51538 55972 51550
rect 56028 51938 56308 51940
rect 56028 51886 56254 51938
rect 56306 51886 56308 51938
rect 56028 51884 56308 51886
rect 55468 51438 55470 51490
rect 55522 51438 55524 51490
rect 55468 51426 55524 51438
rect 55132 51326 55134 51378
rect 55186 51326 55188 51378
rect 55132 51314 55188 51326
rect 55356 51378 55412 51390
rect 55356 51326 55358 51378
rect 55410 51326 55412 51378
rect 55356 51268 55412 51326
rect 55244 50594 55300 50606
rect 55244 50542 55246 50594
rect 55298 50542 55300 50594
rect 54908 50372 54964 50382
rect 55244 50372 55300 50542
rect 54908 50370 55300 50372
rect 54908 50318 54910 50370
rect 54962 50318 55300 50370
rect 54908 50316 55300 50318
rect 54908 50306 54964 50316
rect 54908 49028 54964 49038
rect 54908 48934 54964 48972
rect 55020 49028 55076 50316
rect 55244 49028 55300 49038
rect 55020 49026 55300 49028
rect 55020 48974 55246 49026
rect 55298 48974 55300 49026
rect 55020 48972 55300 48974
rect 54684 48750 54686 48802
rect 54738 48750 54740 48802
rect 53900 48356 53956 48748
rect 54684 48692 54740 48750
rect 54684 48626 54740 48636
rect 54796 48802 54852 48814
rect 54796 48750 54798 48802
rect 54850 48750 54852 48802
rect 53900 48290 53956 48300
rect 54796 48356 54852 48750
rect 54796 48290 54852 48300
rect 52108 46386 52164 46396
rect 52332 47964 53396 48020
rect 53676 48242 53732 48254
rect 53676 48190 53678 48242
rect 53730 48190 53732 48242
rect 53676 48132 53732 48190
rect 54236 48132 54292 48142
rect 53676 48076 54236 48132
rect 51884 44996 51940 45006
rect 51772 44434 51828 44446
rect 51772 44382 51774 44434
rect 51826 44382 51828 44434
rect 51772 43764 51828 44382
rect 51324 43652 51492 43708
rect 50876 40460 51044 40516
rect 51436 42532 51492 43652
rect 50316 40404 50372 40414
rect 49756 39396 49812 39406
rect 49196 39394 49812 39396
rect 49196 39342 49758 39394
rect 49810 39342 49812 39394
rect 49196 39340 49812 39342
rect 48860 39284 48916 39294
rect 48972 39284 49028 39340
rect 48916 39228 49028 39284
rect 48860 39058 48916 39228
rect 48860 39006 48862 39058
rect 48914 39006 48916 39058
rect 48860 38994 48916 39006
rect 47964 28914 48020 28924
rect 48076 38612 48244 38668
rect 48076 26908 48132 38612
rect 48524 37940 48580 37950
rect 48524 37846 48580 37884
rect 48860 35028 48916 35038
rect 48860 34914 48916 34972
rect 48860 34862 48862 34914
rect 48914 34862 48916 34914
rect 48188 34802 48244 34814
rect 48188 34750 48190 34802
rect 48242 34750 48244 34802
rect 48188 34356 48244 34750
rect 48188 34290 48244 34300
rect 48300 33348 48356 33358
rect 48860 33348 48916 34862
rect 48300 33346 48916 33348
rect 48300 33294 48302 33346
rect 48354 33294 48916 33346
rect 48300 33292 48916 33294
rect 48300 31778 48356 33292
rect 49084 33234 49140 33246
rect 49084 33182 49086 33234
rect 49138 33182 49140 33234
rect 49084 32786 49140 33182
rect 49084 32734 49086 32786
rect 49138 32734 49140 32786
rect 49084 32722 49140 32734
rect 49196 32788 49252 39340
rect 49756 39330 49812 39340
rect 50316 38836 50372 40348
rect 50876 39956 50932 40460
rect 50988 40292 51044 40302
rect 50988 40290 51380 40292
rect 50988 40238 50990 40290
rect 51042 40238 51380 40290
rect 50988 40236 51380 40238
rect 50988 40226 51044 40236
rect 50652 39900 51156 39956
rect 50652 39730 50708 39900
rect 50652 39678 50654 39730
rect 50706 39678 50708 39730
rect 50652 39666 50708 39678
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 49756 38834 50372 38836
rect 49756 38782 50318 38834
rect 50370 38782 50372 38834
rect 49756 38780 50372 38782
rect 49420 38724 49476 38734
rect 49420 38630 49476 38668
rect 49308 38050 49364 38062
rect 49308 37998 49310 38050
rect 49362 37998 49364 38050
rect 49308 37828 49364 37998
rect 49756 37828 49812 38780
rect 50316 38770 50372 38780
rect 49308 37826 49812 37828
rect 49308 37774 49758 37826
rect 49810 37774 49812 37826
rect 49308 37772 49812 37774
rect 49308 36482 49364 37772
rect 49756 37762 49812 37772
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 49308 36430 49310 36482
rect 49362 36430 49364 36482
rect 49308 36418 49364 36430
rect 49980 36372 50036 36382
rect 49980 36370 50484 36372
rect 49980 36318 49982 36370
rect 50034 36318 50484 36370
rect 49980 36316 50484 36318
rect 49980 36306 50036 36316
rect 50428 35922 50484 36316
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50428 35870 50430 35922
rect 50482 35870 50484 35922
rect 50428 35858 50484 35870
rect 50764 35810 50820 35822
rect 50764 35758 50766 35810
rect 50818 35758 50820 35810
rect 50652 35700 50708 35710
rect 50764 35700 50820 35758
rect 50652 35698 50820 35700
rect 50652 35646 50654 35698
rect 50706 35646 50820 35698
rect 50652 35644 50820 35646
rect 50652 35634 50708 35644
rect 50316 35476 50372 35486
rect 49756 35028 49812 35038
rect 49980 35028 50036 35038
rect 49812 35026 50036 35028
rect 49812 34974 49982 35026
rect 50034 34974 50036 35026
rect 49812 34972 50036 34974
rect 49756 34962 49812 34972
rect 49980 34962 50036 34972
rect 49420 34804 49476 34814
rect 49420 34710 49476 34748
rect 49532 34804 49588 34814
rect 50316 34804 50372 35420
rect 50876 35252 50932 39900
rect 50988 39730 51044 39742
rect 50988 39678 50990 39730
rect 51042 39678 51044 39730
rect 50988 38946 51044 39678
rect 51100 39506 51156 39900
rect 51324 39842 51380 40236
rect 51324 39790 51326 39842
rect 51378 39790 51380 39842
rect 51324 39778 51380 39790
rect 51100 39454 51102 39506
rect 51154 39454 51156 39506
rect 51100 39442 51156 39454
rect 50988 38894 50990 38946
rect 51042 38894 51044 38946
rect 50988 38882 51044 38894
rect 51436 38668 51492 42476
rect 51548 43652 51828 43708
rect 51884 44322 51940 44940
rect 51884 44270 51886 44322
rect 51938 44270 51940 44322
rect 51548 42754 51604 43652
rect 51548 42702 51550 42754
rect 51602 42702 51604 42754
rect 51548 41074 51604 42702
rect 51660 42866 51716 42878
rect 51660 42814 51662 42866
rect 51714 42814 51716 42866
rect 51660 42644 51716 42814
rect 51772 42756 51828 42766
rect 51884 42756 51940 44270
rect 51772 42754 51940 42756
rect 51772 42702 51774 42754
rect 51826 42702 51940 42754
rect 51772 42700 51940 42702
rect 51772 42690 51828 42700
rect 51660 41636 51716 42588
rect 51660 41580 51828 41636
rect 51548 41022 51550 41074
rect 51602 41022 51604 41074
rect 51548 41010 51604 41022
rect 51660 40964 51716 40974
rect 51660 40870 51716 40908
rect 51660 40516 51716 40526
rect 51660 40402 51716 40460
rect 51660 40350 51662 40402
rect 51714 40350 51716 40402
rect 51660 40338 51716 40350
rect 51772 40290 51828 41580
rect 51884 41412 51940 42700
rect 51884 41186 51940 41356
rect 51884 41134 51886 41186
rect 51938 41134 51940 41186
rect 51884 41122 51940 41134
rect 51996 42530 52052 42542
rect 51996 42478 51998 42530
rect 52050 42478 52052 42530
rect 51996 41858 52052 42478
rect 51996 41806 51998 41858
rect 52050 41806 52052 41858
rect 51996 41300 52052 41806
rect 51996 41186 52052 41244
rect 51996 41134 51998 41186
rect 52050 41134 52052 41186
rect 51996 41122 52052 41134
rect 51772 40238 51774 40290
rect 51826 40238 51828 40290
rect 51772 40226 51828 40238
rect 51212 38612 51492 38668
rect 50988 35924 51044 35934
rect 51212 35924 51268 38612
rect 52332 36708 52388 47964
rect 52668 47460 52724 47470
rect 52668 47366 52724 47404
rect 53676 47460 53732 48076
rect 54236 48038 54292 48076
rect 54908 48132 54964 48142
rect 55020 48132 55076 48972
rect 55244 48962 55300 48972
rect 55356 49028 55412 51212
rect 56028 50706 56084 51884
rect 56252 51874 56308 51884
rect 56700 51602 56756 52332
rect 56700 51550 56702 51602
rect 56754 51550 56756 51602
rect 56700 51538 56756 51550
rect 56812 51492 56868 51502
rect 56476 51380 56532 51390
rect 56476 51286 56532 51324
rect 56812 51378 56868 51436
rect 56812 51326 56814 51378
rect 56866 51326 56868 51378
rect 56812 51314 56868 51326
rect 56028 50654 56030 50706
rect 56082 50654 56084 50706
rect 56028 50642 56084 50654
rect 55356 48962 55412 48972
rect 56140 49140 56196 49150
rect 56028 48916 56084 48926
rect 55916 48914 56084 48916
rect 55916 48862 56030 48914
rect 56082 48862 56084 48914
rect 55916 48860 56084 48862
rect 55692 48692 55748 48702
rect 55468 48356 55524 48366
rect 55468 48262 55524 48300
rect 55692 48354 55748 48636
rect 55916 48466 55972 48860
rect 56028 48850 56084 48860
rect 55916 48414 55918 48466
rect 55970 48414 55972 48466
rect 55916 48402 55972 48414
rect 55692 48302 55694 48354
rect 55746 48302 55748 48354
rect 55692 48290 55748 48302
rect 56140 48242 56196 49084
rect 56924 48468 56980 55412
rect 57708 55410 57764 55422
rect 57708 55358 57710 55410
rect 57762 55358 57764 55410
rect 57708 54628 57764 55358
rect 57708 54562 57764 54572
rect 57148 54514 57204 54526
rect 57148 54462 57150 54514
rect 57202 54462 57204 54514
rect 57148 54292 57204 54462
rect 57148 54226 57204 54236
rect 57372 52836 57428 52846
rect 57372 52742 57428 52780
rect 57596 52834 57652 52846
rect 57596 52782 57598 52834
rect 57650 52782 57652 52834
rect 57596 52276 57652 52782
rect 57596 52210 57652 52220
rect 57036 51604 57092 51614
rect 57036 51378 57092 51548
rect 57036 51326 57038 51378
rect 57090 51326 57092 51378
rect 57036 51314 57092 51326
rect 56924 48412 57092 48468
rect 56140 48190 56142 48242
rect 56194 48190 56196 48242
rect 56140 48178 56196 48190
rect 54964 48076 55076 48132
rect 54908 48038 54964 48076
rect 53676 47394 53732 47404
rect 56252 47460 56308 47470
rect 56252 47366 56308 47404
rect 53452 47348 53508 47358
rect 53452 47346 53620 47348
rect 53452 47294 53454 47346
rect 53506 47294 53620 47346
rect 53452 47292 53620 47294
rect 53452 47282 53508 47292
rect 53564 46898 53620 47292
rect 53564 46846 53566 46898
rect 53618 46846 53620 46898
rect 53564 46834 53620 46846
rect 55692 47234 55748 47246
rect 55692 47182 55694 47234
rect 55746 47182 55748 47234
rect 53340 46674 53396 46686
rect 53340 46622 53342 46674
rect 53394 46622 53396 46674
rect 53004 46564 53060 46574
rect 53340 46564 53396 46622
rect 53676 46676 53732 46686
rect 54124 46676 54180 46686
rect 53676 46674 54180 46676
rect 53676 46622 53678 46674
rect 53730 46622 54126 46674
rect 54178 46622 54180 46674
rect 53676 46620 54180 46622
rect 53676 46610 53732 46620
rect 54124 46610 54180 46620
rect 55020 46674 55076 46686
rect 55020 46622 55022 46674
rect 55074 46622 55076 46674
rect 53060 46508 53396 46564
rect 54908 46564 54964 46574
rect 53004 46470 53060 46508
rect 54908 46470 54964 46508
rect 54908 45892 54964 45902
rect 54908 45666 54964 45836
rect 54908 45614 54910 45666
rect 54962 45614 54964 45666
rect 53340 45108 53396 45118
rect 54908 45108 54964 45614
rect 55020 45332 55076 46622
rect 55692 46564 55748 47182
rect 55748 46508 55860 46564
rect 55692 46498 55748 46508
rect 55020 45266 55076 45276
rect 55244 46002 55300 46014
rect 55244 45950 55246 46002
rect 55298 45950 55300 46002
rect 53340 45014 53396 45052
rect 54796 45052 54908 45108
rect 55244 45108 55300 45950
rect 55692 45332 55748 45342
rect 55692 45218 55748 45276
rect 55692 45166 55694 45218
rect 55746 45166 55748 45218
rect 55692 45154 55748 45166
rect 55468 45108 55524 45118
rect 55244 45106 55524 45108
rect 55244 45054 55470 45106
rect 55522 45054 55524 45106
rect 55244 45052 55524 45054
rect 55804 45108 55860 46508
rect 55916 45332 55972 45342
rect 56924 45332 56980 45342
rect 55916 45330 56868 45332
rect 55916 45278 55918 45330
rect 55970 45278 56868 45330
rect 55916 45276 56868 45278
rect 55916 45266 55972 45276
rect 56028 45108 56084 45118
rect 56588 45108 56644 45118
rect 55804 45106 56084 45108
rect 55804 45054 56030 45106
rect 56082 45054 56084 45106
rect 55804 45052 56084 45054
rect 52892 44996 52948 45006
rect 52892 44902 52948 44940
rect 54572 44548 54628 44558
rect 54572 44454 54628 44492
rect 54236 44436 54292 44446
rect 53676 44434 54292 44436
rect 53676 44382 54238 44434
rect 54290 44382 54292 44434
rect 53676 44380 54292 44382
rect 53564 43652 53620 43662
rect 52780 43540 52836 43550
rect 52780 43446 52836 43484
rect 53228 43540 53284 43550
rect 53228 43446 53284 43484
rect 53564 42978 53620 43596
rect 53564 42926 53566 42978
rect 53618 42926 53620 42978
rect 53564 42914 53620 42926
rect 53676 42978 53732 44380
rect 54236 44370 54292 44380
rect 54348 44100 54404 44110
rect 54348 44006 54404 44044
rect 53676 42926 53678 42978
rect 53730 42926 53732 42978
rect 53676 42914 53732 42926
rect 54796 43426 54852 45052
rect 54908 45042 54964 45052
rect 55132 44996 55188 45006
rect 54908 44098 54964 44110
rect 54908 44046 54910 44098
rect 54962 44046 54964 44098
rect 54908 43764 54964 44046
rect 54908 43698 54964 43708
rect 54796 43374 54798 43426
rect 54850 43374 54852 43426
rect 53900 42754 53956 42766
rect 53900 42702 53902 42754
rect 53954 42702 53956 42754
rect 53116 42532 53172 42542
rect 53116 42438 53172 42476
rect 53900 42532 53956 42702
rect 53900 42466 53956 42476
rect 54012 42642 54068 42654
rect 54012 42590 54014 42642
rect 54066 42590 54068 42642
rect 54012 42196 54068 42590
rect 53788 42140 54068 42196
rect 53788 42082 53844 42140
rect 53788 42030 53790 42082
rect 53842 42030 53844 42082
rect 53788 42018 53844 42030
rect 52444 41972 52500 41982
rect 52444 41878 52500 41916
rect 53116 41972 53172 41982
rect 53116 41878 53172 41916
rect 53564 41972 53620 41982
rect 54796 41972 54852 43374
rect 55132 42532 55188 44940
rect 55244 44548 55300 44558
rect 55244 44454 55300 44492
rect 55356 44324 55412 45052
rect 55468 45042 55524 45052
rect 55356 42644 55412 44268
rect 55468 44322 55524 44334
rect 55468 44270 55470 44322
rect 55522 44270 55524 44322
rect 55468 44100 55524 44270
rect 56028 44212 56084 45052
rect 56140 45106 56644 45108
rect 56140 45054 56590 45106
rect 56642 45054 56644 45106
rect 56140 45052 56644 45054
rect 56140 44548 56196 45052
rect 56588 45042 56644 45052
rect 56812 45106 56868 45276
rect 56812 45054 56814 45106
rect 56866 45054 56868 45106
rect 56812 45042 56868 45054
rect 56924 44548 56980 45276
rect 57036 45108 57092 48412
rect 57372 45780 57428 45790
rect 57148 45778 57428 45780
rect 57148 45726 57374 45778
rect 57426 45726 57428 45778
rect 57148 45724 57428 45726
rect 57148 45218 57204 45724
rect 57372 45714 57428 45724
rect 57148 45166 57150 45218
rect 57202 45166 57204 45218
rect 57148 45154 57204 45166
rect 57036 45014 57092 45052
rect 56140 44454 56196 44492
rect 56364 44492 56980 44548
rect 56028 44146 56084 44156
rect 56252 44436 56308 44446
rect 55468 43708 55524 44044
rect 56252 43708 56308 44380
rect 55468 43652 55972 43708
rect 55916 42754 55972 43652
rect 55916 42702 55918 42754
rect 55970 42702 55972 42754
rect 55468 42644 55524 42654
rect 55356 42642 55524 42644
rect 55356 42590 55470 42642
rect 55522 42590 55524 42642
rect 55356 42588 55524 42590
rect 55468 42578 55524 42588
rect 55132 42466 55188 42476
rect 53620 41916 53732 41972
rect 53564 41906 53620 41916
rect 52892 41412 52948 41422
rect 52892 41318 52948 41356
rect 52668 41300 52724 41310
rect 52668 41206 52724 41244
rect 53116 41186 53172 41198
rect 53116 41134 53118 41186
rect 53170 41134 53172 41186
rect 53116 40516 53172 41134
rect 53564 40964 53620 40974
rect 53564 40870 53620 40908
rect 53116 38722 53172 40460
rect 53676 40404 53732 41916
rect 54796 41906 54852 41916
rect 55356 41860 55412 41870
rect 55356 41074 55412 41804
rect 55916 41858 55972 42702
rect 55916 41806 55918 41858
rect 55970 41806 55972 41858
rect 55916 41794 55972 41806
rect 56140 43652 56308 43708
rect 55356 41022 55358 41074
rect 55410 41022 55412 41074
rect 55356 41010 55412 41022
rect 55692 41186 55748 41198
rect 55692 41134 55694 41186
rect 55746 41134 55748 41186
rect 55692 40626 55748 41134
rect 55692 40574 55694 40626
rect 55746 40574 55748 40626
rect 55692 40562 55748 40574
rect 55916 40964 55972 40974
rect 55916 40516 55972 40908
rect 56028 40962 56084 40974
rect 56028 40910 56030 40962
rect 56082 40910 56084 40962
rect 56028 40628 56084 40910
rect 56028 40562 56084 40572
rect 55916 40422 55972 40460
rect 53676 39618 53732 40348
rect 53676 39566 53678 39618
rect 53730 39566 53732 39618
rect 53564 39060 53620 39070
rect 53676 39060 53732 39566
rect 53116 38670 53118 38722
rect 53170 38670 53172 38722
rect 53116 38658 53172 38670
rect 53340 39058 53732 39060
rect 53340 39006 53566 39058
rect 53618 39006 53732 39058
rect 53340 39004 53732 39006
rect 54012 40404 54068 40414
rect 52332 36642 52388 36652
rect 50988 35922 51268 35924
rect 50988 35870 50990 35922
rect 51042 35870 51214 35922
rect 51266 35870 51268 35922
rect 50988 35868 51268 35870
rect 50988 35858 51044 35868
rect 51212 35858 51268 35868
rect 52108 36594 52164 36606
rect 52108 36542 52110 36594
rect 52162 36542 52164 36594
rect 52108 35700 52164 36542
rect 52892 36596 52948 36606
rect 53340 36596 53396 39004
rect 53564 38994 53620 39004
rect 53676 38724 53732 38734
rect 53900 38724 53956 38734
rect 53732 38722 53956 38724
rect 53732 38670 53902 38722
rect 53954 38670 53956 38722
rect 53732 38668 53956 38670
rect 53564 37828 53620 37838
rect 53676 37828 53732 38668
rect 53900 38658 53956 38668
rect 53564 37826 53732 37828
rect 53564 37774 53566 37826
rect 53618 37774 53732 37826
rect 53564 37772 53732 37774
rect 53564 37762 53620 37772
rect 52892 36594 53396 36596
rect 52892 36542 52894 36594
rect 52946 36542 53396 36594
rect 52892 36540 53396 36542
rect 52892 36530 52948 36540
rect 53340 36482 53396 36540
rect 53340 36430 53342 36482
rect 53394 36430 53396 36482
rect 53340 36418 53396 36430
rect 52892 35700 52948 35710
rect 52108 35698 52948 35700
rect 52108 35646 52110 35698
rect 52162 35646 52894 35698
rect 52946 35646 52948 35698
rect 52108 35644 52948 35646
rect 52108 35634 52164 35644
rect 52892 35634 52948 35644
rect 51996 35586 52052 35598
rect 51996 35534 51998 35586
rect 52050 35534 52052 35586
rect 51772 35476 51828 35486
rect 51772 35382 51828 35420
rect 50876 35186 50932 35196
rect 49532 34802 50372 34804
rect 49532 34750 49534 34802
rect 49586 34750 50372 34802
rect 49532 34748 50372 34750
rect 49532 34738 49588 34748
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 51212 33460 51268 33470
rect 51996 33460 52052 35534
rect 53116 35476 53172 35486
rect 53452 35476 53508 35486
rect 53116 35382 53172 35420
rect 53228 35474 53508 35476
rect 53228 35422 53454 35474
rect 53506 35422 53508 35474
rect 53228 35420 53508 35422
rect 53228 34914 53284 35420
rect 53452 35410 53508 35420
rect 53228 34862 53230 34914
rect 53282 34862 53284 34914
rect 51212 33458 51716 33460
rect 51212 33406 51214 33458
rect 51266 33406 51716 33458
rect 51212 33404 51716 33406
rect 51996 33404 52276 33460
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51212 32788 51268 33404
rect 49196 32732 49588 32788
rect 48972 32564 49028 32574
rect 48972 32470 49028 32508
rect 49196 32562 49252 32574
rect 49196 32510 49198 32562
rect 49250 32510 49252 32562
rect 48300 31726 48302 31778
rect 48354 31726 48356 31778
rect 48300 31556 48356 31726
rect 49196 31780 49252 32510
rect 49532 31892 49588 32732
rect 50652 32732 51268 32788
rect 51548 33234 51604 33246
rect 51548 33182 51550 33234
rect 51602 33182 51604 33234
rect 50652 32674 50708 32732
rect 50652 32622 50654 32674
rect 50706 32622 50708 32674
rect 50652 32610 50708 32622
rect 49644 32564 49700 32574
rect 49644 32470 49700 32508
rect 50316 32562 50372 32574
rect 50316 32510 50318 32562
rect 50370 32510 50372 32562
rect 49868 32002 49924 32014
rect 49868 31950 49870 32002
rect 49922 31950 49924 32002
rect 49532 31836 49700 31892
rect 49308 31780 49364 31790
rect 49196 31724 49308 31780
rect 49308 31686 49364 31724
rect 49420 31668 49476 31678
rect 49420 31574 49476 31612
rect 49532 31666 49588 31678
rect 49532 31614 49534 31666
rect 49586 31614 49588 31666
rect 48748 31556 48804 31566
rect 48300 31554 48804 31556
rect 48300 31502 48750 31554
rect 48802 31502 48804 31554
rect 48300 31500 48804 31502
rect 48748 30212 48804 31500
rect 48972 31556 49028 31566
rect 48972 31218 49028 31500
rect 49532 31556 49588 31614
rect 49532 31490 49588 31500
rect 48972 31166 48974 31218
rect 49026 31166 49028 31218
rect 48972 31154 49028 31166
rect 48748 30146 48804 30156
rect 49084 30098 49140 30110
rect 49084 30046 49086 30098
rect 49138 30046 49140 30098
rect 49084 29652 49140 30046
rect 49084 29586 49140 29596
rect 49644 28868 49700 31836
rect 49868 30882 49924 31950
rect 50316 31948 50372 32510
rect 50428 32564 50484 32574
rect 50428 32470 50484 32508
rect 50876 32562 50932 32574
rect 50876 32510 50878 32562
rect 50930 32510 50932 32562
rect 50092 31892 50148 31902
rect 50316 31892 50484 31948
rect 50092 31778 50148 31836
rect 50092 31726 50094 31778
rect 50146 31726 50148 31778
rect 50092 31714 50148 31726
rect 50428 31780 50484 31892
rect 50876 31892 50932 32510
rect 51436 32450 51492 32462
rect 51436 32398 51438 32450
rect 51490 32398 51492 32450
rect 51436 32116 51492 32398
rect 51436 32050 51492 32060
rect 51548 31892 51604 33182
rect 51660 32564 51716 33404
rect 51884 33348 51940 33358
rect 51884 33254 51940 33292
rect 51996 33236 52052 33246
rect 51996 33142 52052 33180
rect 52108 33234 52164 33246
rect 52108 33182 52110 33234
rect 52162 33182 52164 33234
rect 52108 32900 52164 33182
rect 51772 32844 52164 32900
rect 51772 32786 51828 32844
rect 51772 32734 51774 32786
rect 51826 32734 51828 32786
rect 51772 32722 51828 32734
rect 51996 32674 52052 32686
rect 51996 32622 51998 32674
rect 52050 32622 52052 32674
rect 51996 32564 52052 32622
rect 52108 32676 52164 32686
rect 52220 32676 52276 33404
rect 52780 33346 52836 33358
rect 52780 33294 52782 33346
rect 52834 33294 52836 33346
rect 52108 32674 52220 32676
rect 52108 32622 52110 32674
rect 52162 32622 52220 32674
rect 52108 32620 52220 32622
rect 52108 32610 52164 32620
rect 52220 32582 52276 32620
rect 52668 32676 52724 32686
rect 51660 32508 52052 32564
rect 51772 31892 51828 31902
rect 51548 31836 51772 31892
rect 50876 31826 50932 31836
rect 50428 31554 50484 31724
rect 50428 31502 50430 31554
rect 50482 31502 50484 31554
rect 49868 30830 49870 30882
rect 49922 30830 49924 30882
rect 49868 30818 49924 30830
rect 49980 31106 50036 31118
rect 49980 31054 49982 31106
rect 50034 31054 50036 31106
rect 49980 30324 50036 31054
rect 50204 30772 50260 30782
rect 50204 30678 50260 30716
rect 50428 30548 50484 31502
rect 50764 31556 50820 31594
rect 50820 31500 50932 31556
rect 50764 31490 50820 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50876 30772 50932 31500
rect 50876 30706 50932 30716
rect 49868 30212 49924 30222
rect 49868 30118 49924 30156
rect 49980 29988 50036 30268
rect 50204 30492 50484 30548
rect 50204 30210 50260 30492
rect 51548 30436 51604 30446
rect 50204 30158 50206 30210
rect 50258 30158 50260 30210
rect 50204 30146 50260 30158
rect 50876 30212 50932 30222
rect 50876 30100 50932 30156
rect 51548 30212 51604 30380
rect 51772 30324 51828 31836
rect 52668 31332 52724 32620
rect 52780 32116 52836 33294
rect 52892 32676 52948 32686
rect 52892 32674 53172 32676
rect 52892 32622 52894 32674
rect 52946 32622 53172 32674
rect 52892 32620 53172 32622
rect 52892 32610 52948 32620
rect 52780 32050 52836 32060
rect 53116 31556 53172 32620
rect 53228 32674 53284 34862
rect 53452 34692 53508 34702
rect 53452 34598 53508 34636
rect 53452 33236 53508 33246
rect 53452 33142 53508 33180
rect 53228 32622 53230 32674
rect 53282 32622 53284 32674
rect 53228 32610 53284 32622
rect 52668 31276 52836 31332
rect 51548 30210 51716 30212
rect 51548 30158 51550 30210
rect 51602 30158 51716 30210
rect 51548 30156 51716 30158
rect 51548 30146 51604 30156
rect 50876 30044 51380 30100
rect 50316 29988 50372 29998
rect 49980 29986 50372 29988
rect 49980 29934 50318 29986
rect 50370 29934 50372 29986
rect 49980 29932 50372 29934
rect 50316 29922 50372 29932
rect 50540 29988 50596 29998
rect 50540 29986 51268 29988
rect 50540 29934 50542 29986
rect 50594 29934 51268 29986
rect 50540 29932 51268 29934
rect 50540 29922 50596 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 51100 29652 51156 29662
rect 51100 29558 51156 29596
rect 50988 29428 51044 29438
rect 50988 29334 51044 29372
rect 51212 29426 51268 29932
rect 51212 29374 51214 29426
rect 51266 29374 51268 29426
rect 51212 29362 51268 29374
rect 48524 28756 48580 28766
rect 48524 28662 48580 28700
rect 49532 28756 49588 28766
rect 49644 28756 49700 28812
rect 50652 28868 50708 28878
rect 49532 28754 49700 28756
rect 49532 28702 49534 28754
rect 49586 28702 49700 28754
rect 49532 28700 49700 28702
rect 49756 28756 49812 28766
rect 49532 28690 49588 28700
rect 49756 28662 49812 28700
rect 50652 28754 50708 28812
rect 50652 28702 50654 28754
rect 50706 28702 50708 28754
rect 50652 28690 50708 28702
rect 51324 28756 51380 30044
rect 51548 29540 51604 29550
rect 51548 29446 51604 29484
rect 51436 28756 51492 28766
rect 51324 28700 51436 28756
rect 50092 28420 50148 28430
rect 50092 28326 50148 28364
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50316 27860 50372 27870
rect 48076 26852 48356 26908
rect 47852 26450 47908 26460
rect 48188 26292 48244 26302
rect 47628 26290 48244 26292
rect 47628 26238 47630 26290
rect 47682 26238 48190 26290
rect 48242 26238 48244 26290
rect 47628 26236 48244 26238
rect 47628 26226 47684 26236
rect 48188 26226 48244 26236
rect 47292 26066 47348 26078
rect 47292 26014 47294 26066
rect 47346 26014 47348 26066
rect 46956 25618 47012 25630
rect 46956 25566 46958 25618
rect 47010 25566 47012 25618
rect 46620 25508 46676 25518
rect 46620 25414 46676 25452
rect 46956 25396 47012 25566
rect 47292 25508 47348 26014
rect 47628 26068 47684 26078
rect 47628 25974 47684 26012
rect 47292 25442 47348 25452
rect 46956 25330 47012 25340
rect 46172 24894 46174 24946
rect 46226 24894 46228 24946
rect 45276 24610 45780 24612
rect 45276 24558 45278 24610
rect 45330 24558 45780 24610
rect 45276 24556 45780 24558
rect 45276 24500 45332 24556
rect 45276 24434 45332 24444
rect 44604 24052 44660 24062
rect 44604 23378 44660 23996
rect 45500 24052 45556 24062
rect 45500 23938 45556 23996
rect 45500 23886 45502 23938
rect 45554 23886 45556 23938
rect 45500 23874 45556 23886
rect 46172 23938 46228 24894
rect 48300 24612 48356 26852
rect 49084 26068 49140 26078
rect 49084 25618 49140 26012
rect 50316 25620 50372 27804
rect 51436 27860 51492 28700
rect 51660 28420 51716 30156
rect 51772 30098 51828 30268
rect 52668 30324 52724 30334
rect 52668 30210 52724 30268
rect 52668 30158 52670 30210
rect 52722 30158 52724 30210
rect 52668 30146 52724 30158
rect 51772 30046 51774 30098
rect 51826 30046 51828 30098
rect 51772 30034 51828 30046
rect 51660 28354 51716 28364
rect 52780 28642 52836 31276
rect 53004 29986 53060 29998
rect 53004 29934 53006 29986
rect 53058 29934 53060 29986
rect 53004 29540 53060 29934
rect 53116 29652 53172 31500
rect 53228 29988 53284 29998
rect 53228 29652 53284 29932
rect 53116 29650 53284 29652
rect 53116 29598 53118 29650
rect 53170 29598 53284 29650
rect 53116 29596 53284 29598
rect 53116 29586 53172 29596
rect 53452 29540 53508 29550
rect 53004 28756 53060 29484
rect 53340 29538 53508 29540
rect 53340 29486 53454 29538
rect 53506 29486 53508 29538
rect 53340 29484 53508 29486
rect 53228 29428 53284 29438
rect 53004 28700 53172 28756
rect 52780 28590 52782 28642
rect 52834 28590 52836 28642
rect 52780 27972 52836 28590
rect 52780 27906 52836 27916
rect 53004 28532 53060 28542
rect 53004 28418 53060 28476
rect 53004 28366 53006 28418
rect 53058 28366 53060 28418
rect 51436 27766 51492 27804
rect 52108 27746 52164 27758
rect 52108 27694 52110 27746
rect 52162 27694 52164 27746
rect 52108 26964 52164 27694
rect 53004 27524 53060 28366
rect 53116 28308 53172 28700
rect 53228 28642 53284 29372
rect 53228 28590 53230 28642
rect 53282 28590 53284 28642
rect 53228 28578 53284 28590
rect 53116 28252 53284 28308
rect 52668 27468 53060 27524
rect 52556 27074 52612 27086
rect 52556 27022 52558 27074
rect 52610 27022 52612 27074
rect 52556 26908 52612 27022
rect 52108 26898 52164 26908
rect 52332 26852 52612 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 52332 26514 52388 26852
rect 52668 26628 52724 27468
rect 53228 27188 53284 28252
rect 53340 27860 53396 29484
rect 53452 29474 53508 29484
rect 53564 28532 53620 28542
rect 53564 28438 53620 28476
rect 53340 27794 53396 27804
rect 53452 28418 53508 28430
rect 53452 28366 53454 28418
rect 53506 28366 53508 28418
rect 53452 27748 53508 28366
rect 53676 28308 53732 37772
rect 54012 37044 54068 40348
rect 56028 40402 56084 40414
rect 56028 40350 56030 40402
rect 56082 40350 56084 40402
rect 56028 40292 56084 40350
rect 56028 40226 56084 40236
rect 54348 39508 54404 39518
rect 54236 39506 54404 39508
rect 54236 39454 54350 39506
rect 54402 39454 54404 39506
rect 54236 39452 54404 39454
rect 54124 39060 54180 39070
rect 54124 38966 54180 39004
rect 54236 38722 54292 39452
rect 54348 39442 54404 39452
rect 54236 38670 54238 38722
rect 54290 38670 54292 38722
rect 54236 38658 54292 38670
rect 56140 38668 56196 43652
rect 56364 39508 56420 44492
rect 56588 44324 56644 44334
rect 56588 44230 56644 44268
rect 56924 44322 56980 44492
rect 57596 44994 57652 45006
rect 57596 44942 57598 44994
rect 57650 44942 57652 44994
rect 57596 44436 57652 44942
rect 57596 44370 57652 44380
rect 57708 44546 57764 44558
rect 57708 44494 57710 44546
rect 57762 44494 57764 44546
rect 56924 44270 56926 44322
rect 56978 44270 56980 44322
rect 56924 44258 56980 44270
rect 56700 44212 56756 44222
rect 56700 43708 56756 44156
rect 57596 44212 57652 44222
rect 57708 44212 57764 44494
rect 57596 44210 57764 44212
rect 57596 44158 57598 44210
rect 57650 44158 57764 44210
rect 57596 44156 57764 44158
rect 57596 43708 57652 44156
rect 56476 43652 56756 43708
rect 57372 43652 57652 43708
rect 56476 42754 56532 43652
rect 57372 43650 57428 43652
rect 57372 43598 57374 43650
rect 57426 43598 57428 43650
rect 57372 43586 57428 43598
rect 57820 43650 57876 59052
rect 57932 55468 57988 60732
rect 58044 60564 58100 60574
rect 58044 60470 58100 60508
rect 58044 60004 58100 60014
rect 58044 59910 58100 59948
rect 58156 59220 58212 59230
rect 58156 58548 58212 59164
rect 58268 58548 58324 58558
rect 58156 58546 58324 58548
rect 58156 58494 58270 58546
rect 58322 58494 58324 58546
rect 58156 58492 58324 58494
rect 58268 58482 58324 58492
rect 57932 55412 58324 55468
rect 58156 55300 58212 55310
rect 58156 55206 58212 55244
rect 58156 54292 58212 54302
rect 58156 53842 58212 54236
rect 58156 53790 58158 53842
rect 58210 53790 58212 53842
rect 58156 53778 58212 53790
rect 58156 52946 58212 52958
rect 58156 52894 58158 52946
rect 58210 52894 58212 52946
rect 58156 52836 58212 52894
rect 58156 52276 58212 52780
rect 58156 52210 58212 52220
rect 58156 51604 58212 51614
rect 58156 50706 58212 51548
rect 58156 50654 58158 50706
rect 58210 50654 58212 50706
rect 58156 50642 58212 50654
rect 58156 49140 58212 49150
rect 58156 49046 58212 49084
rect 58044 45892 58100 45902
rect 58044 45798 58100 45836
rect 58268 45556 58324 55412
rect 58044 45500 58324 45556
rect 58044 44546 58100 45500
rect 58156 45332 58212 45342
rect 58212 45276 58324 45332
rect 58156 45238 58212 45276
rect 58044 44494 58046 44546
rect 58098 44494 58100 44546
rect 58044 44482 58100 44494
rect 58268 44434 58324 45276
rect 58268 44382 58270 44434
rect 58322 44382 58324 44434
rect 58268 44370 58324 44382
rect 57820 43598 57822 43650
rect 57874 43598 57876 43650
rect 57148 43426 57204 43438
rect 57148 43374 57150 43426
rect 57202 43374 57204 43426
rect 56476 42702 56478 42754
rect 56530 42702 56532 42754
rect 56476 42690 56532 42702
rect 57036 42866 57092 42878
rect 57036 42814 57038 42866
rect 57090 42814 57092 42866
rect 56924 42644 56980 42654
rect 56588 42642 56980 42644
rect 56588 42590 56926 42642
rect 56978 42590 56980 42642
rect 56588 42588 56980 42590
rect 56476 39732 56532 39742
rect 56588 39732 56644 42588
rect 56924 42578 56980 42588
rect 57036 42082 57092 42814
rect 57036 42030 57038 42082
rect 57090 42030 57092 42082
rect 56700 41860 56756 41870
rect 57036 41860 57092 42030
rect 57148 42084 57204 43374
rect 57148 42028 57652 42084
rect 57372 41970 57428 42028
rect 57372 41918 57374 41970
rect 57426 41918 57428 41970
rect 57372 41906 57428 41918
rect 56756 41804 56868 41860
rect 56700 41766 56756 41804
rect 56700 40516 56756 40526
rect 56700 40422 56756 40460
rect 56812 40292 56868 41804
rect 57036 41794 57092 41804
rect 57484 41858 57540 41870
rect 57484 41806 57486 41858
rect 57538 41806 57540 41858
rect 57260 41188 57316 41198
rect 57260 41074 57316 41132
rect 57260 41022 57262 41074
rect 57314 41022 57316 41074
rect 57260 41010 57316 41022
rect 56476 39730 56644 39732
rect 56476 39678 56478 39730
rect 56530 39678 56644 39730
rect 56476 39676 56644 39678
rect 56476 39666 56532 39676
rect 56588 39620 56644 39676
rect 56588 39554 56644 39564
rect 56700 40236 56868 40292
rect 56924 40404 56980 40414
rect 56924 40290 56980 40348
rect 56924 40238 56926 40290
rect 56978 40238 56980 40290
rect 56364 39442 56420 39452
rect 55692 38612 56196 38668
rect 56700 38722 56756 40236
rect 56924 40226 56980 40238
rect 57036 40402 57092 40414
rect 57036 40350 57038 40402
rect 57090 40350 57092 40402
rect 57036 40292 57092 40350
rect 57484 40402 57540 41806
rect 57484 40350 57486 40402
rect 57538 40350 57540 40402
rect 57484 40338 57540 40350
rect 57596 41186 57652 42028
rect 57596 41134 57598 41186
rect 57650 41134 57652 41186
rect 57036 39844 57092 40236
rect 57484 39844 57540 39854
rect 57036 39842 57540 39844
rect 57036 39790 57486 39842
rect 57538 39790 57540 39842
rect 57036 39788 57540 39790
rect 57484 39778 57540 39788
rect 57036 39620 57092 39630
rect 57036 39526 57092 39564
rect 56812 39508 56868 39518
rect 56812 39414 56868 39452
rect 57596 39506 57652 41134
rect 57708 41972 57764 41982
rect 57820 41972 57876 43598
rect 58156 41972 58212 41982
rect 57708 41970 58212 41972
rect 57708 41918 57710 41970
rect 57762 41918 58158 41970
rect 58210 41918 58212 41970
rect 57708 41916 58212 41918
rect 57708 41188 57764 41916
rect 57764 41132 57876 41188
rect 57708 41122 57764 41132
rect 57820 39842 57876 41132
rect 58156 40626 58212 41916
rect 58156 40574 58158 40626
rect 58210 40574 58212 40626
rect 58156 40562 58212 40574
rect 57820 39790 57822 39842
rect 57874 39790 57876 39842
rect 57820 39778 57876 39790
rect 57596 39454 57598 39506
rect 57650 39454 57652 39506
rect 57596 39442 57652 39454
rect 57820 38946 57876 38958
rect 57820 38894 57822 38946
rect 57874 38894 57876 38946
rect 56700 38670 56702 38722
rect 56754 38670 56756 38722
rect 54908 38052 54964 38062
rect 54908 37958 54964 37996
rect 55356 38052 55412 38062
rect 55356 37958 55412 37996
rect 54012 36978 54068 36988
rect 54012 36372 54068 36382
rect 54012 36370 55188 36372
rect 54012 36318 54014 36370
rect 54066 36318 55188 36370
rect 54012 36316 55188 36318
rect 54012 36306 54068 36316
rect 55132 35922 55188 36316
rect 55132 35870 55134 35922
rect 55186 35870 55188 35922
rect 55132 35858 55188 35870
rect 54908 35700 54964 35710
rect 54684 35698 54964 35700
rect 54684 35646 54910 35698
rect 54962 35646 54964 35698
rect 54684 35644 54964 35646
rect 54012 34692 54068 34702
rect 53788 33348 53844 33358
rect 53788 32340 53844 33292
rect 53900 32788 53956 32798
rect 53900 32694 53956 32732
rect 54012 32674 54068 34636
rect 54684 34354 54740 35644
rect 54908 35634 54964 35644
rect 55356 35698 55412 35710
rect 55356 35646 55358 35698
rect 55410 35646 55412 35698
rect 55356 34916 55412 35646
rect 55580 35698 55636 35710
rect 55580 35646 55582 35698
rect 55634 35646 55636 35698
rect 55580 35588 55636 35646
rect 55580 35522 55636 35532
rect 55692 35252 55748 38612
rect 56700 38052 56756 38670
rect 57596 38724 57652 38734
rect 57596 38630 57652 38668
rect 57820 38388 57876 38894
rect 58156 38834 58212 38846
rect 58156 38782 58158 38834
rect 58210 38782 58212 38834
rect 58156 38724 58212 38782
rect 58156 38612 58212 38668
rect 58156 38546 58212 38556
rect 57820 38332 58324 38388
rect 56028 37940 56084 37950
rect 56028 37938 56644 37940
rect 56028 37886 56030 37938
rect 56082 37886 56644 37938
rect 56028 37884 56644 37886
rect 56028 37874 56084 37884
rect 56140 36596 56196 36606
rect 56140 36594 56420 36596
rect 56140 36542 56142 36594
rect 56194 36542 56420 36594
rect 56140 36540 56420 36542
rect 56140 36530 56196 36540
rect 55580 35196 55748 35252
rect 55468 34916 55524 34926
rect 55356 34914 55524 34916
rect 55356 34862 55470 34914
rect 55522 34862 55524 34914
rect 55356 34860 55524 34862
rect 55468 34850 55524 34860
rect 54684 34302 54686 34354
rect 54738 34302 54740 34354
rect 54684 34290 54740 34302
rect 54908 34242 54964 34254
rect 54908 34190 54910 34242
rect 54962 34190 54964 34242
rect 54908 32788 54964 34190
rect 55020 34244 55076 34254
rect 55020 34130 55076 34188
rect 55020 34078 55022 34130
rect 55074 34078 55076 34130
rect 55020 33348 55076 34078
rect 55580 33684 55636 35196
rect 56364 35028 56420 36540
rect 56588 35924 56644 37884
rect 56700 36594 56756 37996
rect 56700 36542 56702 36594
rect 56754 36542 56756 36594
rect 56700 36530 56756 36542
rect 58156 38218 58212 38230
rect 58156 38166 58158 38218
rect 58210 38166 58212 38218
rect 56812 35924 56868 35934
rect 56588 35922 56868 35924
rect 56588 35870 56814 35922
rect 56866 35870 56868 35922
rect 56588 35868 56868 35870
rect 56812 35858 56868 35868
rect 56924 35924 56980 35934
rect 56028 34972 56420 35028
rect 55804 34802 55860 34814
rect 55804 34750 55806 34802
rect 55858 34750 55860 34802
rect 55692 34690 55748 34702
rect 55692 34638 55694 34690
rect 55746 34638 55748 34690
rect 55692 34468 55748 34638
rect 55804 34692 55860 34750
rect 55804 34626 55860 34636
rect 56028 34468 56084 34972
rect 55692 34412 56084 34468
rect 56252 34804 56308 34814
rect 56252 34244 56308 34748
rect 56364 34802 56420 34972
rect 56588 35698 56644 35710
rect 56588 35646 56590 35698
rect 56642 35646 56644 35698
rect 56588 34914 56644 35646
rect 56588 34862 56590 34914
rect 56642 34862 56644 34914
rect 56588 34850 56644 34862
rect 56364 34750 56366 34802
rect 56418 34750 56420 34802
rect 56364 34738 56420 34750
rect 56924 34802 56980 35868
rect 57708 35924 57764 35934
rect 58156 35924 58212 38166
rect 57764 35868 58212 35924
rect 57708 35830 57764 35868
rect 57036 35700 57092 35710
rect 57036 35606 57092 35644
rect 57148 35698 57204 35710
rect 57148 35646 57150 35698
rect 57202 35646 57204 35698
rect 57148 35588 57204 35646
rect 56924 34750 56926 34802
rect 56978 34750 56980 34802
rect 56924 34738 56980 34750
rect 57036 34804 57092 34814
rect 57036 34710 57092 34748
rect 56252 34178 56308 34188
rect 56700 34690 56756 34702
rect 56700 34638 56702 34690
rect 56754 34638 56756 34690
rect 56700 34242 56756 34638
rect 57148 34356 57204 35532
rect 57596 35698 57652 35710
rect 57596 35646 57598 35698
rect 57650 35646 57652 35698
rect 56700 34190 56702 34242
rect 56754 34190 56756 34242
rect 56700 34178 56756 34190
rect 56924 34300 57204 34356
rect 56812 34020 56868 34030
rect 55020 32788 55076 33292
rect 55468 33628 55636 33684
rect 56140 34018 56868 34020
rect 56140 33966 56814 34018
rect 56866 33966 56868 34018
rect 56140 33964 56868 33966
rect 55132 32788 55188 32798
rect 55020 32786 55188 32788
rect 55020 32734 55134 32786
rect 55186 32734 55188 32786
rect 55020 32732 55188 32734
rect 54908 32722 54964 32732
rect 55132 32722 55188 32732
rect 54012 32622 54014 32674
rect 54066 32622 54068 32674
rect 54012 32610 54068 32622
rect 54796 32676 54852 32686
rect 54796 32582 54852 32620
rect 53900 32340 53956 32350
rect 53788 32338 53956 32340
rect 53788 32286 53902 32338
rect 53954 32286 53956 32338
rect 53788 32284 53956 32286
rect 53900 32274 53956 32284
rect 55244 32116 55300 32126
rect 55244 31778 55300 32060
rect 55244 31726 55246 31778
rect 55298 31726 55300 31778
rect 55132 30994 55188 31006
rect 55132 30942 55134 30994
rect 55186 30942 55188 30994
rect 55132 30436 55188 30942
rect 54572 29988 54628 29998
rect 54572 29894 54628 29932
rect 54908 29988 54964 29998
rect 54908 29894 54964 29932
rect 53900 29314 53956 29326
rect 53900 29262 53902 29314
rect 53954 29262 53956 29314
rect 53900 28644 53956 29262
rect 53900 28578 53956 28588
rect 54236 28644 54292 28654
rect 54236 28550 54292 28588
rect 55132 28532 55188 30380
rect 55244 30212 55300 31726
rect 55356 31106 55412 31118
rect 55356 31054 55358 31106
rect 55410 31054 55412 31106
rect 55356 30996 55412 31054
rect 55356 30930 55412 30940
rect 55356 30212 55412 30222
rect 55244 30210 55412 30212
rect 55244 30158 55358 30210
rect 55410 30158 55412 30210
rect 55244 30156 55412 30158
rect 55132 28466 55188 28476
rect 55356 28756 55412 30156
rect 53452 27682 53508 27692
rect 53564 28252 53732 28308
rect 52892 27132 53284 27188
rect 52780 26964 52836 27002
rect 52780 26898 52836 26908
rect 52332 26462 52334 26514
rect 52386 26462 52388 26514
rect 52332 26450 52388 26462
rect 52444 26572 52724 26628
rect 52444 26180 52500 26572
rect 49084 25566 49086 25618
rect 49138 25566 49140 25618
rect 49084 25554 49140 25566
rect 49868 25618 50372 25620
rect 49868 25566 50318 25618
rect 50370 25566 50372 25618
rect 49868 25564 50372 25566
rect 49868 25508 49924 25564
rect 49532 25506 49924 25508
rect 49532 25454 49870 25506
rect 49922 25454 49924 25506
rect 49532 25452 49924 25454
rect 49532 24722 49588 25452
rect 49868 25442 49924 25452
rect 50204 25284 50260 25294
rect 50204 24834 50260 25228
rect 50204 24782 50206 24834
rect 50258 24782 50260 24834
rect 50204 24770 50260 24782
rect 49532 24670 49534 24722
rect 49586 24670 49588 24722
rect 49532 24658 49588 24670
rect 48300 24546 48356 24556
rect 48748 24612 48804 24622
rect 46172 23886 46174 23938
rect 46226 23886 46228 23938
rect 46172 23874 46228 23886
rect 44940 23714 44996 23726
rect 44940 23662 44942 23714
rect 44994 23662 44996 23714
rect 44940 23604 44996 23662
rect 45836 23714 45892 23726
rect 45836 23662 45838 23714
rect 45890 23662 45892 23714
rect 44940 23538 44996 23548
rect 45388 23604 45444 23614
rect 44604 23326 44606 23378
rect 44658 23326 44660 23378
rect 44604 23314 44660 23326
rect 45052 23380 45108 23390
rect 44940 23268 44996 23278
rect 44940 23174 44996 23212
rect 45052 22482 45108 23324
rect 45052 22430 45054 22482
rect 45106 22430 45108 22482
rect 45052 22418 45108 22430
rect 45388 23154 45444 23548
rect 45836 23492 45892 23662
rect 45836 23426 45892 23436
rect 46508 23714 46564 23726
rect 46508 23662 46510 23714
rect 46562 23662 46564 23714
rect 45388 23102 45390 23154
rect 45442 23102 45444 23154
rect 45388 22484 45444 23102
rect 45612 23268 45668 23278
rect 45500 22484 45556 22494
rect 45388 22482 45556 22484
rect 45388 22430 45502 22482
rect 45554 22430 45556 22482
rect 45388 22428 45556 22430
rect 45500 22418 45556 22428
rect 45612 22372 45668 23212
rect 46060 23044 46116 23054
rect 45836 23042 46116 23044
rect 45836 22990 46062 23042
rect 46114 22990 46116 23042
rect 45836 22988 46116 22990
rect 45388 22260 45444 22270
rect 45388 21474 45444 22204
rect 45388 21422 45390 21474
rect 45442 21422 45444 21474
rect 44492 18358 44548 18396
rect 44604 20020 44660 20030
rect 44604 19348 44660 19964
rect 45276 20020 45332 20030
rect 45388 20020 45444 21422
rect 45332 19964 45444 20020
rect 45276 19954 45332 19964
rect 43932 18162 43988 18172
rect 44268 17892 44324 17902
rect 44268 17778 44324 17836
rect 44268 17726 44270 17778
rect 44322 17726 44324 17778
rect 44268 17714 44324 17726
rect 44268 17444 44324 17454
rect 43708 14306 43876 14308
rect 43708 14254 43710 14306
rect 43762 14254 43876 14306
rect 43708 14252 43876 14254
rect 43708 14242 43764 14252
rect 43708 13636 43764 13646
rect 43708 13542 43764 13580
rect 43820 13636 43876 14252
rect 44044 14532 44100 14542
rect 44044 13858 44100 14476
rect 44044 13806 44046 13858
rect 44098 13806 44100 13858
rect 44044 13794 44100 13806
rect 44156 13858 44212 13870
rect 44156 13806 44158 13858
rect 44210 13806 44212 13858
rect 44156 13636 44212 13806
rect 43820 13580 44212 13636
rect 43708 12964 43764 12974
rect 43708 12870 43764 12908
rect 43820 12516 43876 13580
rect 44156 13412 44212 13422
rect 43484 12338 43540 12348
rect 43708 12460 43876 12516
rect 43932 13356 44156 13412
rect 42588 11732 42980 11788
rect 43260 11732 43428 11788
rect 42588 9940 42644 11732
rect 43036 11508 43092 11518
rect 42812 11452 43036 11508
rect 42812 10834 42868 11452
rect 42812 10782 42814 10834
rect 42866 10782 42868 10834
rect 42812 10770 42868 10782
rect 43036 10612 43092 11452
rect 43148 10612 43204 10622
rect 43036 10556 43148 10612
rect 43148 10518 43204 10556
rect 42588 9846 42644 9884
rect 43036 10164 43092 10174
rect 43036 9826 43092 10108
rect 43036 9774 43038 9826
rect 43090 9774 43092 9826
rect 43036 9762 43092 9774
rect 42476 9650 42532 9660
rect 43260 9380 43316 11732
rect 43484 9828 43540 9838
rect 43708 9828 43764 12460
rect 43932 12068 43988 13356
rect 44156 13346 44212 13356
rect 44044 12738 44100 12750
rect 44044 12686 44046 12738
rect 44098 12686 44100 12738
rect 44044 12628 44100 12686
rect 44044 12562 44100 12572
rect 43820 12012 43988 12068
rect 43820 10052 43876 12012
rect 44156 11956 44212 11966
rect 43932 11954 44212 11956
rect 43932 11902 44158 11954
rect 44210 11902 44212 11954
rect 43932 11900 44212 11902
rect 43932 10722 43988 11900
rect 44156 11890 44212 11900
rect 44268 10836 44324 17388
rect 44380 13746 44436 13758
rect 44380 13694 44382 13746
rect 44434 13694 44436 13746
rect 44380 13188 44436 13694
rect 44604 13524 44660 19292
rect 44716 19906 44772 19918
rect 44716 19854 44718 19906
rect 44770 19854 44772 19906
rect 44716 19012 44772 19854
rect 45612 19234 45668 22316
rect 45612 19182 45614 19234
rect 45666 19182 45668 19234
rect 45612 19170 45668 19182
rect 45724 22484 45780 22494
rect 44716 18564 44772 18956
rect 45276 19010 45332 19022
rect 45276 18958 45278 19010
rect 45330 18958 45332 19010
rect 45276 18676 45332 18958
rect 45276 18610 45332 18620
rect 44716 18498 44772 18508
rect 45052 18452 45108 18462
rect 44940 18450 45108 18452
rect 44940 18398 45054 18450
rect 45106 18398 45108 18450
rect 44940 18396 45108 18398
rect 44940 17668 44996 18396
rect 45052 18386 45108 18396
rect 45724 18116 45780 22428
rect 45836 22482 45892 22988
rect 46060 22978 46116 22988
rect 46508 23044 46564 23662
rect 46508 22978 46564 22988
rect 46620 23714 46676 23726
rect 46620 23662 46622 23714
rect 46674 23662 46676 23714
rect 45836 22430 45838 22482
rect 45890 22430 45892 22482
rect 45836 22418 45892 22430
rect 45948 22370 46004 22382
rect 45948 22318 45950 22370
rect 46002 22318 46004 22370
rect 45948 22260 46004 22318
rect 46284 22372 46340 22382
rect 46620 22372 46676 23662
rect 46732 23716 46788 23726
rect 46732 23714 46900 23716
rect 46732 23662 46734 23714
rect 46786 23662 46900 23714
rect 46732 23660 46900 23662
rect 46732 23650 46788 23660
rect 46844 23492 46900 23660
rect 46284 22370 46676 22372
rect 46284 22318 46286 22370
rect 46338 22318 46676 22370
rect 46284 22316 46676 22318
rect 46732 22372 46788 22382
rect 46284 22306 46340 22316
rect 45948 22194 46004 22204
rect 46396 22148 46452 22158
rect 46396 21810 46452 22092
rect 46396 21758 46398 21810
rect 46450 21758 46452 21810
rect 46284 20020 46340 20030
rect 46284 19906 46340 19964
rect 46284 19854 46286 19906
rect 46338 19854 46340 19906
rect 46172 19460 46228 19470
rect 46172 19234 46228 19404
rect 46172 19182 46174 19234
rect 46226 19182 46228 19234
rect 46172 19170 46228 19182
rect 45948 19122 46004 19134
rect 45948 19070 45950 19122
rect 46002 19070 46004 19122
rect 45836 19010 45892 19022
rect 45836 18958 45838 19010
rect 45890 18958 45892 19010
rect 45836 18562 45892 18958
rect 45948 18676 46004 19070
rect 45948 18610 46004 18620
rect 45836 18510 45838 18562
rect 45890 18510 45892 18562
rect 45836 18498 45892 18510
rect 45724 18050 45780 18060
rect 44940 17574 44996 17612
rect 45276 17892 45332 17902
rect 45052 15876 45108 15886
rect 45052 15426 45108 15820
rect 45052 15374 45054 15426
rect 45106 15374 45108 15426
rect 45052 15362 45108 15374
rect 45276 15314 45332 17836
rect 45388 15876 45444 15886
rect 45388 15782 45444 15820
rect 45724 15876 45780 15886
rect 45724 15782 45780 15820
rect 45276 15262 45278 15314
rect 45330 15262 45332 15314
rect 45276 15250 45332 15262
rect 45612 15316 45668 15326
rect 45724 15316 45780 15326
rect 45612 15314 45724 15316
rect 45612 15262 45614 15314
rect 45666 15262 45724 15314
rect 45612 15260 45724 15262
rect 44716 15204 44772 15242
rect 45164 15202 45220 15214
rect 45164 15150 45166 15202
rect 45218 15150 45220 15202
rect 45164 15148 45220 15150
rect 44716 15138 44772 15148
rect 45052 15092 45220 15148
rect 44716 14532 44772 14542
rect 44716 14438 44772 14476
rect 45052 14532 45108 15092
rect 45052 14530 45220 14532
rect 45052 14478 45054 14530
rect 45106 14478 45220 14530
rect 45052 14476 45220 14478
rect 45052 14466 45108 14476
rect 44940 14306 44996 14318
rect 44940 14254 44942 14306
rect 44994 14254 44996 14306
rect 44940 13860 44996 14254
rect 44940 13794 44996 13804
rect 45164 13858 45220 14476
rect 45164 13806 45166 13858
rect 45218 13806 45220 13858
rect 45164 13794 45220 13806
rect 44604 13458 44660 13468
rect 44940 13634 44996 13646
rect 44940 13582 44942 13634
rect 44994 13582 44996 13634
rect 44828 13188 44884 13198
rect 44380 13186 44884 13188
rect 44380 13134 44830 13186
rect 44882 13134 44884 13186
rect 44380 13132 44884 13134
rect 44828 13122 44884 13132
rect 44940 13186 44996 13582
rect 44940 13134 44942 13186
rect 44994 13134 44996 13186
rect 44940 13122 44996 13134
rect 45612 12964 45668 15260
rect 45724 15250 45780 15260
rect 46284 15148 46340 19854
rect 46396 15540 46452 21758
rect 46620 20132 46676 20142
rect 46732 20132 46788 22316
rect 46844 21588 46900 23436
rect 48748 23380 48804 24556
rect 50316 23604 50372 25564
rect 52220 26124 52500 26180
rect 52556 26402 52612 26414
rect 52556 26350 52558 26402
rect 52610 26350 52612 26402
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 52220 24724 52276 26124
rect 52556 25956 52612 26350
rect 52668 26402 52724 26572
rect 52668 26350 52670 26402
rect 52722 26350 52724 26402
rect 52668 26338 52724 26350
rect 52220 24658 52276 24668
rect 52332 25900 52612 25956
rect 52332 25396 52388 25900
rect 52332 24610 52388 25340
rect 52556 25506 52612 25518
rect 52892 25508 52948 27132
rect 53228 27074 53284 27132
rect 53228 27022 53230 27074
rect 53282 27022 53284 27074
rect 53228 27010 53284 27022
rect 53004 26962 53060 26974
rect 53004 26910 53006 26962
rect 53058 26910 53060 26962
rect 53004 26908 53060 26910
rect 53452 26962 53508 26974
rect 53452 26910 53454 26962
rect 53506 26910 53508 26962
rect 53452 26908 53508 26910
rect 53004 26852 53508 26908
rect 52556 25454 52558 25506
rect 52610 25454 52612 25506
rect 52556 24946 52612 25454
rect 52556 24894 52558 24946
rect 52610 24894 52612 24946
rect 52556 24882 52612 24894
rect 52668 25452 52948 25508
rect 52332 24558 52334 24610
rect 52386 24558 52388 24610
rect 52332 24546 52388 24558
rect 52668 23938 52724 25452
rect 52780 25284 52836 25294
rect 52892 25284 52948 25452
rect 53004 25564 53396 25620
rect 53004 25506 53060 25564
rect 53004 25454 53006 25506
rect 53058 25454 53060 25506
rect 53004 25442 53060 25454
rect 53340 25508 53396 25564
rect 53452 25508 53508 25518
rect 53340 25506 53508 25508
rect 53340 25454 53454 25506
rect 53506 25454 53508 25506
rect 53340 25452 53508 25454
rect 53452 25442 53508 25452
rect 53228 25394 53284 25406
rect 53228 25342 53230 25394
rect 53282 25342 53284 25394
rect 53228 25284 53284 25342
rect 52892 25228 53284 25284
rect 52780 25190 52836 25228
rect 52780 24834 52836 24846
rect 53564 24836 53620 28252
rect 54684 28084 54740 28094
rect 55356 28084 55412 28700
rect 55468 28196 55524 33628
rect 55580 33458 55636 33470
rect 55580 33406 55582 33458
rect 55634 33406 55636 33458
rect 55580 32788 55636 33406
rect 55580 32722 55636 32732
rect 56028 33122 56084 33134
rect 56028 33070 56030 33122
rect 56082 33070 56084 33122
rect 56028 32116 56084 33070
rect 56028 32050 56084 32060
rect 56028 31892 56084 31902
rect 56140 31892 56196 33964
rect 56812 33954 56868 33964
rect 56924 32900 56980 34300
rect 57036 34130 57092 34142
rect 57036 34078 57038 34130
rect 57090 34078 57092 34130
rect 57036 33570 57092 34078
rect 57148 34130 57204 34300
rect 57148 34078 57150 34130
rect 57202 34078 57204 34130
rect 57148 34066 57204 34078
rect 57260 34692 57316 34702
rect 57260 33908 57316 34636
rect 57596 34692 57652 35646
rect 57932 35700 57988 35710
rect 57932 35606 57988 35644
rect 57596 34626 57652 34636
rect 57036 33518 57038 33570
rect 57090 33518 57092 33570
rect 57036 33506 57092 33518
rect 57148 33852 57316 33908
rect 57148 33346 57204 33852
rect 57596 33572 57652 33582
rect 57148 33294 57150 33346
rect 57202 33294 57204 33346
rect 57148 33282 57204 33294
rect 57260 33570 57652 33572
rect 57260 33518 57598 33570
rect 57650 33518 57652 33570
rect 57260 33516 57652 33518
rect 57036 33124 57092 33134
rect 57036 33030 57092 33068
rect 56924 32844 57092 32900
rect 56028 31890 56196 31892
rect 56028 31838 56030 31890
rect 56082 31838 56196 31890
rect 56028 31836 56196 31838
rect 56028 31826 56084 31836
rect 56924 31220 56980 31230
rect 56028 31218 56980 31220
rect 56028 31166 56926 31218
rect 56978 31166 56980 31218
rect 56028 31164 56980 31166
rect 56028 30322 56084 31164
rect 56924 31154 56980 31164
rect 56588 30996 56644 31006
rect 56812 30996 56868 31006
rect 56588 30902 56644 30940
rect 56700 30994 56868 30996
rect 56700 30942 56814 30994
rect 56866 30942 56868 30994
rect 56700 30940 56868 30942
rect 56028 30270 56030 30322
rect 56082 30270 56084 30322
rect 56028 30258 56084 30270
rect 56700 29650 56756 30940
rect 56812 30930 56868 30940
rect 56924 30996 56980 31006
rect 57036 30996 57092 32844
rect 56980 30940 57092 30996
rect 57260 30994 57316 33516
rect 57596 33506 57652 33516
rect 57484 33348 57540 33358
rect 57484 33254 57540 33292
rect 57596 33124 57652 33134
rect 57596 31892 57652 33068
rect 58156 32450 58212 32462
rect 58156 32398 58158 32450
rect 58210 32398 58212 32450
rect 58156 32116 58212 32398
rect 58156 32050 58212 32060
rect 58156 31892 58212 31902
rect 57596 31890 58212 31892
rect 57596 31838 58158 31890
rect 58210 31838 58212 31890
rect 57596 31836 58212 31838
rect 58156 31826 58212 31836
rect 58156 31444 58212 31454
rect 57820 31108 57876 31118
rect 58156 31108 58212 31388
rect 57820 31014 57876 31052
rect 57932 31106 58212 31108
rect 57932 31054 58158 31106
rect 58210 31054 58212 31106
rect 57932 31052 58212 31054
rect 57260 30942 57262 30994
rect 57314 30942 57316 30994
rect 56924 30930 56980 30940
rect 57260 30930 57316 30942
rect 57036 29988 57092 29998
rect 56700 29598 56702 29650
rect 56754 29598 56756 29650
rect 56700 29586 56756 29598
rect 56924 29652 56980 29662
rect 56924 29558 56980 29596
rect 57036 29538 57092 29932
rect 57484 29988 57540 29998
rect 57540 29932 57652 29988
rect 57484 29922 57540 29932
rect 57036 29486 57038 29538
rect 57090 29486 57092 29538
rect 57036 29474 57092 29486
rect 57372 29652 57428 29662
rect 56588 28756 56644 28794
rect 56588 28690 56644 28700
rect 55468 28130 55524 28140
rect 56588 28532 56644 28542
rect 54684 28082 55412 28084
rect 54684 28030 54686 28082
rect 54738 28030 55412 28082
rect 54684 28028 55412 28030
rect 54684 28018 54740 28028
rect 53676 27860 53732 27870
rect 53676 27076 53732 27804
rect 55132 27860 55188 27870
rect 55132 27766 55188 27804
rect 54236 27748 54292 27758
rect 53788 27076 53844 27086
rect 53676 27074 53844 27076
rect 53676 27022 53790 27074
rect 53842 27022 53844 27074
rect 53676 27020 53844 27022
rect 53676 26852 53732 26862
rect 53676 26758 53732 26796
rect 53788 25506 53844 27020
rect 54236 26964 54292 27692
rect 54236 26898 54292 26908
rect 55020 27300 55076 27310
rect 53788 25454 53790 25506
rect 53842 25454 53844 25506
rect 53676 25396 53732 25406
rect 53676 25302 53732 25340
rect 52780 24782 52782 24834
rect 52834 24782 52836 24834
rect 52780 24052 52836 24782
rect 53116 24780 53620 24836
rect 52892 24724 52948 24734
rect 52892 24630 52948 24668
rect 52780 23986 52836 23996
rect 52668 23886 52670 23938
rect 52722 23886 52724 23938
rect 52668 23874 52724 23886
rect 52892 23828 52948 23838
rect 52892 23734 52948 23772
rect 51436 23716 51492 23726
rect 50316 23548 50484 23604
rect 48748 23314 48804 23324
rect 47964 23156 48020 23166
rect 47516 22482 47572 22494
rect 47516 22430 47518 22482
rect 47570 22430 47572 22482
rect 47068 22258 47124 22270
rect 47068 22206 47070 22258
rect 47122 22206 47124 22258
rect 46956 22146 47012 22158
rect 46956 22094 46958 22146
rect 47010 22094 47012 22146
rect 46956 21812 47012 22094
rect 46956 21746 47012 21756
rect 47068 21810 47124 22206
rect 47180 22258 47236 22270
rect 47180 22206 47182 22258
rect 47234 22206 47236 22258
rect 47180 22148 47236 22206
rect 47516 22148 47572 22430
rect 47964 22370 48020 23100
rect 50428 23156 50484 23548
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 51436 23266 51492 23660
rect 53004 23716 53060 23726
rect 53004 23622 53060 23660
rect 53116 23548 53172 24780
rect 53340 24610 53396 24622
rect 53340 24558 53342 24610
rect 53394 24558 53396 24610
rect 53228 23940 53284 23950
rect 53228 23846 53284 23884
rect 53004 23492 53172 23548
rect 51436 23214 51438 23266
rect 51490 23214 51492 23266
rect 51436 23202 51492 23214
rect 52220 23268 52276 23278
rect 50428 23090 50484 23100
rect 50764 23154 50820 23166
rect 50764 23102 50766 23154
rect 50818 23102 50820 23154
rect 48188 23044 48244 23054
rect 48188 22484 48244 22988
rect 50764 23044 50820 23102
rect 50764 22978 50820 22988
rect 51212 23044 51268 23054
rect 48188 22418 48244 22428
rect 50204 22484 50260 22494
rect 47964 22318 47966 22370
rect 48018 22318 48020 22370
rect 47964 22306 48020 22318
rect 48636 22260 48692 22270
rect 48076 22258 48692 22260
rect 48076 22206 48638 22258
rect 48690 22206 48692 22258
rect 48076 22204 48692 22206
rect 48076 22148 48132 22204
rect 48636 22194 48692 22204
rect 47516 22092 48132 22148
rect 47180 22082 47236 22092
rect 49084 21924 49140 21934
rect 47068 21758 47070 21810
rect 47122 21758 47124 21810
rect 47068 21746 47124 21758
rect 47292 21812 47348 21822
rect 47292 21810 47908 21812
rect 47292 21758 47294 21810
rect 47346 21758 47908 21810
rect 47292 21756 47908 21758
rect 47292 21746 47348 21756
rect 47404 21588 47460 21598
rect 46844 21586 47572 21588
rect 46844 21534 47406 21586
rect 47458 21534 47572 21586
rect 46844 21532 47572 21534
rect 47404 21522 47460 21532
rect 46620 20130 46788 20132
rect 46620 20078 46622 20130
rect 46674 20078 46788 20130
rect 46620 20076 46788 20078
rect 47292 20578 47348 20590
rect 47292 20526 47294 20578
rect 47346 20526 47348 20578
rect 46620 20066 46676 20076
rect 46844 20020 46900 20030
rect 46844 19926 46900 19964
rect 47068 20018 47124 20030
rect 47068 19966 47070 20018
rect 47122 19966 47124 20018
rect 46732 19908 46788 19918
rect 46732 19814 46788 19852
rect 46956 19796 47012 19806
rect 46732 18564 46788 18574
rect 46620 17444 46676 17454
rect 46620 17350 46676 17388
rect 46396 15484 46564 15540
rect 46172 15092 46340 15148
rect 45724 12964 45780 12974
rect 45612 12962 46116 12964
rect 45612 12910 45726 12962
rect 45778 12910 46116 12962
rect 45612 12908 46116 12910
rect 45724 12898 45780 12908
rect 45500 12852 45556 12862
rect 45500 12758 45556 12796
rect 45276 12738 45332 12750
rect 45276 12686 45278 12738
rect 45330 12686 45332 12738
rect 45276 12628 45332 12686
rect 45276 12562 45332 12572
rect 45612 12738 45668 12750
rect 45612 12686 45614 12738
rect 45666 12686 45668 12738
rect 44716 12292 44772 12302
rect 44716 12198 44772 12236
rect 45612 12292 45668 12686
rect 45612 12226 45668 12236
rect 44380 11956 44436 11966
rect 44604 11956 44660 11966
rect 44380 11954 44660 11956
rect 44380 11902 44382 11954
rect 44434 11902 44606 11954
rect 44658 11902 44660 11954
rect 44380 11900 44660 11902
rect 44380 11890 44436 11900
rect 44604 11890 44660 11900
rect 43932 10670 43934 10722
rect 43986 10670 43988 10722
rect 43932 10658 43988 10670
rect 44156 10780 44324 10836
rect 43820 9996 43988 10052
rect 43484 9826 43764 9828
rect 43484 9774 43486 9826
rect 43538 9774 43764 9826
rect 43484 9772 43764 9774
rect 43820 9828 43876 9838
rect 43484 9762 43540 9772
rect 41916 9324 42308 9380
rect 41916 9266 41972 9324
rect 41916 9214 41918 9266
rect 41970 9214 41972 9266
rect 41916 9202 41972 9214
rect 42140 9154 42196 9166
rect 42140 9102 42142 9154
rect 42194 9102 42196 9154
rect 42140 8260 42196 9102
rect 42252 9044 42308 9324
rect 42924 9324 43316 9380
rect 42812 9156 42868 9166
rect 42812 9062 42868 9100
rect 42364 9044 42420 9054
rect 42252 9042 42420 9044
rect 42252 8990 42366 9042
rect 42418 8990 42420 9042
rect 42252 8988 42420 8990
rect 42364 8978 42420 8988
rect 42140 8194 42196 8204
rect 41468 7858 41524 7868
rect 42924 8148 42980 9324
rect 43596 9268 43652 9772
rect 43820 9734 43876 9772
rect 43596 9202 43652 9212
rect 43148 9156 43204 9166
rect 40908 7756 41412 7812
rect 40012 7700 40068 7710
rect 40012 7606 40068 7644
rect 40124 7588 40180 7598
rect 40124 7494 40180 7532
rect 39900 7410 39956 7420
rect 40348 7474 40404 7486
rect 40348 7422 40350 7474
rect 40402 7422 40404 7474
rect 39676 7186 39732 7196
rect 40236 6692 40292 6702
rect 40236 6598 40292 6636
rect 40012 6578 40068 6590
rect 40012 6526 40014 6578
rect 40066 6526 40068 6578
rect 40012 6356 40068 6526
rect 40012 6290 40068 6300
rect 40124 6466 40180 6478
rect 40124 6414 40126 6466
rect 40178 6414 40180 6466
rect 40124 5796 40180 6414
rect 40348 6356 40404 7422
rect 40796 7476 40852 7486
rect 40796 7382 40852 7420
rect 40796 6916 40852 6926
rect 40796 6822 40852 6860
rect 40908 6914 40964 7756
rect 41356 7698 41412 7756
rect 41356 7646 41358 7698
rect 41410 7646 41412 7698
rect 41356 7634 41412 7646
rect 41468 7700 41524 7710
rect 42588 7700 42644 7710
rect 42924 7700 42980 8092
rect 41524 7644 41636 7700
rect 41468 7606 41524 7644
rect 41244 7476 41300 7514
rect 41244 7410 41300 7420
rect 40908 6862 40910 6914
rect 40962 6862 40964 6914
rect 40908 6850 40964 6862
rect 41580 6914 41636 7644
rect 42588 7698 42980 7700
rect 42588 7646 42590 7698
rect 42642 7646 42926 7698
rect 42978 7646 42980 7698
rect 42588 7644 42980 7646
rect 42588 7634 42644 7644
rect 42924 7634 42980 7644
rect 43036 9154 43204 9156
rect 43036 9102 43150 9154
rect 43202 9102 43204 9154
rect 43036 9100 43204 9102
rect 41580 6862 41582 6914
rect 41634 6862 41636 6914
rect 41580 6850 41636 6862
rect 41692 7588 41748 7598
rect 41244 6804 41300 6814
rect 41244 6710 41300 6748
rect 40572 6692 40628 6702
rect 40572 6578 40628 6636
rect 40572 6526 40574 6578
rect 40626 6526 40628 6578
rect 40572 6514 40628 6526
rect 40348 6290 40404 6300
rect 40124 5740 40740 5796
rect 39452 5282 39508 5292
rect 39900 5348 39956 5358
rect 39900 5236 39956 5292
rect 40348 5236 40404 5246
rect 39900 5234 40404 5236
rect 39900 5182 40350 5234
rect 40402 5182 40404 5234
rect 39900 5180 40404 5182
rect 38220 5124 38276 5134
rect 38220 4562 38276 5068
rect 39116 5124 39172 5134
rect 39116 5030 39172 5068
rect 39900 5122 39956 5180
rect 40348 5170 40404 5180
rect 40684 5234 40740 5740
rect 41244 5794 41300 5806
rect 41244 5742 41246 5794
rect 41298 5742 41300 5794
rect 40684 5182 40686 5234
rect 40738 5182 40740 5234
rect 40684 5170 40740 5182
rect 40908 5348 40964 5358
rect 39900 5070 39902 5122
rect 39954 5070 39956 5122
rect 39900 5058 39956 5070
rect 38220 4510 38222 4562
rect 38274 4510 38276 4562
rect 38220 4498 38276 4510
rect 40796 4898 40852 4910
rect 40796 4846 40798 4898
rect 40850 4846 40852 4898
rect 38108 4398 38110 4450
rect 38162 4398 38164 4450
rect 38108 4386 38164 4398
rect 40796 4452 40852 4846
rect 40796 4386 40852 4396
rect 37212 4286 37214 4338
rect 37266 4286 37268 4338
rect 37212 4274 37268 4286
rect 40908 4338 40964 5292
rect 41244 5348 41300 5742
rect 41580 5796 41636 5806
rect 41692 5796 41748 7532
rect 41804 7476 41860 7486
rect 41804 6802 41860 7420
rect 41804 6750 41806 6802
rect 41858 6750 41860 6802
rect 41804 6580 41860 6750
rect 42924 6692 42980 6702
rect 43036 6692 43092 9100
rect 43148 9090 43204 9100
rect 43484 9156 43540 9166
rect 43820 9156 43876 9166
rect 43484 9062 43540 9100
rect 43708 9154 43876 9156
rect 43708 9102 43822 9154
rect 43874 9102 43876 9154
rect 43708 9100 43876 9102
rect 43708 8036 43764 9100
rect 43820 9090 43876 9100
rect 43596 7700 43652 7710
rect 43708 7700 43764 7980
rect 43596 7698 43764 7700
rect 43596 7646 43598 7698
rect 43650 7646 43764 7698
rect 43596 7644 43764 7646
rect 43596 7634 43652 7644
rect 43260 7586 43316 7598
rect 43260 7534 43262 7586
rect 43314 7534 43316 7586
rect 43260 7140 43316 7534
rect 43820 7588 43876 7598
rect 43820 7494 43876 7532
rect 43260 6804 43316 7084
rect 43708 7362 43764 7374
rect 43708 7310 43710 7362
rect 43762 7310 43764 7362
rect 43708 6916 43764 7310
rect 43260 6738 43316 6748
rect 43484 6860 43764 6916
rect 42924 6690 43036 6692
rect 42924 6638 42926 6690
rect 42978 6638 43036 6690
rect 42924 6636 43036 6638
rect 42924 6626 42980 6636
rect 43036 6598 43092 6636
rect 43484 6690 43540 6860
rect 43932 6692 43988 9996
rect 44156 9714 44212 10780
rect 44156 9662 44158 9714
rect 44210 9662 44212 9714
rect 44156 7474 44212 9662
rect 44268 10612 44324 10622
rect 44268 9268 44324 10556
rect 46060 10498 46116 12908
rect 46060 10446 46062 10498
rect 46114 10446 46116 10498
rect 46060 10434 46116 10446
rect 46172 10276 46228 15092
rect 45612 10220 46228 10276
rect 44268 9266 44660 9268
rect 44268 9214 44270 9266
rect 44322 9214 44660 9266
rect 44268 9212 44660 9214
rect 44268 9202 44324 9212
rect 44156 7422 44158 7474
rect 44210 7422 44212 7474
rect 44156 7362 44212 7422
rect 44156 7310 44158 7362
rect 44210 7310 44212 7362
rect 44156 7298 44212 7310
rect 43484 6638 43486 6690
rect 43538 6638 43540 6690
rect 43484 6626 43540 6638
rect 43596 6690 43988 6692
rect 43596 6638 43934 6690
rect 43986 6638 43988 6690
rect 43596 6636 43988 6638
rect 41804 6514 41860 6524
rect 43260 6578 43316 6590
rect 43260 6526 43262 6578
rect 43314 6526 43316 6578
rect 43148 6466 43204 6478
rect 43148 6414 43150 6466
rect 43202 6414 43204 6466
rect 43148 6132 43204 6414
rect 43260 6244 43316 6526
rect 43596 6244 43652 6636
rect 43260 6188 43652 6244
rect 43820 6468 43876 6478
rect 43148 6076 43764 6132
rect 43708 6018 43764 6076
rect 43708 5966 43710 6018
rect 43762 5966 43764 6018
rect 43708 5954 43764 5966
rect 41580 5794 41748 5796
rect 41580 5742 41582 5794
rect 41634 5742 41748 5794
rect 41580 5740 41748 5742
rect 41580 5730 41636 5740
rect 41244 5282 41300 5292
rect 41692 4452 41748 4462
rect 41692 4358 41748 4396
rect 40908 4286 40910 4338
rect 40962 4286 40964 4338
rect 40908 4274 40964 4286
rect 34300 4226 35140 4228
rect 34300 4174 34302 4226
rect 34354 4174 35140 4226
rect 34300 4172 35140 4174
rect 43820 4226 43876 6412
rect 43932 6244 43988 6636
rect 43932 6178 43988 6188
rect 44380 5908 44436 9212
rect 44604 9042 44660 9212
rect 44604 8990 44606 9042
rect 44658 8990 44660 9042
rect 44604 8978 44660 8990
rect 45388 8930 45444 8942
rect 45388 8878 45390 8930
rect 45442 8878 45444 8930
rect 44940 8372 44996 8382
rect 44940 8278 44996 8316
rect 45388 8370 45444 8878
rect 45388 8318 45390 8370
rect 45442 8318 45444 8370
rect 45388 8306 45444 8318
rect 45612 8372 45668 10220
rect 45164 8258 45220 8270
rect 45164 8206 45166 8258
rect 45218 8206 45220 8258
rect 44604 7474 44660 7486
rect 44604 7422 44606 7474
rect 44658 7422 44660 7474
rect 44492 7364 44548 7374
rect 44604 7364 44660 7422
rect 44492 7362 44660 7364
rect 44492 7310 44494 7362
rect 44546 7310 44660 7362
rect 44492 7308 44660 7310
rect 44492 7298 44548 7308
rect 43820 4174 43822 4226
rect 43874 4174 43876 4226
rect 34300 4162 34356 4172
rect 43820 4162 43876 4174
rect 44044 5906 44436 5908
rect 44044 5854 44382 5906
rect 44434 5854 44436 5906
rect 44044 5852 44436 5854
rect 44044 5234 44100 5852
rect 44380 5842 44436 5852
rect 44044 5182 44046 5234
rect 44098 5182 44100 5234
rect 44044 4340 44100 5182
rect 44604 5236 44660 7308
rect 45164 6692 45220 8206
rect 45612 8258 45668 8316
rect 45612 8206 45614 8258
rect 45666 8206 45668 8258
rect 45612 8194 45668 8206
rect 45724 8260 45780 8270
rect 45724 7700 45780 8204
rect 45836 8260 45892 8270
rect 46284 8260 46340 8270
rect 45836 8258 46340 8260
rect 45836 8206 45838 8258
rect 45890 8206 46286 8258
rect 46338 8206 46340 8258
rect 45836 8204 46340 8206
rect 45836 8194 45892 8204
rect 46284 8194 46340 8204
rect 46396 8260 46452 8270
rect 46396 8166 46452 8204
rect 46172 8036 46228 8046
rect 45836 7700 45892 7710
rect 45724 7698 45892 7700
rect 45724 7646 45838 7698
rect 45890 7646 45892 7698
rect 45724 7644 45892 7646
rect 45836 7634 45892 7644
rect 45052 6636 45164 6692
rect 45052 6132 45108 6636
rect 45164 6626 45220 6636
rect 45052 6018 45108 6076
rect 46172 6020 46228 7980
rect 46396 6692 46452 6702
rect 46508 6692 46564 15484
rect 46620 15204 46676 15242
rect 46620 15138 46676 15148
rect 46732 14532 46788 18508
rect 46956 17666 47012 19740
rect 47068 17778 47124 19966
rect 47292 20020 47348 20526
rect 47180 19236 47236 19246
rect 47180 19142 47236 19180
rect 47068 17726 47070 17778
rect 47122 17726 47124 17778
rect 47068 17714 47124 17726
rect 46956 17614 46958 17666
rect 47010 17614 47012 17666
rect 46956 17602 47012 17614
rect 47180 17668 47236 17678
rect 47180 17574 47236 17612
rect 47292 17444 47348 19964
rect 47516 20018 47572 21532
rect 47852 21474 47908 21756
rect 47852 21422 47854 21474
rect 47906 21422 47908 21474
rect 47852 20356 47908 21422
rect 47852 20300 48132 20356
rect 47964 20130 48020 20142
rect 47964 20078 47966 20130
rect 48018 20078 48020 20130
rect 47516 19966 47518 20018
rect 47570 19966 47572 20018
rect 47516 19796 47572 19966
rect 47740 20018 47796 20030
rect 47740 19966 47742 20018
rect 47794 19966 47796 20018
rect 47516 19730 47572 19740
rect 47628 19906 47684 19918
rect 47628 19854 47630 19906
rect 47682 19854 47684 19906
rect 47628 19460 47684 19854
rect 47628 19394 47684 19404
rect 47740 19124 47796 19966
rect 47964 20020 48020 20078
rect 47964 19954 48020 19964
rect 47852 19908 47908 19918
rect 47852 19346 47908 19852
rect 47852 19294 47854 19346
rect 47906 19294 47908 19346
rect 47852 19282 47908 19294
rect 47740 18340 47796 19068
rect 47964 18340 48020 18350
rect 47740 18338 48020 18340
rect 47740 18286 47966 18338
rect 48018 18286 48020 18338
rect 47740 18284 48020 18286
rect 47964 18274 48020 18284
rect 47852 18116 47908 18126
rect 47404 17444 47460 17454
rect 47292 17388 47404 17444
rect 47404 17350 47460 17388
rect 47740 15988 47796 15998
rect 47180 15876 47236 15886
rect 46844 15316 46900 15326
rect 46844 15222 46900 15260
rect 47068 15202 47124 15214
rect 47068 15150 47070 15202
rect 47122 15150 47124 15202
rect 47068 15148 47124 15150
rect 46956 15092 47124 15148
rect 46844 14532 46900 14542
rect 46732 14530 46900 14532
rect 46732 14478 46846 14530
rect 46898 14478 46900 14530
rect 46732 14476 46900 14478
rect 46844 14466 46900 14476
rect 46620 14418 46676 14430
rect 46620 14366 46622 14418
rect 46674 14366 46676 14418
rect 46620 14308 46676 14366
rect 46956 14308 47012 15092
rect 47180 14530 47236 15820
rect 47292 15540 47348 15550
rect 47292 15314 47348 15484
rect 47740 15538 47796 15932
rect 47852 15986 47908 18060
rect 47852 15934 47854 15986
rect 47906 15934 47908 15986
rect 47852 15922 47908 15934
rect 47740 15486 47742 15538
rect 47794 15486 47796 15538
rect 47740 15474 47796 15486
rect 47292 15262 47294 15314
rect 47346 15262 47348 15314
rect 47292 15250 47348 15262
rect 48076 15148 48132 20300
rect 48972 16994 49028 17006
rect 48972 16942 48974 16994
rect 49026 16942 49028 16994
rect 48972 15876 49028 16942
rect 48972 15810 49028 15820
rect 48972 15540 49028 15550
rect 48972 15314 49028 15484
rect 49084 15426 49140 21868
rect 49644 21812 49700 21822
rect 49644 21718 49700 21756
rect 49756 21700 49812 21710
rect 49756 21606 49812 21644
rect 50092 19794 50148 19806
rect 50092 19742 50094 19794
rect 50146 19742 50148 19794
rect 49980 19348 50036 19358
rect 49868 19346 50036 19348
rect 49868 19294 49982 19346
rect 50034 19294 50036 19346
rect 49868 19292 50036 19294
rect 49868 17668 49924 19292
rect 49980 19282 50036 19292
rect 50092 19236 50148 19742
rect 50092 19124 50148 19180
rect 49868 17602 49924 17612
rect 49980 19068 50148 19124
rect 49308 17556 49364 17566
rect 49308 16882 49364 17500
rect 49308 16830 49310 16882
rect 49362 16830 49364 16882
rect 49308 16210 49364 16830
rect 49308 16158 49310 16210
rect 49362 16158 49364 16210
rect 49308 16146 49364 16158
rect 49532 16098 49588 16110
rect 49532 16046 49534 16098
rect 49586 16046 49588 16098
rect 49084 15374 49086 15426
rect 49138 15374 49140 15426
rect 49084 15362 49140 15374
rect 49420 15876 49476 15886
rect 49420 15426 49476 15820
rect 49420 15374 49422 15426
rect 49474 15374 49476 15426
rect 49420 15362 49476 15374
rect 48972 15262 48974 15314
rect 49026 15262 49028 15314
rect 48972 15250 49028 15262
rect 49308 15202 49364 15214
rect 49308 15150 49310 15202
rect 49362 15150 49364 15202
rect 48076 15092 48468 15148
rect 47852 14532 47908 14542
rect 47180 14478 47182 14530
rect 47234 14478 47236 14530
rect 47180 14466 47236 14478
rect 47404 14530 47908 14532
rect 47404 14478 47854 14530
rect 47906 14478 47908 14530
rect 47404 14476 47908 14478
rect 46620 14252 47012 14308
rect 47068 14308 47124 14318
rect 47404 14308 47460 14476
rect 47068 14306 47460 14308
rect 47068 14254 47070 14306
rect 47122 14254 47460 14306
rect 47068 14252 47460 14254
rect 47516 14306 47572 14318
rect 47516 14254 47518 14306
rect 47570 14254 47572 14306
rect 46620 12964 46676 14252
rect 47068 14242 47124 14252
rect 47516 13860 47572 14254
rect 47628 14308 47684 14318
rect 47628 13970 47684 14252
rect 47628 13918 47630 13970
rect 47682 13918 47684 13970
rect 47628 13906 47684 13918
rect 47852 13970 47908 14476
rect 48076 14532 48132 14542
rect 48076 14438 48132 14476
rect 47852 13918 47854 13970
rect 47906 13918 47908 13970
rect 47852 13906 47908 13918
rect 48300 14420 48356 14430
rect 47292 13748 47348 13758
rect 47180 12964 47236 12974
rect 46620 12962 47236 12964
rect 46620 12910 47182 12962
rect 47234 12910 47236 12962
rect 46620 12908 47236 12910
rect 46732 11506 46788 12908
rect 47180 12898 47236 12908
rect 46732 11454 46734 11506
rect 46786 11454 46788 11506
rect 46732 11442 46788 11454
rect 46620 10724 46676 10734
rect 47180 10724 47236 10734
rect 47292 10724 47348 13692
rect 47516 13076 47572 13804
rect 47740 13634 47796 13646
rect 47740 13582 47742 13634
rect 47794 13582 47796 13634
rect 47740 13300 47796 13582
rect 47740 13244 48244 13300
rect 48188 13186 48244 13244
rect 48188 13134 48190 13186
rect 48242 13134 48244 13186
rect 48188 13122 48244 13134
rect 48076 13076 48132 13086
rect 47516 13074 48132 13076
rect 47516 13022 48078 13074
rect 48130 13022 48132 13074
rect 47516 13020 48132 13022
rect 48076 13010 48132 13020
rect 48300 12964 48356 14364
rect 48188 12908 48356 12964
rect 47516 12852 47572 12862
rect 47516 12758 47572 12796
rect 47852 12852 47908 12862
rect 48188 12852 48244 12908
rect 47852 12850 48244 12852
rect 47852 12798 47854 12850
rect 47906 12798 48244 12850
rect 47852 12796 48244 12798
rect 47404 12738 47460 12750
rect 47404 12686 47406 12738
rect 47458 12686 47460 12738
rect 47404 12404 47460 12686
rect 47852 12628 47908 12796
rect 47852 12562 47908 12572
rect 47404 12348 47796 12404
rect 47740 12290 47796 12348
rect 47740 12238 47742 12290
rect 47794 12238 47796 12290
rect 47740 12226 47796 12238
rect 47852 11954 47908 11966
rect 47852 11902 47854 11954
rect 47906 11902 47908 11954
rect 47852 11508 47908 11902
rect 47852 11442 47908 11452
rect 46676 10668 46788 10724
rect 46620 10658 46676 10668
rect 46620 8148 46676 8158
rect 46620 8054 46676 8092
rect 46732 6692 46788 10668
rect 47180 10722 47348 10724
rect 47180 10670 47182 10722
rect 47234 10670 47348 10722
rect 47180 10668 47348 10670
rect 48300 10724 48356 10734
rect 48412 10724 48468 15092
rect 49308 14756 49364 15150
rect 49308 14690 49364 14700
rect 49532 13300 49588 16046
rect 49980 15148 50036 19068
rect 50204 18564 50260 22428
rect 50764 22484 50820 22494
rect 50764 22482 51044 22484
rect 50764 22430 50766 22482
rect 50818 22430 51044 22482
rect 50764 22428 51044 22430
rect 50764 22418 50820 22428
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50988 21700 51044 22428
rect 51212 22482 51268 22988
rect 51212 22430 51214 22482
rect 51266 22430 51268 22482
rect 51212 22418 51268 22430
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50316 19906 50372 19918
rect 50316 19854 50318 19906
rect 50370 19854 50372 19906
rect 50316 19794 50372 19854
rect 50316 19742 50318 19794
rect 50370 19742 50372 19794
rect 50316 19730 50372 19742
rect 50428 19234 50484 19246
rect 50428 19182 50430 19234
rect 50482 19182 50484 19234
rect 50204 18508 50372 18564
rect 50092 15876 50148 15886
rect 50092 15426 50148 15820
rect 50092 15374 50094 15426
rect 50146 15374 50148 15426
rect 50092 15362 50148 15374
rect 50316 15428 50372 18508
rect 50428 18450 50484 19182
rect 50876 19124 50932 19134
rect 50764 19012 50820 19050
rect 50876 19030 50932 19068
rect 50764 18946 50820 18956
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50876 18564 50932 18574
rect 50988 18564 51044 21644
rect 52220 21474 52276 23212
rect 52220 21422 52222 21474
rect 52274 21422 52276 21474
rect 52220 21410 52276 21422
rect 51212 19906 51268 19918
rect 51212 19854 51214 19906
rect 51266 19854 51268 19906
rect 50876 18562 51044 18564
rect 50876 18510 50878 18562
rect 50930 18510 51044 18562
rect 50876 18508 51044 18510
rect 51100 19122 51156 19134
rect 51100 19070 51102 19122
rect 51154 19070 51156 19122
rect 51100 18564 51156 19070
rect 51212 19012 51268 19854
rect 51212 18946 51268 18956
rect 51436 19010 51492 19022
rect 51436 18958 51438 19010
rect 51490 18958 51492 19010
rect 50876 18498 50932 18508
rect 51100 18498 51156 18508
rect 50428 18398 50430 18450
rect 50482 18398 50484 18450
rect 50428 17666 50484 18398
rect 51324 18450 51380 18462
rect 51324 18398 51326 18450
rect 51378 18398 51380 18450
rect 51100 18338 51156 18350
rect 51100 18286 51102 18338
rect 51154 18286 51156 18338
rect 50652 18004 50708 18014
rect 50540 17948 50652 18004
rect 50540 17778 50596 17948
rect 50652 17938 50708 17948
rect 50540 17726 50542 17778
rect 50594 17726 50596 17778
rect 50540 17714 50596 17726
rect 50988 17780 51044 17790
rect 50428 17614 50430 17666
rect 50482 17614 50484 17666
rect 50428 17556 50484 17614
rect 50652 17668 50708 17678
rect 50652 17574 50708 17612
rect 50988 17666 51044 17724
rect 50988 17614 50990 17666
rect 51042 17614 51044 17666
rect 50988 17602 51044 17614
rect 50428 17490 50484 17500
rect 51100 17444 51156 18286
rect 51324 18228 51380 18398
rect 51324 18162 51380 18172
rect 51436 18004 51492 18958
rect 51548 19010 51604 19022
rect 51548 18958 51550 19010
rect 51602 18958 51604 19010
rect 51548 18452 51604 18958
rect 51548 18386 51604 18396
rect 51660 19010 51716 19022
rect 51660 18958 51662 19010
rect 51714 18958 51716 19010
rect 51436 17892 51492 17948
rect 51548 17892 51604 17902
rect 51436 17890 51604 17892
rect 51436 17838 51550 17890
rect 51602 17838 51604 17890
rect 51436 17836 51604 17838
rect 51548 17826 51604 17836
rect 51100 17378 51156 17388
rect 51324 17668 51380 17678
rect 51660 17668 51716 18958
rect 51884 19012 51940 19022
rect 51884 18918 51940 18956
rect 52780 19010 52836 19022
rect 52780 18958 52782 19010
rect 52834 18958 52836 19010
rect 52556 18564 52612 18574
rect 52780 18564 52836 18958
rect 52556 18562 52836 18564
rect 52556 18510 52558 18562
rect 52610 18510 52836 18562
rect 52556 18508 52836 18510
rect 52220 18452 52276 18462
rect 52220 18358 52276 18396
rect 52556 18340 52612 18508
rect 51324 17666 51716 17668
rect 51324 17614 51326 17666
rect 51378 17614 51716 17666
rect 51324 17612 51716 17614
rect 51772 18228 51828 18238
rect 52332 18228 52388 18238
rect 51324 17444 51380 17612
rect 51324 17378 51380 17388
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 51436 16884 51492 16894
rect 51212 16772 51268 16782
rect 51436 16772 51492 16828
rect 51100 16770 51492 16772
rect 51100 16718 51214 16770
rect 51266 16718 51492 16770
rect 51100 16716 51492 16718
rect 51660 16884 51716 16894
rect 50540 15988 50596 15998
rect 50540 15894 50596 15932
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50428 15428 50484 15438
rect 50316 15426 50484 15428
rect 50316 15374 50430 15426
rect 50482 15374 50484 15426
rect 50316 15372 50484 15374
rect 50428 15362 50484 15372
rect 50652 15314 50708 15326
rect 50652 15262 50654 15314
rect 50706 15262 50708 15314
rect 50204 15204 50260 15242
rect 49980 15092 50148 15148
rect 50204 15138 50260 15148
rect 49532 13234 49588 13244
rect 49868 12404 49924 12414
rect 49868 12178 49924 12348
rect 49868 12126 49870 12178
rect 49922 12126 49924 12178
rect 49868 12114 49924 12126
rect 50092 11732 50148 15092
rect 50652 15092 50708 15262
rect 50652 15026 50708 15036
rect 51100 14980 51156 16716
rect 51212 16706 51268 16716
rect 51660 16098 51716 16828
rect 51772 16772 51828 18172
rect 51884 18172 52332 18228
rect 51884 17890 51940 18172
rect 52332 18134 52388 18172
rect 52556 18004 52612 18284
rect 52332 17948 52612 18004
rect 52892 18450 52948 18462
rect 52892 18398 52894 18450
rect 52946 18398 52948 18450
rect 51884 17838 51886 17890
rect 51938 17838 51940 17890
rect 51884 17106 51940 17838
rect 52108 17892 52164 17902
rect 51884 17054 51886 17106
rect 51938 17054 51940 17106
rect 51884 17042 51940 17054
rect 51996 17108 52052 17118
rect 51772 16706 51828 16716
rect 51996 16770 52052 17052
rect 52108 17106 52164 17836
rect 52332 17444 52388 17948
rect 52780 17892 52836 17902
rect 52332 17378 52388 17388
rect 52444 17836 52780 17892
rect 52108 17054 52110 17106
rect 52162 17054 52164 17106
rect 52108 17042 52164 17054
rect 51996 16718 51998 16770
rect 52050 16718 52052 16770
rect 51996 16706 52052 16718
rect 52332 16772 52388 16782
rect 51660 16046 51662 16098
rect 51714 16046 51716 16098
rect 51660 16034 51716 16046
rect 52108 15876 52164 15886
rect 51996 15874 52164 15876
rect 51996 15822 52110 15874
rect 52162 15822 52164 15874
rect 51996 15820 52164 15822
rect 51772 15428 51828 15438
rect 51772 15314 51828 15372
rect 51772 15262 51774 15314
rect 51826 15262 51828 15314
rect 51772 15250 51828 15262
rect 51996 15314 52052 15820
rect 52108 15810 52164 15820
rect 51996 15262 51998 15314
rect 52050 15262 52052 15314
rect 51548 15204 51604 15242
rect 51548 15138 51604 15148
rect 51100 14914 51156 14924
rect 51212 15090 51268 15102
rect 51212 15038 51214 15090
rect 51266 15038 51268 15090
rect 50540 14756 50596 14766
rect 51212 14756 51268 15038
rect 51996 14980 52052 15262
rect 51996 14914 52052 14924
rect 52108 15540 52164 15550
rect 50428 14644 50484 14654
rect 50204 14532 50260 14542
rect 50204 14438 50260 14476
rect 50428 13972 50484 14588
rect 50540 14308 50596 14700
rect 50764 14700 51212 14756
rect 50764 14644 50820 14700
rect 51212 14690 51268 14700
rect 50764 14550 50820 14588
rect 51100 14532 51156 14542
rect 50540 14242 50596 14252
rect 50876 14530 51156 14532
rect 50876 14478 51102 14530
rect 51154 14478 51156 14530
rect 50876 14476 51156 14478
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50652 13972 50708 13982
rect 50428 13970 50708 13972
rect 50428 13918 50654 13970
rect 50706 13918 50708 13970
rect 50428 13916 50708 13918
rect 50652 13906 50708 13916
rect 50764 13972 50820 13982
rect 50876 13972 50932 14476
rect 51100 14466 51156 14476
rect 51212 14532 51268 14542
rect 51212 14438 51268 14476
rect 52108 14530 52164 15484
rect 52108 14478 52110 14530
rect 52162 14478 52164 14530
rect 51772 14420 51828 14430
rect 51660 14364 51772 14420
rect 50764 13970 50932 13972
rect 50764 13918 50766 13970
rect 50818 13918 50932 13970
rect 50764 13916 50932 13918
rect 50988 14308 51044 14318
rect 50764 13906 50820 13916
rect 50204 13748 50260 13758
rect 50204 13654 50260 13692
rect 50876 13748 50932 13758
rect 50988 13748 51044 14252
rect 51548 14308 51604 14318
rect 51548 14214 51604 14252
rect 50876 13746 51044 13748
rect 50876 13694 50878 13746
rect 50930 13694 51044 13746
rect 50876 13692 51044 13694
rect 50876 13682 50932 13692
rect 50316 13636 50372 13646
rect 48860 11508 48916 11518
rect 50092 11508 50148 11676
rect 48860 11414 48916 11452
rect 49644 11506 50148 11508
rect 49644 11454 50094 11506
rect 50146 11454 50148 11506
rect 49644 11452 50148 11454
rect 49644 11394 49700 11452
rect 50092 11442 50148 11452
rect 50204 12852 50260 12862
rect 49644 11342 49646 11394
rect 49698 11342 49700 11394
rect 49644 11330 49700 11342
rect 48356 10668 48468 10724
rect 50204 10834 50260 12796
rect 50316 12292 50372 13580
rect 50876 13524 50932 13534
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50316 12178 50372 12236
rect 50316 12126 50318 12178
rect 50370 12126 50372 12178
rect 50316 12114 50372 12126
rect 50652 12404 50708 12414
rect 50652 11506 50708 12348
rect 50652 11454 50654 11506
rect 50706 11454 50708 11506
rect 50652 11442 50708 11454
rect 50764 11844 50820 11854
rect 50764 11172 50820 11788
rect 50876 11396 50932 13468
rect 51100 12738 51156 12750
rect 51100 12686 51102 12738
rect 51154 12686 51156 12738
rect 50988 12290 51044 12302
rect 50988 12238 50990 12290
rect 51042 12238 51044 12290
rect 50988 11844 51044 12238
rect 51100 12180 51156 12686
rect 51436 12738 51492 12750
rect 51436 12686 51438 12738
rect 51490 12686 51492 12738
rect 51436 12404 51492 12686
rect 51436 12338 51492 12348
rect 51660 12402 51716 14364
rect 51772 14326 51828 14364
rect 51884 14306 51940 14318
rect 51884 14254 51886 14306
rect 51938 14254 51940 14306
rect 51884 13748 51940 14254
rect 51884 13682 51940 13692
rect 52108 13636 52164 14478
rect 52220 13636 52276 13646
rect 52108 13580 52220 13636
rect 52220 13570 52276 13580
rect 52332 12516 52388 16716
rect 52444 15538 52500 17836
rect 52780 17798 52836 17836
rect 52668 17666 52724 17678
rect 52668 17614 52670 17666
rect 52722 17614 52724 17666
rect 52556 17444 52612 17454
rect 52556 16884 52612 17388
rect 52668 17108 52724 17614
rect 52892 17556 52948 18398
rect 52892 17490 52948 17500
rect 53004 17332 53060 23492
rect 53340 23044 53396 24558
rect 53452 24052 53508 24062
rect 53508 23996 53732 24052
rect 53452 23986 53508 23996
rect 53452 23828 53508 23838
rect 53452 23734 53508 23772
rect 53340 22978 53396 22988
rect 53564 23042 53620 23996
rect 53676 23826 53732 23996
rect 53788 23940 53844 25454
rect 54124 24724 54180 24734
rect 53788 23938 54068 23940
rect 53788 23886 53790 23938
rect 53842 23886 54068 23938
rect 53788 23884 54068 23886
rect 53788 23874 53844 23884
rect 53676 23774 53678 23826
rect 53730 23774 53732 23826
rect 53676 23762 53732 23774
rect 54012 23266 54068 23884
rect 54124 23938 54180 24668
rect 54124 23886 54126 23938
rect 54178 23886 54180 23938
rect 54124 23874 54180 23886
rect 54460 23940 54516 23950
rect 54460 23846 54516 23884
rect 54236 23714 54292 23726
rect 54236 23662 54238 23714
rect 54290 23662 54292 23714
rect 54012 23214 54014 23266
rect 54066 23214 54068 23266
rect 54012 23202 54068 23214
rect 54124 23268 54180 23278
rect 54236 23268 54292 23662
rect 54180 23212 54292 23268
rect 54348 23268 54404 23278
rect 54348 23266 54964 23268
rect 54348 23214 54350 23266
rect 54402 23214 54964 23266
rect 54348 23212 54964 23214
rect 54124 23174 54180 23212
rect 54348 23202 54404 23212
rect 53564 22990 53566 23042
rect 53618 22990 53620 23042
rect 53564 22978 53620 22990
rect 54684 23044 54740 23054
rect 54740 22988 54852 23044
rect 54684 22950 54740 22988
rect 54572 22260 54628 22270
rect 54572 22166 54628 22204
rect 54684 22146 54740 22158
rect 54684 22094 54686 22146
rect 54738 22094 54740 22146
rect 54684 21812 54740 22094
rect 54348 21756 54740 21812
rect 54348 21698 54404 21756
rect 54348 21646 54350 21698
rect 54402 21646 54404 21698
rect 54348 21634 54404 21646
rect 54796 21588 54852 22988
rect 54908 22370 54964 23212
rect 54908 22318 54910 22370
rect 54962 22318 54964 22370
rect 54908 22306 54964 22318
rect 54796 21522 54852 21532
rect 53116 18450 53172 18462
rect 53116 18398 53118 18450
rect 53170 18398 53172 18450
rect 53116 18004 53172 18398
rect 53452 18452 53508 18462
rect 53228 18340 53284 18350
rect 53228 18246 53284 18284
rect 53116 17938 53172 17948
rect 53452 17668 53508 18396
rect 53564 18338 53620 18350
rect 53564 18286 53566 18338
rect 53618 18286 53620 18338
rect 53564 18228 53620 18286
rect 54460 18340 54516 18350
rect 54460 18246 54516 18284
rect 53564 18162 53620 18172
rect 53788 18226 53844 18238
rect 53788 18174 53790 18226
rect 53842 18174 53844 18226
rect 53788 18116 53844 18174
rect 53788 18050 53844 18060
rect 54124 18226 54180 18238
rect 54124 18174 54126 18226
rect 54178 18174 54180 18226
rect 54124 17892 54180 18174
rect 54572 18228 54628 18238
rect 54572 18134 54628 18172
rect 54124 17826 54180 17836
rect 54348 17778 54404 17790
rect 54348 17726 54350 17778
rect 54402 17726 54404 17778
rect 53564 17668 53620 17678
rect 54348 17668 54404 17726
rect 53452 17666 53844 17668
rect 53452 17614 53566 17666
rect 53618 17614 53844 17666
rect 53452 17612 53844 17614
rect 53564 17602 53620 17612
rect 53228 17556 53284 17566
rect 53340 17556 53396 17566
rect 53284 17554 53396 17556
rect 53284 17502 53342 17554
rect 53394 17502 53396 17554
rect 53284 17500 53396 17502
rect 53116 17444 53172 17454
rect 53116 17350 53172 17388
rect 52668 17042 52724 17052
rect 52780 17276 53060 17332
rect 52668 16884 52724 16894
rect 52556 16882 52724 16884
rect 52556 16830 52670 16882
rect 52722 16830 52724 16882
rect 52556 16828 52724 16830
rect 52668 16818 52724 16828
rect 52780 16660 52836 17276
rect 52892 16884 52948 16894
rect 52892 16790 52948 16828
rect 52780 16604 52948 16660
rect 52444 15486 52446 15538
rect 52498 15486 52500 15538
rect 52444 15428 52500 15486
rect 52444 15362 52500 15372
rect 52668 15314 52724 15326
rect 52668 15262 52670 15314
rect 52722 15262 52724 15314
rect 52556 15202 52612 15214
rect 52556 15150 52558 15202
rect 52610 15150 52612 15202
rect 52556 14756 52612 15150
rect 52668 15204 52724 15262
rect 52668 15138 52724 15148
rect 52668 14756 52724 14766
rect 52556 14754 52724 14756
rect 52556 14702 52670 14754
rect 52722 14702 52724 14754
rect 52556 14700 52724 14702
rect 52668 14690 52724 14700
rect 52780 14756 52836 14766
rect 52780 14662 52836 14700
rect 52780 13860 52836 13870
rect 52780 13766 52836 13804
rect 52668 13748 52724 13758
rect 52668 13654 52724 13692
rect 51660 12350 51662 12402
rect 51714 12350 51716 12402
rect 51660 12338 51716 12350
rect 52108 12460 52612 12516
rect 52108 12402 52164 12460
rect 52108 12350 52110 12402
rect 52162 12350 52164 12402
rect 52108 12338 52164 12350
rect 52220 12292 52276 12302
rect 52220 12198 52276 12236
rect 51324 12180 51380 12190
rect 51100 12178 51380 12180
rect 51100 12126 51326 12178
rect 51378 12126 51380 12178
rect 51100 12124 51380 12126
rect 50988 11778 51044 11788
rect 50988 11396 51044 11406
rect 50876 11394 51044 11396
rect 50876 11342 50990 11394
rect 51042 11342 51044 11394
rect 50876 11340 51044 11342
rect 50988 11330 51044 11340
rect 50764 11116 50932 11172
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50204 10782 50206 10834
rect 50258 10782 50260 10834
rect 46844 10610 46900 10622
rect 46844 10558 46846 10610
rect 46898 10558 46900 10610
rect 46844 10164 46900 10558
rect 46844 10098 46900 10108
rect 47180 9156 47236 10668
rect 48300 10658 48356 10668
rect 49868 10612 49924 10622
rect 49532 10500 49588 10510
rect 49868 10500 49924 10556
rect 47180 9090 47236 9100
rect 49420 10498 49924 10500
rect 49420 10446 49534 10498
rect 49586 10446 49924 10498
rect 49420 10444 49924 10446
rect 47516 8930 47572 8942
rect 47516 8878 47518 8930
rect 47570 8878 47572 8930
rect 47404 8372 47460 8382
rect 47404 8278 47460 8316
rect 47180 8258 47236 8270
rect 47180 8206 47182 8258
rect 47234 8206 47236 8258
rect 47180 8036 47236 8206
rect 47516 8260 47572 8878
rect 47516 8166 47572 8204
rect 48412 8258 48468 8270
rect 48412 8206 48414 8258
rect 48466 8206 48468 8258
rect 47852 8148 47908 8158
rect 47852 8054 47908 8092
rect 48188 8146 48244 8158
rect 48188 8094 48190 8146
rect 48242 8094 48244 8146
rect 47180 7812 47236 7980
rect 47180 7746 47236 7756
rect 46844 6692 46900 6702
rect 46396 6690 46508 6692
rect 46396 6638 46398 6690
rect 46450 6638 46508 6690
rect 46396 6636 46508 6638
rect 46396 6626 46452 6636
rect 46508 6598 46564 6636
rect 46620 6690 46900 6692
rect 46620 6638 46846 6690
rect 46898 6638 46900 6690
rect 46620 6636 46900 6638
rect 46620 6468 46676 6636
rect 46844 6626 46900 6636
rect 47292 6692 47348 6702
rect 46284 6412 46676 6468
rect 46284 6130 46340 6412
rect 46620 6356 46676 6412
rect 46620 6290 46676 6300
rect 46284 6078 46286 6130
rect 46338 6078 46340 6130
rect 46284 6066 46340 6078
rect 46732 6132 46788 6142
rect 46732 6038 46788 6076
rect 45052 5966 45054 6018
rect 45106 5966 45108 6018
rect 45052 5954 45108 5966
rect 46060 6018 46228 6020
rect 46060 5966 46174 6018
rect 46226 5966 46228 6018
rect 46060 5964 46228 5966
rect 45276 5906 45332 5918
rect 45276 5854 45278 5906
rect 45330 5854 45332 5906
rect 45164 5794 45220 5806
rect 45164 5742 45166 5794
rect 45218 5742 45220 5794
rect 44604 5170 44660 5180
rect 44940 5684 44996 5694
rect 44940 5234 44996 5628
rect 44940 5182 44942 5234
rect 44994 5182 44996 5234
rect 44940 5170 44996 5182
rect 44940 4452 44996 4462
rect 45164 4452 45220 5742
rect 45276 5684 45332 5854
rect 45612 5908 45668 5918
rect 45612 5906 45780 5908
rect 45612 5854 45614 5906
rect 45666 5854 45780 5906
rect 45612 5852 45780 5854
rect 45612 5842 45668 5852
rect 45276 5618 45332 5628
rect 45500 5236 45556 5246
rect 45500 5142 45556 5180
rect 45724 4900 45780 5852
rect 45836 5124 45892 5134
rect 46060 5124 46116 5964
rect 46172 5954 46228 5964
rect 46508 6020 46564 6030
rect 46508 5926 46564 5964
rect 46956 6018 47012 6030
rect 46956 5966 46958 6018
rect 47010 5966 47012 6018
rect 45836 5122 46116 5124
rect 45836 5070 45838 5122
rect 45890 5070 46116 5122
rect 45836 5068 46116 5070
rect 46508 5236 46564 5246
rect 46508 5122 46564 5180
rect 46508 5070 46510 5122
rect 46562 5070 46564 5122
rect 45836 5058 45892 5068
rect 46508 5058 46564 5070
rect 45948 4900 46004 4910
rect 45724 4898 46004 4900
rect 45724 4846 45950 4898
rect 46002 4846 46004 4898
rect 45724 4844 46004 4846
rect 45948 4834 46004 4844
rect 46060 4898 46116 4910
rect 46060 4846 46062 4898
rect 46114 4846 46116 4898
rect 44940 4450 45220 4452
rect 44940 4398 44942 4450
rect 44994 4398 45220 4450
rect 44940 4396 45220 4398
rect 44940 4386 44996 4396
rect 44156 4340 44212 4350
rect 44044 4338 44212 4340
rect 44044 4286 44158 4338
rect 44210 4286 44212 4338
rect 44044 4284 44212 4286
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 21532 3614 21534 3666
rect 21586 3614 21588 3666
rect 21532 3602 21588 3614
rect 43932 3668 43988 3678
rect 44044 3668 44100 4284
rect 44156 4274 44212 4284
rect 46060 4228 46116 4846
rect 46956 4564 47012 5966
rect 47068 6020 47124 6030
rect 47068 5926 47124 5964
rect 47292 6018 47348 6636
rect 48188 6468 48244 8094
rect 48188 6402 48244 6412
rect 48412 6690 48468 8206
rect 48636 8258 48692 8270
rect 48636 8206 48638 8258
rect 48690 8206 48692 8258
rect 48636 8148 48692 8206
rect 48860 8260 48916 8270
rect 48860 8166 48916 8204
rect 48524 8036 48580 8046
rect 48524 6804 48580 7980
rect 48636 7364 48692 8092
rect 49308 8034 49364 8046
rect 49308 7982 49310 8034
rect 49362 7982 49364 8034
rect 49308 7924 49364 7982
rect 49308 7858 49364 7868
rect 48636 7298 48692 7308
rect 49420 7252 49476 10444
rect 49532 10434 49588 10444
rect 50204 10052 50260 10782
rect 50876 10724 50932 11116
rect 50876 10658 50932 10668
rect 51100 11170 51156 11182
rect 51100 11118 51102 11170
rect 51154 11118 51156 11170
rect 50652 10500 50708 10510
rect 51100 10500 51156 11118
rect 51212 10612 51268 12124
rect 51324 12114 51380 12124
rect 51884 12178 51940 12190
rect 51884 12126 51886 12178
rect 51938 12126 51940 12178
rect 51660 11508 51716 11518
rect 51660 11414 51716 11452
rect 51884 11394 51940 12126
rect 52556 11508 52612 12460
rect 52668 12292 52724 12302
rect 52668 12198 52724 12236
rect 52668 11508 52724 11518
rect 52556 11506 52724 11508
rect 52556 11454 52670 11506
rect 52722 11454 52724 11506
rect 52556 11452 52724 11454
rect 52668 11442 52724 11452
rect 52108 11396 52164 11406
rect 51884 11342 51886 11394
rect 51938 11342 51940 11394
rect 51884 11330 51940 11342
rect 51996 11340 52108 11396
rect 51324 11284 51380 11294
rect 51548 11284 51604 11294
rect 51324 11282 51604 11284
rect 51324 11230 51326 11282
rect 51378 11230 51550 11282
rect 51602 11230 51604 11282
rect 51324 11228 51604 11230
rect 51324 11218 51380 11228
rect 51548 11218 51604 11228
rect 51996 10834 52052 11340
rect 52108 11302 52164 11340
rect 52892 11396 52948 16604
rect 53228 14420 53284 17500
rect 53340 17490 53396 17500
rect 53452 17442 53508 17454
rect 53452 17390 53454 17442
rect 53506 17390 53508 17442
rect 53452 17220 53508 17390
rect 53452 17154 53508 17164
rect 53564 17332 53620 17342
rect 53564 16882 53620 17276
rect 53564 16830 53566 16882
rect 53618 16830 53620 16882
rect 53564 16818 53620 16830
rect 53788 16884 53844 17612
rect 54348 17602 54404 17612
rect 55020 17556 55076 27244
rect 55356 27074 55412 28028
rect 56588 28082 56644 28476
rect 56588 28030 56590 28082
rect 56642 28030 56644 28082
rect 56588 28018 56644 28030
rect 57372 28082 57428 29596
rect 57372 28030 57374 28082
rect 57426 28030 57428 28082
rect 57372 28018 57428 28030
rect 55468 27972 55524 27982
rect 56924 27972 56980 27982
rect 55468 27878 55524 27916
rect 56700 27970 56980 27972
rect 56700 27918 56926 27970
rect 56978 27918 56980 27970
rect 56700 27916 56980 27918
rect 56700 27412 56756 27916
rect 56924 27906 56980 27916
rect 57260 27972 57316 27982
rect 57260 27878 57316 27916
rect 57596 27860 57652 29932
rect 57820 29652 57876 29662
rect 57932 29652 57988 31052
rect 58156 31042 58212 31052
rect 57820 29650 57988 29652
rect 57820 29598 57822 29650
rect 57874 29598 57988 29650
rect 57820 29596 57988 29598
rect 58156 30322 58212 30334
rect 58156 30270 58158 30322
rect 58210 30270 58212 30322
rect 58156 29652 58212 30270
rect 57820 29586 57876 29596
rect 58156 29586 58212 29596
rect 58156 29316 58212 29326
rect 58044 29314 58212 29316
rect 58044 29262 58158 29314
rect 58210 29262 58212 29314
rect 58044 29260 58212 29262
rect 58044 28756 58100 29260
rect 58156 29250 58212 29260
rect 57932 27972 57988 27982
rect 57932 27878 57988 27916
rect 57820 27860 57876 27870
rect 57596 27858 57876 27860
rect 57596 27806 57822 27858
rect 57874 27806 57876 27858
rect 57596 27804 57876 27806
rect 55356 27022 55358 27074
rect 55410 27022 55412 27074
rect 55356 27010 55412 27022
rect 56588 27356 56756 27412
rect 56812 27748 56868 27758
rect 56028 26962 56084 26974
rect 56028 26910 56030 26962
rect 56082 26910 56084 26962
rect 56028 26516 56084 26910
rect 56028 26450 56084 26460
rect 56588 26292 56644 27356
rect 56476 26290 56644 26292
rect 56476 26238 56590 26290
rect 56642 26238 56644 26290
rect 56476 26236 56644 26238
rect 56364 25282 56420 25294
rect 56364 25230 56366 25282
rect 56418 25230 56420 25282
rect 56364 24724 56420 25230
rect 56476 25172 56532 26236
rect 56588 26226 56644 26236
rect 56700 27188 56756 27198
rect 56700 26068 56756 27132
rect 56588 26012 56756 26068
rect 56588 25394 56644 26012
rect 56588 25342 56590 25394
rect 56642 25342 56644 25394
rect 56588 25330 56644 25342
rect 56700 25508 56756 25518
rect 56812 25508 56868 27692
rect 56924 27636 56980 27646
rect 56924 26290 56980 27580
rect 57372 27634 57428 27646
rect 57372 27582 57374 27634
rect 57426 27582 57428 27634
rect 57036 26516 57092 26526
rect 57036 26422 57092 26460
rect 56924 26238 56926 26290
rect 56978 26238 56980 26290
rect 56924 26226 56980 26238
rect 57260 26292 57316 26302
rect 57372 26292 57428 27582
rect 57820 26908 57876 27804
rect 57932 27636 57988 27646
rect 57932 27542 57988 27580
rect 57820 26852 57988 26908
rect 57260 26290 57428 26292
rect 57260 26238 57262 26290
rect 57314 26238 57428 26290
rect 57260 26236 57428 26238
rect 57260 26226 57316 26236
rect 56700 25506 56868 25508
rect 56700 25454 56702 25506
rect 56754 25454 56868 25506
rect 56700 25452 56868 25454
rect 56476 25116 56644 25172
rect 56476 24724 56532 24734
rect 56364 24722 56532 24724
rect 56364 24670 56478 24722
rect 56530 24670 56532 24722
rect 56364 24668 56532 24670
rect 56476 24658 56532 24668
rect 56588 24724 56644 25116
rect 56588 24658 56644 24668
rect 56700 24164 56756 25452
rect 57596 25284 57652 25294
rect 57596 25190 57652 25228
rect 57820 25282 57876 25294
rect 57820 25230 57822 25282
rect 57874 25230 57876 25282
rect 56812 24948 56868 24958
rect 56812 24946 57316 24948
rect 56812 24894 56814 24946
rect 56866 24894 57316 24946
rect 56812 24892 57316 24894
rect 56812 24882 56868 24892
rect 56924 24722 56980 24734
rect 56924 24670 56926 24722
rect 56978 24670 56980 24722
rect 56700 24108 56868 24164
rect 55132 24050 55188 24062
rect 55132 23998 55134 24050
rect 55186 23998 55188 24050
rect 55132 23380 55188 23998
rect 55132 23314 55188 23324
rect 56700 23380 56756 23390
rect 56588 23268 56644 23278
rect 56588 23174 56644 23212
rect 55132 22258 55188 22270
rect 55132 22206 55134 22258
rect 55186 22206 55188 22258
rect 55132 22036 55188 22206
rect 56700 22258 56756 23324
rect 56812 22372 56868 24108
rect 56924 23378 56980 24670
rect 56924 23326 56926 23378
rect 56978 23326 56980 23378
rect 56924 23314 56980 23326
rect 57148 24724 57204 24734
rect 56812 22278 56868 22316
rect 56700 22206 56702 22258
rect 56754 22206 56756 22258
rect 56700 22194 56756 22206
rect 57036 22260 57092 22270
rect 57036 22166 57092 22204
rect 55132 21970 55188 21980
rect 56476 22146 56532 22158
rect 56476 22094 56478 22146
rect 56530 22094 56532 22146
rect 55132 21588 55188 21598
rect 55580 21588 55636 21598
rect 55188 21586 55636 21588
rect 55188 21534 55582 21586
rect 55634 21534 55636 21586
rect 55188 21532 55636 21534
rect 55132 21494 55188 21532
rect 55244 20802 55300 21532
rect 55580 21522 55636 21532
rect 56476 21586 56532 22094
rect 56924 22148 56980 22158
rect 56924 21698 56980 22092
rect 56924 21646 56926 21698
rect 56978 21646 56980 21698
rect 56924 21634 56980 21646
rect 57148 22036 57204 24668
rect 57260 24050 57316 24892
rect 57820 24834 57876 25230
rect 57820 24782 57822 24834
rect 57874 24782 57876 24834
rect 57820 24770 57876 24782
rect 57484 24612 57540 24622
rect 57484 24518 57540 24556
rect 57260 23998 57262 24050
rect 57314 23998 57316 24050
rect 57260 23986 57316 23998
rect 57932 23268 57988 26852
rect 57372 22372 57428 22382
rect 57372 22278 57428 22316
rect 57932 22370 57988 23212
rect 58044 26180 58100 28700
rect 58156 27972 58212 27982
rect 58156 27188 58212 27916
rect 58156 27094 58212 27132
rect 58156 26180 58212 26190
rect 58044 26178 58212 26180
rect 58044 26126 58158 26178
rect 58210 26126 58212 26178
rect 58044 26124 58212 26126
rect 58044 23938 58100 26124
rect 58156 26114 58212 26124
rect 58268 25620 58324 38332
rect 58268 25554 58324 25564
rect 58156 25394 58212 25406
rect 58156 25342 58158 25394
rect 58210 25342 58212 25394
rect 58156 25284 58212 25342
rect 58156 24500 58212 25228
rect 58156 24434 58212 24444
rect 58044 23886 58046 23938
rect 58098 23886 58100 23938
rect 58044 23044 58100 23886
rect 58156 23044 58212 23054
rect 58044 23042 58324 23044
rect 58044 22990 58158 23042
rect 58210 22990 58324 23042
rect 58044 22988 58324 22990
rect 58156 22978 58212 22988
rect 57932 22318 57934 22370
rect 57986 22318 57988 22370
rect 57932 22306 57988 22318
rect 57148 21698 57204 21980
rect 57260 22146 57316 22158
rect 57260 22094 57262 22146
rect 57314 22094 57316 22146
rect 57260 21924 57316 22094
rect 57596 22148 57652 22158
rect 57596 22054 57652 22092
rect 57820 22146 57876 22158
rect 57820 22094 57822 22146
rect 57874 22094 57876 22146
rect 57820 21924 57876 22094
rect 57260 21868 57876 21924
rect 57148 21646 57150 21698
rect 57202 21646 57204 21698
rect 57148 21634 57204 21646
rect 56476 21534 56478 21586
rect 56530 21534 56532 21586
rect 56476 21522 56532 21534
rect 56700 21476 56756 21486
rect 56588 21474 56756 21476
rect 56588 21422 56702 21474
rect 56754 21422 56756 21474
rect 56588 21420 56756 21422
rect 56588 21028 56644 21420
rect 56700 21410 56756 21420
rect 56028 20972 56644 21028
rect 56028 20914 56084 20972
rect 56028 20862 56030 20914
rect 56082 20862 56084 20914
rect 56028 20850 56084 20862
rect 57820 20916 57876 21868
rect 58156 20916 58212 20926
rect 57820 20914 58212 20916
rect 57820 20862 58158 20914
rect 58210 20862 58212 20914
rect 57820 20860 58212 20862
rect 58156 20850 58212 20860
rect 55244 20750 55246 20802
rect 55298 20750 55300 20802
rect 55244 20738 55300 20750
rect 58156 20244 58212 20254
rect 58268 20244 58324 22988
rect 58156 20242 58324 20244
rect 58156 20190 58158 20242
rect 58210 20190 58324 20242
rect 58156 20188 58324 20190
rect 58156 20178 58212 20188
rect 55020 17490 55076 17500
rect 55132 18338 55188 18350
rect 55132 18286 55134 18338
rect 55186 18286 55188 18338
rect 55132 17220 55188 18286
rect 55132 17154 55188 17164
rect 55244 18226 55300 18238
rect 55244 18174 55246 18226
rect 55298 18174 55300 18226
rect 53340 16772 53396 16782
rect 53340 16678 53396 16716
rect 53788 16770 53844 16828
rect 55132 16884 55188 16894
rect 53788 16718 53790 16770
rect 53842 16718 53844 16770
rect 53788 16706 53844 16718
rect 54012 16770 54068 16782
rect 54012 16718 54014 16770
rect 54066 16718 54068 16770
rect 53564 15092 53620 15102
rect 53564 14530 53620 15036
rect 54012 15092 54068 16718
rect 55132 16212 55188 16828
rect 55244 16772 55300 18174
rect 56476 18228 56532 18238
rect 56476 17778 56532 18172
rect 56476 17726 56478 17778
rect 56530 17726 56532 17778
rect 56476 17714 56532 17726
rect 57260 17668 57316 17678
rect 57260 17666 57540 17668
rect 57260 17614 57262 17666
rect 57314 17614 57540 17666
rect 57260 17612 57540 17614
rect 57260 17602 57316 17612
rect 57484 17108 57540 17612
rect 57820 17556 57876 17566
rect 57820 17462 57876 17500
rect 58156 17556 58212 17566
rect 58212 17500 58324 17556
rect 58156 17462 58212 17500
rect 57484 17106 58100 17108
rect 57484 17054 57486 17106
rect 57538 17054 58100 17106
rect 57484 17052 58100 17054
rect 57484 17042 57540 17052
rect 55244 16706 55300 16716
rect 57036 16996 57092 17006
rect 55244 16212 55300 16222
rect 55132 16210 55300 16212
rect 55132 16158 55246 16210
rect 55298 16158 55300 16210
rect 55132 16156 55300 16158
rect 55244 16146 55300 16156
rect 54012 15026 54068 15036
rect 54460 15092 54516 15102
rect 53676 14644 53732 14654
rect 54012 14644 54068 14654
rect 53676 14642 54068 14644
rect 53676 14590 53678 14642
rect 53730 14590 54014 14642
rect 54066 14590 54068 14642
rect 53676 14588 54068 14590
rect 53676 14578 53732 14588
rect 54012 14578 54068 14588
rect 54460 14642 54516 15036
rect 54460 14590 54462 14642
rect 54514 14590 54516 14642
rect 54460 14578 54516 14590
rect 53564 14478 53566 14530
rect 53618 14478 53620 14530
rect 53564 14466 53620 14478
rect 53340 14420 53396 14430
rect 53228 14364 53340 14420
rect 53340 14326 53396 14364
rect 54124 14420 54180 14430
rect 54124 14326 54180 14364
rect 56588 14420 56644 14430
rect 56588 14326 56644 14364
rect 53116 14308 53172 14318
rect 53116 14214 53172 14252
rect 55244 13860 55300 13870
rect 55244 13766 55300 13804
rect 55916 13746 55972 13758
rect 55916 13694 55918 13746
rect 55970 13694 55972 13746
rect 53116 13636 53172 13646
rect 53116 13542 53172 13580
rect 54460 13636 54516 13646
rect 53004 12740 53060 12750
rect 53060 12684 53396 12740
rect 53004 12646 53060 12684
rect 53340 12178 53396 12684
rect 53340 12126 53342 12178
rect 53394 12126 53396 12178
rect 53340 12114 53396 12126
rect 54460 12066 54516 13580
rect 55916 13636 55972 13694
rect 55916 13570 55972 13580
rect 56700 13636 56756 13646
rect 56700 13542 56756 13580
rect 54460 12014 54462 12066
rect 54514 12014 54516 12066
rect 54460 11732 54516 12014
rect 54460 11666 54516 11676
rect 55580 11732 55636 11742
rect 57036 11732 57092 16940
rect 57372 16772 57428 16782
rect 57372 16210 57428 16716
rect 57372 16158 57374 16210
rect 57426 16158 57428 16210
rect 57372 16146 57428 16158
rect 58044 16098 58100 17052
rect 58268 17106 58324 17500
rect 58268 17054 58270 17106
rect 58322 17054 58324 17106
rect 58268 17042 58324 17054
rect 58044 16046 58046 16098
rect 58098 16046 58100 16098
rect 58044 15540 58100 16046
rect 58156 15540 58212 15550
rect 58044 15538 58212 15540
rect 58044 15486 58158 15538
rect 58210 15486 58212 15538
rect 58044 15484 58212 15486
rect 57260 14530 57316 14542
rect 57260 14478 57262 14530
rect 57314 14478 57316 14530
rect 57260 14420 57316 14478
rect 57260 13636 57316 14364
rect 57820 14420 57876 14430
rect 58156 14420 58212 15484
rect 57876 14364 58212 14420
rect 57820 14326 57876 14364
rect 57260 13570 57316 13580
rect 57036 11676 57316 11732
rect 54796 11508 54852 11518
rect 54796 11414 54852 11452
rect 52892 11330 52948 11340
rect 55580 11394 55636 11676
rect 57260 11618 57316 11676
rect 57260 11566 57262 11618
rect 57314 11566 57316 11618
rect 57260 11554 57316 11566
rect 55580 11342 55582 11394
rect 55634 11342 55636 11394
rect 51996 10782 51998 10834
rect 52050 10782 52052 10834
rect 51324 10724 51380 10734
rect 51324 10630 51380 10668
rect 51436 10724 51492 10734
rect 51436 10722 51604 10724
rect 51436 10670 51438 10722
rect 51490 10670 51604 10722
rect 51436 10668 51604 10670
rect 51436 10658 51492 10668
rect 51212 10546 51268 10556
rect 50708 10444 51156 10500
rect 50652 10406 50708 10444
rect 50204 9986 50260 9996
rect 50764 9828 50820 9838
rect 50316 9826 50820 9828
rect 50316 9774 50766 9826
rect 50818 9774 50820 9826
rect 50316 9772 50820 9774
rect 50204 9268 50260 9278
rect 50316 9268 50372 9772
rect 50764 9762 50820 9772
rect 50876 9714 50932 10444
rect 50876 9662 50878 9714
rect 50930 9662 50932 9714
rect 50428 9604 50484 9614
rect 50876 9604 50932 9662
rect 50428 9602 50932 9604
rect 50428 9550 50430 9602
rect 50482 9550 50932 9602
rect 50428 9548 50932 9550
rect 50988 10052 51044 10062
rect 50428 9538 50484 9548
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50204 9266 50596 9268
rect 50204 9214 50206 9266
rect 50258 9214 50596 9266
rect 50204 9212 50596 9214
rect 50204 9202 50260 9212
rect 49980 9156 50036 9166
rect 49980 8932 50036 9100
rect 50428 9042 50484 9054
rect 50428 8990 50430 9042
rect 50482 8990 50484 9042
rect 49980 8876 50260 8932
rect 49532 8258 49588 8270
rect 49532 8206 49534 8258
rect 49586 8206 49588 8258
rect 49532 8036 49588 8206
rect 49868 8148 49924 8158
rect 49868 8054 49924 8092
rect 49532 7970 49588 7980
rect 49644 7700 49700 7710
rect 49420 7186 49476 7196
rect 49532 7698 49700 7700
rect 49532 7646 49646 7698
rect 49698 7646 49700 7698
rect 49532 7644 49700 7646
rect 48748 6804 48804 6814
rect 48524 6748 48692 6804
rect 48412 6638 48414 6690
rect 48466 6638 48468 6690
rect 48412 6132 48468 6638
rect 48412 6066 48468 6076
rect 48524 6578 48580 6590
rect 48524 6526 48526 6578
rect 48578 6526 48580 6578
rect 47292 5966 47294 6018
rect 47346 5966 47348 6018
rect 47292 5954 47348 5966
rect 47516 5796 47572 5806
rect 47516 5794 47796 5796
rect 47516 5742 47518 5794
rect 47570 5742 47796 5794
rect 47516 5740 47796 5742
rect 47516 5730 47572 5740
rect 47740 5234 47796 5740
rect 47740 5182 47742 5234
rect 47794 5182 47796 5234
rect 47740 5170 47796 5182
rect 47068 5124 47124 5134
rect 47068 5030 47124 5068
rect 46956 4498 47012 4508
rect 46060 4162 46116 4172
rect 47068 4228 47124 4238
rect 47068 4134 47124 4172
rect 48524 4228 48580 6526
rect 48636 6580 48692 6748
rect 48748 6710 48804 6748
rect 49532 6692 49588 7644
rect 49644 7634 49700 7644
rect 49756 7700 49812 7710
rect 49756 7698 50036 7700
rect 49756 7646 49758 7698
rect 49810 7646 50036 7698
rect 49756 7644 50036 7646
rect 49756 7634 49812 7644
rect 49868 7476 49924 7486
rect 49868 7382 49924 7420
rect 49980 7252 50036 7644
rect 50204 7474 50260 8876
rect 50204 7422 50206 7474
rect 50258 7422 50260 7474
rect 50204 7410 50260 7422
rect 50316 8930 50372 8942
rect 50316 8878 50318 8930
rect 50370 8878 50372 8930
rect 50316 7476 50372 8878
rect 50428 8484 50484 8990
rect 50428 8418 50484 8428
rect 50428 8260 50484 8270
rect 50428 8166 50484 8204
rect 50540 8260 50596 9212
rect 50988 8428 51044 9996
rect 51548 9940 51604 10668
rect 51660 10612 51716 10622
rect 51660 10610 51828 10612
rect 51660 10558 51662 10610
rect 51714 10558 51828 10610
rect 51660 10556 51828 10558
rect 51660 10546 51716 10556
rect 51100 9828 51156 9838
rect 51436 9828 51492 9838
rect 51100 9826 51492 9828
rect 51100 9774 51102 9826
rect 51154 9774 51438 9826
rect 51490 9774 51492 9826
rect 51100 9772 51492 9774
rect 51100 9762 51156 9772
rect 51436 9762 51492 9772
rect 51324 9268 51380 9278
rect 51324 9174 51380 9212
rect 51548 8428 51604 9884
rect 51772 9826 51828 10556
rect 51772 9774 51774 9826
rect 51826 9774 51828 9826
rect 51772 9762 51828 9774
rect 51996 10388 52052 10782
rect 52444 10724 52500 10734
rect 52444 10630 52500 10668
rect 51996 9826 52052 10332
rect 52668 9940 52724 9950
rect 52668 9846 52724 9884
rect 51996 9774 51998 9826
rect 52050 9774 52052 9826
rect 51660 9716 51716 9726
rect 51660 9622 51716 9660
rect 51996 9268 52052 9774
rect 55580 9826 55636 11342
rect 57372 11284 57428 11294
rect 57820 11284 57876 11294
rect 57372 11282 57876 11284
rect 57372 11230 57374 11282
rect 57426 11230 57822 11282
rect 57874 11230 57876 11282
rect 57372 11228 57876 11230
rect 57372 11218 57428 11228
rect 57820 11218 57876 11228
rect 58156 11282 58212 11294
rect 58156 11230 58158 11282
rect 58210 11230 58212 11282
rect 55580 9774 55582 9826
rect 55634 9774 55636 9826
rect 54796 9716 54852 9726
rect 54796 9622 54852 9660
rect 55580 9604 55636 9774
rect 56028 11170 56084 11182
rect 56028 11118 56030 11170
rect 56082 11118 56084 11170
rect 56028 9604 56084 11118
rect 58156 10612 58212 11230
rect 58156 10518 58212 10556
rect 55580 9602 56084 9604
rect 55580 9550 56030 9602
rect 56082 9550 56084 9602
rect 55580 9548 56084 9550
rect 51996 9202 52052 9212
rect 50988 8372 51156 8428
rect 50988 8260 51044 8270
rect 50540 8258 51044 8260
rect 50540 8206 50990 8258
rect 51042 8206 51044 8258
rect 50540 8204 51044 8206
rect 50540 8034 50596 8204
rect 50988 8194 51044 8204
rect 50540 7982 50542 8034
rect 50594 7982 50596 8034
rect 50540 7970 50596 7982
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50652 7588 50708 7598
rect 50540 7476 50596 7486
rect 50316 7474 50596 7476
rect 50316 7422 50542 7474
rect 50594 7422 50596 7474
rect 50316 7420 50596 7422
rect 50540 7410 50596 7420
rect 50652 7474 50708 7532
rect 50652 7422 50654 7474
rect 50706 7422 50708 7474
rect 50652 7252 50708 7422
rect 50876 7586 50932 7598
rect 50876 7534 50878 7586
rect 50930 7534 50932 7586
rect 50876 7364 50932 7534
rect 49980 7196 50372 7252
rect 50316 6914 50372 7196
rect 50652 7186 50708 7196
rect 50764 7308 50876 7364
rect 50316 6862 50318 6914
rect 50370 6862 50372 6914
rect 50316 6850 50372 6862
rect 49980 6804 50036 6814
rect 49980 6710 50036 6748
rect 50428 6802 50484 6814
rect 50428 6750 50430 6802
rect 50482 6750 50484 6802
rect 49756 6692 49812 6702
rect 49532 6636 49756 6692
rect 49756 6598 49812 6636
rect 48860 6580 48916 6590
rect 48636 6578 48916 6580
rect 48636 6526 48862 6578
rect 48914 6526 48916 6578
rect 48636 6524 48916 6526
rect 48860 6514 48916 6524
rect 49420 6580 49476 6590
rect 49420 6486 49476 6524
rect 50428 6580 50484 6750
rect 50428 6514 50484 6524
rect 50764 6578 50820 7308
rect 50876 7298 50932 7308
rect 51100 7588 51156 8372
rect 51212 8372 51268 8382
rect 51212 8278 51268 8316
rect 51324 8372 51604 8428
rect 51324 8260 51380 8372
rect 51324 8194 51380 8204
rect 51548 8034 51604 8046
rect 51548 7982 51550 8034
rect 51602 7982 51604 8034
rect 51212 7588 51268 7598
rect 51100 7586 51268 7588
rect 51100 7534 51214 7586
rect 51266 7534 51268 7586
rect 51100 7532 51268 7534
rect 50988 6692 51044 6702
rect 51100 6692 51156 7532
rect 51212 7522 51268 7532
rect 51548 7588 51604 7982
rect 51548 7522 51604 7532
rect 51436 7476 51492 7486
rect 51436 6804 51492 7420
rect 51548 7364 51604 7374
rect 51548 7270 51604 7308
rect 52444 7364 52500 7374
rect 52444 7270 52500 7308
rect 52556 7250 52612 7262
rect 52556 7198 52558 7250
rect 52610 7198 52612 7250
rect 51548 6804 51604 6814
rect 51436 6748 51548 6804
rect 51548 6738 51604 6748
rect 50988 6690 51156 6692
rect 50988 6638 50990 6690
rect 51042 6638 51156 6690
rect 50988 6636 51156 6638
rect 52556 6692 52612 7198
rect 52668 6804 52724 6814
rect 52668 6710 52724 6748
rect 50988 6626 51044 6636
rect 52556 6626 52612 6636
rect 54796 6692 54852 6702
rect 54796 6598 54852 6636
rect 55468 6692 55524 6702
rect 56028 6692 56084 9548
rect 55468 6690 56084 6692
rect 55468 6638 55470 6690
rect 55522 6638 56030 6690
rect 56082 6638 56084 6690
rect 55468 6636 56084 6638
rect 50764 6526 50766 6578
rect 50818 6526 50820 6578
rect 50764 6514 50820 6526
rect 51212 6578 51268 6590
rect 51212 6526 51214 6578
rect 51266 6526 51268 6578
rect 51100 6466 51156 6478
rect 51100 6414 51102 6466
rect 51154 6414 51156 6466
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50428 6132 50484 6142
rect 49868 5908 49924 5918
rect 48860 5236 48916 5246
rect 48748 4564 48804 4574
rect 48748 4470 48804 4508
rect 48860 4450 48916 5180
rect 49868 5236 49924 5852
rect 49868 5142 49924 5180
rect 50316 5124 50372 5134
rect 50316 5030 50372 5068
rect 48860 4398 48862 4450
rect 48914 4398 48916 4450
rect 48860 4386 48916 4398
rect 50428 4228 50484 6076
rect 51100 5236 51156 6414
rect 51212 6132 51268 6526
rect 51212 6066 51268 6076
rect 54012 6468 54068 6478
rect 51212 5236 51268 5246
rect 51100 5234 51268 5236
rect 51100 5182 51214 5234
rect 51266 5182 51268 5234
rect 51100 5180 51268 5182
rect 51212 5170 51268 5180
rect 53340 5012 53396 5022
rect 51324 4900 51380 4910
rect 51324 4806 51380 4844
rect 52668 4900 52724 4910
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 52668 4450 52724 4844
rect 52668 4398 52670 4450
rect 52722 4398 52724 4450
rect 52668 4386 52724 4398
rect 53340 4564 53396 4956
rect 53900 4564 53956 4574
rect 53340 4562 53956 4564
rect 53340 4510 53902 4562
rect 53954 4510 53956 4562
rect 53340 4508 53956 4510
rect 53340 4338 53396 4508
rect 53900 4498 53956 4508
rect 53340 4286 53342 4338
rect 53394 4286 53396 4338
rect 53340 4274 53396 4286
rect 54012 4340 54068 6412
rect 55468 5012 55524 6636
rect 56028 6626 56084 6636
rect 55468 4946 55524 4956
rect 54012 4274 54068 4284
rect 57596 4340 57652 4350
rect 57596 4246 57652 4284
rect 58156 4338 58212 4350
rect 58156 4286 58158 4338
rect 58210 4286 58212 4338
rect 50540 4228 50596 4238
rect 50428 4226 50596 4228
rect 50428 4174 50542 4226
rect 50594 4174 50596 4226
rect 50428 4172 50596 4174
rect 48524 4162 48580 4172
rect 50540 4162 50596 4172
rect 57372 4228 57428 4238
rect 57372 4134 57428 4172
rect 58156 4228 58212 4286
rect 43932 3666 44100 3668
rect 43932 3614 43934 3666
rect 43986 3614 44100 3666
rect 43932 3612 44100 3614
rect 58156 3668 58212 4172
rect 43932 3602 43988 3612
rect 58156 3602 58212 3612
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
<< via2 >>
rect 4732 66780 4788 66836
rect 5516 66780 5572 66836
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 5740 64706 5796 64708
rect 5740 64654 5742 64706
rect 5742 64654 5794 64706
rect 5794 64654 5796 64706
rect 5740 64652 5796 64654
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 1708 58322 1764 58324
rect 1708 58270 1710 58322
rect 1710 58270 1762 58322
rect 1762 58270 1764 58322
rect 1708 58268 1764 58270
rect 1820 58604 1876 58660
rect 5628 60674 5684 60676
rect 5628 60622 5630 60674
rect 5630 60622 5682 60674
rect 5682 60622 5684 60674
rect 5628 60620 5684 60622
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 3500 59388 3556 59444
rect 8876 64652 8932 64708
rect 9324 64706 9380 64708
rect 9324 64654 9326 64706
rect 9326 64654 9378 64706
rect 9378 64654 9380 64706
rect 9324 64652 9380 64654
rect 6524 63026 6580 63028
rect 6524 62974 6526 63026
rect 6526 62974 6578 63026
rect 6578 62974 6580 63026
rect 6524 62972 6580 62974
rect 7308 62972 7364 63028
rect 7644 63026 7700 63028
rect 7644 62974 7646 63026
rect 7646 62974 7698 63026
rect 7698 62974 7700 63026
rect 7644 62972 7700 62974
rect 6748 62300 6804 62356
rect 7084 62354 7140 62356
rect 7084 62302 7086 62354
rect 7086 62302 7138 62354
rect 7138 62302 7140 62354
rect 7084 62300 7140 62302
rect 11788 64540 11844 64596
rect 11452 64034 11508 64036
rect 11452 63982 11454 64034
rect 11454 63982 11506 64034
rect 11506 63982 11508 64034
rect 11452 63980 11508 63982
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 20188 65490 20244 65492
rect 20188 65438 20190 65490
rect 20190 65438 20242 65490
rect 20242 65438 20244 65490
rect 20188 65436 20244 65438
rect 17612 65324 17668 65380
rect 12572 64652 12628 64708
rect 12124 63980 12180 64036
rect 9996 63308 10052 63364
rect 12236 64428 12292 64484
rect 12348 63362 12404 63364
rect 12348 63310 12350 63362
rect 12350 63310 12402 63362
rect 12402 63310 12404 63362
rect 12348 63308 12404 63310
rect 12684 64594 12740 64596
rect 12684 64542 12686 64594
rect 12686 64542 12738 64594
rect 12738 64542 12740 64594
rect 12684 64540 12740 64542
rect 12796 64482 12852 64484
rect 12796 64430 12798 64482
rect 12798 64430 12850 64482
rect 12850 64430 12852 64482
rect 12796 64428 12852 64430
rect 12572 63868 12628 63924
rect 12460 62914 12516 62916
rect 12460 62862 12462 62914
rect 12462 62862 12514 62914
rect 12514 62862 12516 62914
rect 12460 62860 12516 62862
rect 8540 62466 8596 62468
rect 8540 62414 8542 62466
rect 8542 62414 8594 62466
rect 8594 62414 8596 62466
rect 8540 62412 8596 62414
rect 10892 62466 10948 62468
rect 10892 62414 10894 62466
rect 10894 62414 10946 62466
rect 10946 62414 10948 62466
rect 10892 62412 10948 62414
rect 8092 62300 8148 62356
rect 10220 62354 10276 62356
rect 10220 62302 10222 62354
rect 10222 62302 10274 62354
rect 10274 62302 10276 62354
rect 10220 62300 10276 62302
rect 7868 62188 7924 62244
rect 10556 62242 10612 62244
rect 10556 62190 10558 62242
rect 10558 62190 10610 62242
rect 10610 62190 10612 62242
rect 10556 62188 10612 62190
rect 6188 61346 6244 61348
rect 6188 61294 6190 61346
rect 6190 61294 6242 61346
rect 6242 61294 6244 61346
rect 6188 61292 6244 61294
rect 6300 60620 6356 60676
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4844 58716 4900 58772
rect 2828 58604 2884 58660
rect 1820 47516 1876 47572
rect 3836 58322 3892 58324
rect 3836 58270 3838 58322
rect 3838 58270 3890 58322
rect 3890 58270 3892 58322
rect 3836 58268 3892 58270
rect 4060 58268 4116 58324
rect 2492 58156 2548 58212
rect 3948 58210 4004 58212
rect 3948 58158 3950 58210
rect 3950 58158 4002 58210
rect 4002 58158 4004 58210
rect 3948 58156 4004 58158
rect 4620 57538 4676 57540
rect 4620 57486 4622 57538
rect 4622 57486 4674 57538
rect 4674 57486 4676 57538
rect 4620 57484 4676 57486
rect 6860 61346 6916 61348
rect 6860 61294 6862 61346
rect 6862 61294 6914 61346
rect 6914 61294 6916 61346
rect 6860 61292 6916 61294
rect 5852 58716 5908 58772
rect 6636 58716 6692 58772
rect 4956 58268 5012 58324
rect 5628 57484 5684 57540
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4844 56924 4900 56980
rect 5516 56924 5572 56980
rect 4620 55970 4676 55972
rect 4620 55918 4622 55970
rect 4622 55918 4674 55970
rect 4674 55918 4676 55970
rect 4620 55916 4676 55918
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 5292 56812 5348 56868
rect 5180 55970 5236 55972
rect 5180 55918 5182 55970
rect 5182 55918 5234 55970
rect 5234 55918 5236 55970
rect 5180 55916 5236 55918
rect 3164 55020 3220 55076
rect 3836 55074 3892 55076
rect 3836 55022 3838 55074
rect 3838 55022 3890 55074
rect 3890 55022 3892 55074
rect 3836 55020 3892 55022
rect 3276 54572 3332 54628
rect 4060 54572 4116 54628
rect 4620 54460 4676 54516
rect 3388 53900 3444 53956
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4284 53900 4340 53956
rect 4284 53004 4340 53060
rect 5180 54514 5236 54516
rect 5180 54462 5182 54514
rect 5182 54462 5234 54514
rect 5234 54462 5236 54514
rect 5180 54460 5236 54462
rect 5852 57036 5908 57092
rect 6188 57036 6244 57092
rect 6748 56866 6804 56868
rect 6748 56814 6750 56866
rect 6750 56814 6802 56866
rect 6802 56814 6804 56866
rect 6748 56812 6804 56814
rect 6860 56700 6916 56756
rect 6188 55468 6244 55524
rect 6636 55916 6692 55972
rect 7644 59442 7700 59444
rect 7644 59390 7646 59442
rect 7646 59390 7698 59442
rect 7698 59390 7700 59442
rect 7644 59388 7700 59390
rect 7532 59330 7588 59332
rect 7532 59278 7534 59330
rect 7534 59278 7586 59330
rect 7586 59278 7588 59330
rect 7532 59276 7588 59278
rect 10220 60732 10276 60788
rect 9100 60114 9156 60116
rect 9100 60062 9102 60114
rect 9102 60062 9154 60114
rect 9154 60062 9156 60114
rect 9100 60060 9156 60062
rect 8428 60002 8484 60004
rect 8428 59950 8430 60002
rect 8430 59950 8482 60002
rect 8482 59950 8484 60002
rect 8428 59948 8484 59950
rect 8652 59948 8708 60004
rect 8204 59330 8260 59332
rect 8204 59278 8206 59330
rect 8206 59278 8258 59330
rect 8258 59278 8260 59330
rect 8204 59276 8260 59278
rect 8428 57596 8484 57652
rect 8204 56252 8260 56308
rect 8316 56194 8372 56196
rect 8316 56142 8318 56194
rect 8318 56142 8370 56194
rect 8370 56142 8372 56194
rect 8316 56140 8372 56142
rect 13804 64594 13860 64596
rect 13804 64542 13806 64594
rect 13806 64542 13858 64594
rect 13858 64542 13860 64594
rect 13804 64540 13860 64542
rect 13468 64428 13524 64484
rect 13580 63922 13636 63924
rect 13580 63870 13582 63922
rect 13582 63870 13634 63922
rect 13634 63870 13636 63922
rect 13580 63868 13636 63870
rect 19516 65378 19572 65380
rect 19516 65326 19518 65378
rect 19518 65326 19570 65378
rect 19570 65326 19572 65378
rect 19516 65324 19572 65326
rect 17948 64706 18004 64708
rect 17948 64654 17950 64706
rect 17950 64654 18002 64706
rect 18002 64654 18004 64706
rect 17948 64652 18004 64654
rect 20860 65436 20916 65492
rect 20188 64652 20244 64708
rect 16716 63980 16772 64036
rect 13692 62914 13748 62916
rect 13692 62862 13694 62914
rect 13694 62862 13746 62914
rect 13746 62862 13748 62914
rect 13692 62860 13748 62862
rect 13692 62300 13748 62356
rect 13916 63084 13972 63140
rect 15484 63138 15540 63140
rect 15484 63086 15486 63138
rect 15486 63086 15538 63138
rect 15538 63086 15540 63138
rect 15484 63084 15540 63086
rect 16268 62860 16324 62916
rect 15148 62354 15204 62356
rect 15148 62302 15150 62354
rect 15150 62302 15202 62354
rect 15202 62302 15204 62354
rect 15148 62300 15204 62302
rect 16380 63026 16436 63028
rect 16380 62974 16382 63026
rect 16382 62974 16434 63026
rect 16434 62974 16436 63026
rect 16380 62972 16436 62974
rect 17724 64034 17780 64036
rect 17724 63982 17726 64034
rect 17726 63982 17778 64034
rect 17778 63982 17780 64034
rect 17724 63980 17780 63982
rect 16828 63922 16884 63924
rect 16828 63870 16830 63922
rect 16830 63870 16882 63922
rect 16882 63870 16884 63922
rect 16828 63868 16884 63870
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 20860 64428 20916 64484
rect 17276 63084 17332 63140
rect 17612 63026 17668 63028
rect 17612 62974 17614 63026
rect 17614 62974 17666 63026
rect 17666 62974 17668 63026
rect 17612 62972 17668 62974
rect 17388 62914 17444 62916
rect 17388 62862 17390 62914
rect 17390 62862 17442 62914
rect 17442 62862 17444 62914
rect 17388 62860 17444 62862
rect 11004 60898 11060 60900
rect 11004 60846 11006 60898
rect 11006 60846 11058 60898
rect 11058 60846 11060 60898
rect 11004 60844 11060 60846
rect 10780 60786 10836 60788
rect 10780 60734 10782 60786
rect 10782 60734 10834 60786
rect 10834 60734 10836 60786
rect 10780 60732 10836 60734
rect 10556 60172 10612 60228
rect 11340 59948 11396 60004
rect 11788 60114 11844 60116
rect 11788 60062 11790 60114
rect 11790 60062 11842 60114
rect 11842 60062 11844 60114
rect 11788 60060 11844 60062
rect 11340 59276 11396 59332
rect 13244 60898 13300 60900
rect 13244 60846 13246 60898
rect 13246 60846 13298 60898
rect 13298 60846 13300 60898
rect 13244 60844 13300 60846
rect 13356 60786 13412 60788
rect 13356 60734 13358 60786
rect 13358 60734 13410 60786
rect 13410 60734 13412 60786
rect 13356 60732 13412 60734
rect 12908 60002 12964 60004
rect 12908 59950 12910 60002
rect 12910 59950 12962 60002
rect 12962 59950 12964 60002
rect 12908 59948 12964 59950
rect 14588 60732 14644 60788
rect 12460 59724 12516 59780
rect 11004 58268 11060 58324
rect 9436 57650 9492 57652
rect 9436 57598 9438 57650
rect 9438 57598 9490 57650
rect 9490 57598 9492 57650
rect 9436 57596 9492 57598
rect 10108 57650 10164 57652
rect 10108 57598 10110 57650
rect 10110 57598 10162 57650
rect 10162 57598 10164 57650
rect 10108 57596 10164 57598
rect 9996 57036 10052 57092
rect 8652 56812 8708 56868
rect 9772 56812 9828 56868
rect 8764 56700 8820 56756
rect 8764 56306 8820 56308
rect 8764 56254 8766 56306
rect 8766 56254 8818 56306
rect 8818 56254 8820 56306
rect 8764 56252 8820 56254
rect 9884 56754 9940 56756
rect 9884 56702 9886 56754
rect 9886 56702 9938 56754
rect 9938 56702 9940 56754
rect 9884 56700 9940 56702
rect 9212 56140 9268 56196
rect 5404 54626 5460 54628
rect 5404 54574 5406 54626
rect 5406 54574 5458 54626
rect 5458 54574 5460 54626
rect 5404 54572 5460 54574
rect 4956 53004 5012 53060
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 3836 52108 3892 52164
rect 3276 51212 3332 51268
rect 3388 51324 3444 51380
rect 2492 49980 2548 50036
rect 3612 50540 3668 50596
rect 4620 52162 4676 52164
rect 4620 52110 4622 52162
rect 4622 52110 4674 52162
rect 4674 52110 4676 52162
rect 4620 52108 4676 52110
rect 2716 46562 2772 46564
rect 2716 46510 2718 46562
rect 2718 46510 2770 46562
rect 2770 46510 2772 46562
rect 2716 46508 2772 46510
rect 3500 46562 3556 46564
rect 3500 46510 3502 46562
rect 3502 46510 3554 46562
rect 3554 46510 3556 46562
rect 3500 46508 3556 46510
rect 3388 44380 3444 44436
rect 3948 51212 4004 51268
rect 4396 51100 4452 51156
rect 5068 51378 5124 51380
rect 5068 51326 5070 51378
rect 5070 51326 5122 51378
rect 5122 51326 5124 51378
rect 5068 51324 5124 51326
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4060 50428 4116 50484
rect 4284 50316 4340 50372
rect 4732 50204 4788 50260
rect 4508 50034 4564 50036
rect 4508 49982 4510 50034
rect 4510 49982 4562 50034
rect 4562 49982 4564 50034
rect 4508 49980 4564 49982
rect 5964 53452 6020 53508
rect 5516 51266 5572 51268
rect 5516 51214 5518 51266
rect 5518 51214 5570 51266
rect 5570 51214 5572 51266
rect 5516 51212 5572 51214
rect 5516 50652 5572 50708
rect 5628 50594 5684 50596
rect 5628 50542 5630 50594
rect 5630 50542 5682 50594
rect 5682 50542 5684 50594
rect 5628 50540 5684 50542
rect 5740 50482 5796 50484
rect 5740 50430 5742 50482
rect 5742 50430 5794 50482
rect 5794 50430 5796 50482
rect 5740 50428 5796 50430
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 5404 48972 5460 49028
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 6076 49026 6132 49028
rect 6076 48974 6078 49026
rect 6078 48974 6130 49026
rect 6130 48974 6132 49026
rect 6076 48972 6132 48974
rect 5068 47570 5124 47572
rect 5068 47518 5070 47570
rect 5070 47518 5122 47570
rect 5122 47518 5124 47570
rect 5068 47516 5124 47518
rect 4620 47292 4676 47348
rect 5292 47292 5348 47348
rect 2380 43708 2436 43764
rect 1820 42028 1876 42084
rect 1820 37436 1876 37492
rect 1820 35026 1876 35028
rect 1820 34974 1822 35026
rect 1822 34974 1874 35026
rect 1874 34974 1876 35026
rect 1820 34972 1876 34974
rect 2604 43708 2660 43764
rect 3612 43596 3668 43652
rect 2828 41356 2884 41412
rect 3276 41356 3332 41412
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4508 44380 4564 44436
rect 5292 44492 5348 44548
rect 4844 44268 4900 44324
rect 5068 43650 5124 43652
rect 5068 43598 5070 43650
rect 5070 43598 5122 43650
rect 5122 43598 5124 43650
rect 5068 43596 5124 43598
rect 5740 47346 5796 47348
rect 5740 47294 5742 47346
rect 5742 47294 5794 47346
rect 5794 47294 5796 47346
rect 5740 47292 5796 47294
rect 5516 46956 5572 47012
rect 6300 46956 6356 47012
rect 6076 45106 6132 45108
rect 6076 45054 6078 45106
rect 6078 45054 6130 45106
rect 6130 45054 6132 45106
rect 6076 45052 6132 45054
rect 5964 44546 6020 44548
rect 5964 44494 5966 44546
rect 5966 44494 6018 44546
rect 6018 44494 6020 44546
rect 5964 44492 6020 44494
rect 5628 44434 5684 44436
rect 5628 44382 5630 44434
rect 5630 44382 5682 44434
rect 5682 44382 5684 44434
rect 5628 44380 5684 44382
rect 6188 44322 6244 44324
rect 6188 44270 6190 44322
rect 6190 44270 6242 44322
rect 6242 44270 6244 44322
rect 6188 44268 6244 44270
rect 5516 43650 5572 43652
rect 5516 43598 5518 43650
rect 5518 43598 5570 43650
rect 5570 43598 5572 43650
rect 5516 43596 5572 43598
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5068 42028 5124 42084
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 3836 39676 3892 39732
rect 3164 39618 3220 39620
rect 3164 39566 3166 39618
rect 3166 39566 3218 39618
rect 3218 39566 3220 39618
rect 3164 39564 3220 39566
rect 5404 42028 5460 42084
rect 6076 41858 6132 41860
rect 6076 41806 6078 41858
rect 6078 41806 6130 41858
rect 6130 41806 6132 41858
rect 6076 41804 6132 41806
rect 4172 39788 4228 39844
rect 4620 40290 4676 40292
rect 4620 40238 4622 40290
rect 4622 40238 4674 40290
rect 4674 40238 4676 40290
rect 4620 40236 4676 40238
rect 3948 39564 4004 39620
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4396 39676 4452 39732
rect 4620 39730 4676 39732
rect 4620 39678 4622 39730
rect 4622 39678 4674 39730
rect 4674 39678 4676 39730
rect 4620 39676 4676 39678
rect 4396 38668 4452 38724
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4060 38050 4116 38052
rect 4060 37998 4062 38050
rect 4062 37998 4114 38050
rect 4114 37998 4116 38050
rect 4060 37996 4116 37998
rect 2716 37548 2772 37604
rect 3612 37548 3668 37604
rect 3052 37378 3108 37380
rect 3052 37326 3054 37378
rect 3054 37326 3106 37378
rect 3106 37326 3108 37378
rect 3052 37324 3108 37326
rect 3948 37324 4004 37380
rect 3164 37266 3220 37268
rect 3164 37214 3166 37266
rect 3166 37214 3218 37266
rect 3218 37214 3220 37266
rect 3164 37212 3220 37214
rect 3724 37266 3780 37268
rect 3724 37214 3726 37266
rect 3726 37214 3778 37266
rect 3778 37214 3780 37266
rect 3724 37212 3780 37214
rect 4620 37436 4676 37492
rect 5852 40908 5908 40964
rect 5740 40236 5796 40292
rect 5628 39842 5684 39844
rect 5628 39790 5630 39842
rect 5630 39790 5682 39842
rect 5682 39790 5684 39842
rect 5628 39788 5684 39790
rect 6524 40908 6580 40964
rect 6188 39676 6244 39732
rect 6748 54348 6804 54404
rect 7420 53618 7476 53620
rect 7420 53566 7422 53618
rect 7422 53566 7474 53618
rect 7474 53566 7476 53618
rect 7420 53564 7476 53566
rect 7196 53506 7252 53508
rect 7196 53454 7198 53506
rect 7198 53454 7250 53506
rect 7250 53454 7252 53506
rect 7196 53452 7252 53454
rect 7868 53564 7924 53620
rect 9100 53564 9156 53620
rect 7644 53116 7700 53172
rect 7308 52780 7364 52836
rect 6748 52108 6804 52164
rect 8652 53116 8708 53172
rect 8428 52946 8484 52948
rect 8428 52894 8430 52946
rect 8430 52894 8482 52946
rect 8482 52894 8484 52946
rect 8428 52892 8484 52894
rect 8652 52946 8708 52948
rect 8652 52894 8654 52946
rect 8654 52894 8706 52946
rect 8706 52894 8708 52946
rect 8652 52892 8708 52894
rect 8204 52274 8260 52276
rect 8204 52222 8206 52274
rect 8206 52222 8258 52274
rect 8258 52222 8260 52274
rect 8204 52220 8260 52222
rect 7980 51996 8036 52052
rect 7644 51100 7700 51156
rect 6748 48914 6804 48916
rect 6748 48862 6750 48914
rect 6750 48862 6802 48914
rect 6802 48862 6804 48914
rect 6748 48860 6804 48862
rect 7532 45164 7588 45220
rect 7196 44380 7252 44436
rect 7084 40348 7140 40404
rect 6188 39058 6244 39060
rect 6188 39006 6190 39058
rect 6190 39006 6242 39058
rect 6242 39006 6244 39058
rect 6188 39004 6244 39006
rect 6860 39004 6916 39060
rect 5852 38780 5908 38836
rect 6636 38834 6692 38836
rect 6636 38782 6638 38834
rect 6638 38782 6690 38834
rect 6690 38782 6692 38834
rect 6636 38780 6692 38782
rect 6412 38556 6468 38612
rect 7084 38556 7140 38612
rect 7420 38722 7476 38724
rect 7420 38670 7422 38722
rect 7422 38670 7474 38722
rect 7474 38670 7476 38722
rect 7420 38668 7476 38670
rect 9100 52892 9156 52948
rect 10444 57036 10500 57092
rect 10668 57650 10724 57652
rect 10668 57598 10670 57650
rect 10670 57598 10722 57650
rect 10722 57598 10724 57650
rect 10668 57596 10724 57598
rect 10780 57036 10836 57092
rect 10332 55468 10388 55524
rect 11788 58268 11844 58324
rect 12236 58716 12292 58772
rect 11228 56588 11284 56644
rect 11788 56028 11844 56084
rect 11004 55468 11060 55524
rect 11340 55298 11396 55300
rect 11340 55246 11342 55298
rect 11342 55246 11394 55298
rect 11394 55246 11396 55298
rect 11340 55244 11396 55246
rect 9996 53004 10052 53060
rect 8652 52220 8708 52276
rect 8764 52050 8820 52052
rect 8764 51998 8766 52050
rect 8766 51998 8818 52050
rect 8818 51998 8820 52050
rect 8764 51996 8820 51998
rect 8652 49868 8708 49924
rect 8540 49084 8596 49140
rect 8428 48748 8484 48804
rect 8316 48466 8372 48468
rect 8316 48414 8318 48466
rect 8318 48414 8370 48466
rect 8370 48414 8372 48466
rect 8316 48412 8372 48414
rect 8092 48354 8148 48356
rect 8092 48302 8094 48354
rect 8094 48302 8146 48354
rect 8146 48302 8148 48354
rect 8092 48300 8148 48302
rect 8876 49810 8932 49812
rect 8876 49758 8878 49810
rect 8878 49758 8930 49810
rect 8930 49758 8932 49810
rect 8876 49756 8932 49758
rect 9660 52162 9716 52164
rect 9660 52110 9662 52162
rect 9662 52110 9714 52162
rect 9714 52110 9716 52162
rect 9660 52108 9716 52110
rect 10332 53004 10388 53060
rect 10668 52834 10724 52836
rect 10668 52782 10670 52834
rect 10670 52782 10722 52834
rect 10722 52782 10724 52834
rect 10668 52780 10724 52782
rect 10108 52220 10164 52276
rect 10220 52162 10276 52164
rect 10220 52110 10222 52162
rect 10222 52110 10274 52162
rect 10274 52110 10276 52162
rect 10220 52108 10276 52110
rect 11452 52220 11508 52276
rect 11116 51100 11172 51156
rect 11788 51548 11844 51604
rect 11564 50876 11620 50932
rect 9212 49868 9268 49924
rect 11564 50706 11620 50708
rect 11564 50654 11566 50706
rect 11566 50654 11618 50706
rect 11618 50654 11620 50706
rect 11564 50652 11620 50654
rect 9324 49756 9380 49812
rect 8764 48300 8820 48356
rect 9100 49084 9156 49140
rect 8092 44434 8148 44436
rect 8092 44382 8094 44434
rect 8094 44382 8146 44434
rect 8146 44382 8148 44434
rect 8092 44380 8148 44382
rect 8316 45276 8372 45332
rect 8764 45612 8820 45668
rect 8876 45276 8932 45332
rect 8988 45612 9044 45668
rect 8428 43596 8484 43652
rect 8876 42754 8932 42756
rect 8876 42702 8878 42754
rect 8878 42702 8930 42754
rect 8930 42702 8932 42754
rect 8876 42700 8932 42702
rect 8764 42476 8820 42532
rect 8204 41916 8260 41972
rect 8876 41916 8932 41972
rect 8764 41858 8820 41860
rect 8764 41806 8766 41858
rect 8766 41806 8818 41858
rect 8818 41806 8820 41858
rect 8764 41804 8820 41806
rect 8988 41804 9044 41860
rect 8540 41186 8596 41188
rect 8540 41134 8542 41186
rect 8542 41134 8594 41186
rect 8594 41134 8596 41186
rect 8540 41132 8596 41134
rect 7868 40402 7924 40404
rect 7868 40350 7870 40402
rect 7870 40350 7922 40402
rect 7922 40350 7924 40402
rect 7868 40348 7924 40350
rect 8540 40348 8596 40404
rect 8540 39116 8596 39172
rect 7868 38834 7924 38836
rect 7868 38782 7870 38834
rect 7870 38782 7922 38834
rect 7922 38782 7924 38834
rect 7868 38780 7924 38782
rect 9324 48914 9380 48916
rect 9324 48862 9326 48914
rect 9326 48862 9378 48914
rect 9378 48862 9380 48914
rect 9324 48860 9380 48862
rect 10220 49922 10276 49924
rect 10220 49870 10222 49922
rect 10222 49870 10274 49922
rect 10274 49870 10276 49922
rect 10220 49868 10276 49870
rect 10332 49810 10388 49812
rect 10332 49758 10334 49810
rect 10334 49758 10386 49810
rect 10386 49758 10388 49810
rect 10332 49756 10388 49758
rect 10780 49644 10836 49700
rect 9660 48748 9716 48804
rect 10108 48972 10164 49028
rect 9548 48412 9604 48468
rect 9548 47628 9604 47684
rect 9996 48300 10052 48356
rect 9660 47404 9716 47460
rect 10556 48354 10612 48356
rect 10556 48302 10558 48354
rect 10558 48302 10610 48354
rect 10610 48302 10612 48354
rect 10556 48300 10612 48302
rect 9436 45388 9492 45444
rect 9996 45612 10052 45668
rect 9772 45330 9828 45332
rect 9772 45278 9774 45330
rect 9774 45278 9826 45330
rect 9826 45278 9828 45330
rect 9772 45276 9828 45278
rect 9436 45052 9492 45108
rect 10108 45164 10164 45220
rect 9660 42754 9716 42756
rect 9660 42702 9662 42754
rect 9662 42702 9714 42754
rect 9714 42702 9716 42754
rect 9660 42700 9716 42702
rect 9772 42476 9828 42532
rect 9436 41916 9492 41972
rect 9884 42140 9940 42196
rect 10556 42140 10612 42196
rect 10332 41858 10388 41860
rect 10332 41806 10334 41858
rect 10334 41806 10386 41858
rect 10386 41806 10388 41858
rect 10332 41804 10388 41806
rect 10108 41132 10164 41188
rect 9884 38668 9940 38724
rect 7980 38556 8036 38612
rect 5068 37436 5124 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 7868 37490 7924 37492
rect 7868 37438 7870 37490
rect 7870 37438 7922 37490
rect 7922 37438 7924 37490
rect 7868 37436 7924 37438
rect 8428 37378 8484 37380
rect 8428 37326 8430 37378
rect 8430 37326 8482 37378
rect 8482 37326 8484 37378
rect 8428 37324 8484 37326
rect 7980 36988 8036 37044
rect 8204 36428 8260 36484
rect 2268 35810 2324 35812
rect 2268 35758 2270 35810
rect 2270 35758 2322 35810
rect 2322 35758 2324 35810
rect 2268 35756 2324 35758
rect 7868 35644 7924 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 5852 34860 5908 34916
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 5068 28924 5124 28980
rect 4284 28588 4340 28644
rect 4732 28588 4788 28644
rect 5404 27746 5460 27748
rect 5404 27694 5406 27746
rect 5406 27694 5458 27746
rect 5458 27694 5460 27746
rect 5404 27692 5460 27694
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2268 26236 2324 26292
rect 5628 27020 5684 27076
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 7532 34802 7588 34804
rect 7532 34750 7534 34802
rect 7534 34750 7586 34802
rect 7586 34750 7588 34802
rect 7532 34748 7588 34750
rect 8092 35420 8148 35476
rect 7420 33852 7476 33908
rect 6972 28642 7028 28644
rect 6972 28590 6974 28642
rect 6974 28590 7026 28642
rect 7026 28590 7028 28642
rect 6972 28588 7028 28590
rect 6748 27074 6804 27076
rect 6748 27022 6750 27074
rect 6750 27022 6802 27074
rect 6802 27022 6804 27074
rect 6748 27020 6804 27022
rect 7308 31890 7364 31892
rect 7308 31838 7310 31890
rect 7310 31838 7362 31890
rect 7362 31838 7364 31890
rect 7308 31836 7364 31838
rect 7196 29372 7252 29428
rect 8988 37490 9044 37492
rect 8988 37438 8990 37490
rect 8990 37438 9042 37490
rect 9042 37438 9044 37490
rect 8988 37436 9044 37438
rect 9436 37436 9492 37492
rect 8428 36204 8484 36260
rect 9548 37324 9604 37380
rect 9660 37042 9716 37044
rect 9660 36990 9662 37042
rect 9662 36990 9714 37042
rect 9714 36990 9716 37042
rect 9660 36988 9716 36990
rect 8764 36428 8820 36484
rect 8764 36258 8820 36260
rect 8764 36206 8766 36258
rect 8766 36206 8818 36258
rect 8818 36206 8820 36258
rect 8764 36204 8820 36206
rect 8876 35980 8932 36036
rect 7980 33852 8036 33908
rect 7868 31836 7924 31892
rect 7868 31276 7924 31332
rect 7980 32508 8036 32564
rect 9772 36092 9828 36148
rect 9996 37436 10052 37492
rect 11116 48242 11172 48244
rect 11116 48190 11118 48242
rect 11118 48190 11170 48242
rect 11170 48190 11172 48242
rect 11116 48188 11172 48190
rect 11116 47682 11172 47684
rect 11116 47630 11118 47682
rect 11118 47630 11170 47682
rect 11170 47630 11172 47682
rect 11116 47628 11172 47630
rect 11340 48300 11396 48356
rect 11116 47458 11172 47460
rect 11116 47406 11118 47458
rect 11118 47406 11170 47458
rect 11170 47406 11172 47458
rect 11116 47404 11172 47406
rect 11788 47404 11844 47460
rect 11340 47292 11396 47348
rect 11788 46844 11844 46900
rect 11564 42082 11620 42084
rect 11564 42030 11566 42082
rect 11566 42030 11618 42082
rect 11618 42030 11620 42082
rect 11564 42028 11620 42030
rect 11676 41020 11732 41076
rect 11452 38892 11508 38948
rect 11564 38722 11620 38724
rect 11564 38670 11566 38722
rect 11566 38670 11618 38722
rect 11618 38670 11620 38722
rect 11564 38668 11620 38670
rect 12796 59276 12852 59332
rect 12796 58828 12852 58884
rect 14028 59724 14084 59780
rect 13804 57762 13860 57764
rect 13804 57710 13806 57762
rect 13806 57710 13858 57762
rect 13858 57710 13860 57762
rect 13804 57708 13860 57710
rect 13356 57596 13412 57652
rect 13916 57650 13972 57652
rect 13916 57598 13918 57650
rect 13918 57598 13970 57650
rect 13970 57598 13972 57650
rect 13916 57596 13972 57598
rect 12236 57090 12292 57092
rect 12236 57038 12238 57090
rect 12238 57038 12290 57090
rect 12290 57038 12292 57090
rect 12236 57036 12292 57038
rect 12012 56588 12068 56644
rect 12572 56642 12628 56644
rect 12572 56590 12574 56642
rect 12574 56590 12626 56642
rect 12626 56590 12628 56642
rect 12572 56588 12628 56590
rect 12908 56028 12964 56084
rect 12684 55074 12740 55076
rect 12684 55022 12686 55074
rect 12686 55022 12738 55074
rect 12738 55022 12740 55074
rect 12684 55020 12740 55022
rect 12572 54460 12628 54516
rect 13692 56700 13748 56756
rect 15596 60060 15652 60116
rect 15708 60508 15764 60564
rect 15148 59948 15204 60004
rect 15036 59442 15092 59444
rect 15036 59390 15038 59442
rect 15038 59390 15090 59442
rect 15090 59390 15092 59442
rect 15036 59388 15092 59390
rect 14588 58716 14644 58772
rect 17836 62914 17892 62916
rect 17836 62862 17838 62914
rect 17838 62862 17890 62914
rect 17890 62862 17892 62914
rect 17836 62860 17892 62862
rect 18508 62914 18564 62916
rect 18508 62862 18510 62914
rect 18510 62862 18562 62914
rect 18562 62862 18564 62914
rect 18508 62860 18564 62862
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 18956 62466 19012 62468
rect 18956 62414 18958 62466
rect 18958 62414 19010 62466
rect 19010 62414 19012 62466
rect 18956 62412 19012 62414
rect 24892 66444 24948 66500
rect 26124 66498 26180 66500
rect 26124 66446 26126 66498
rect 26126 66446 26178 66498
rect 26178 66446 26180 66498
rect 26124 66444 26180 66446
rect 21420 64482 21476 64484
rect 21420 64430 21422 64482
rect 21422 64430 21474 64482
rect 21474 64430 21476 64482
rect 21420 64428 21476 64430
rect 22540 64876 22596 64932
rect 21868 64428 21924 64484
rect 23548 64930 23604 64932
rect 23548 64878 23550 64930
rect 23550 64878 23602 64930
rect 23602 64878 23604 64930
rect 23548 64876 23604 64878
rect 23212 64482 23268 64484
rect 23212 64430 23214 64482
rect 23214 64430 23266 64482
rect 23266 64430 23268 64482
rect 23212 64428 23268 64430
rect 23996 64428 24052 64484
rect 21084 63308 21140 63364
rect 22316 63362 22372 63364
rect 22316 63310 22318 63362
rect 22318 63310 22370 63362
rect 22370 63310 22372 63362
rect 22316 63308 22372 63310
rect 22092 62860 22148 62916
rect 18172 62300 18228 62356
rect 16268 60844 16324 60900
rect 16156 59890 16212 59892
rect 16156 59838 16158 59890
rect 16158 59838 16210 59890
rect 16210 59838 16212 59890
rect 16156 59836 16212 59838
rect 17500 60898 17556 60900
rect 17500 60846 17502 60898
rect 17502 60846 17554 60898
rect 17554 60846 17556 60898
rect 17500 60844 17556 60846
rect 17612 60226 17668 60228
rect 17612 60174 17614 60226
rect 17614 60174 17666 60226
rect 17666 60174 17668 60226
rect 17612 60172 17668 60174
rect 16716 59724 16772 59780
rect 14924 57708 14980 57764
rect 15372 58210 15428 58212
rect 15372 58158 15374 58210
rect 15374 58158 15426 58210
rect 15426 58158 15428 58210
rect 15372 58156 15428 58158
rect 14252 56754 14308 56756
rect 14252 56702 14254 56754
rect 14254 56702 14306 56754
rect 14306 56702 14308 56754
rect 14252 56700 14308 56702
rect 15148 56754 15204 56756
rect 15148 56702 15150 56754
rect 15150 56702 15202 56754
rect 15202 56702 15204 56754
rect 15148 56700 15204 56702
rect 13916 56588 13972 56644
rect 13356 56194 13412 56196
rect 13356 56142 13358 56194
rect 13358 56142 13410 56194
rect 13410 56142 13412 56194
rect 13356 56140 13412 56142
rect 13132 55916 13188 55972
rect 12348 52780 12404 52836
rect 12236 50652 12292 50708
rect 12684 49810 12740 49812
rect 12684 49758 12686 49810
rect 12686 49758 12738 49810
rect 12738 49758 12740 49810
rect 12684 49756 12740 49758
rect 12348 49698 12404 49700
rect 12348 49646 12350 49698
rect 12350 49646 12402 49698
rect 12402 49646 12404 49698
rect 12348 49644 12404 49646
rect 12572 48188 12628 48244
rect 12236 47458 12292 47460
rect 12236 47406 12238 47458
rect 12238 47406 12290 47458
rect 12290 47406 12292 47458
rect 12236 47404 12292 47406
rect 12908 53004 12964 53060
rect 14700 56642 14756 56644
rect 14700 56590 14702 56642
rect 14702 56590 14754 56642
rect 14754 56590 14756 56642
rect 14700 56588 14756 56590
rect 14028 56194 14084 56196
rect 14028 56142 14030 56194
rect 14030 56142 14082 56194
rect 14082 56142 14084 56194
rect 14028 56140 14084 56142
rect 13468 55244 13524 55300
rect 13580 55074 13636 55076
rect 13580 55022 13582 55074
rect 13582 55022 13634 55074
rect 13634 55022 13636 55074
rect 13580 55020 13636 55022
rect 13356 54124 13412 54180
rect 14588 56082 14644 56084
rect 14588 56030 14590 56082
rect 14590 56030 14642 56082
rect 14642 56030 14644 56082
rect 14588 56028 14644 56030
rect 14252 55916 14308 55972
rect 15260 55970 15316 55972
rect 15260 55918 15262 55970
rect 15262 55918 15314 55970
rect 15314 55918 15316 55970
rect 15260 55916 15316 55918
rect 14476 55298 14532 55300
rect 14476 55246 14478 55298
rect 14478 55246 14530 55298
rect 14530 55246 14532 55298
rect 14476 55244 14532 55246
rect 14476 54514 14532 54516
rect 14476 54462 14478 54514
rect 14478 54462 14530 54514
rect 14530 54462 14532 54514
rect 14476 54460 14532 54462
rect 14140 54124 14196 54180
rect 15484 54514 15540 54516
rect 15484 54462 15486 54514
rect 15486 54462 15538 54514
rect 15538 54462 15540 54514
rect 15484 54460 15540 54462
rect 14812 53058 14868 53060
rect 14812 53006 14814 53058
rect 14814 53006 14866 53058
rect 14866 53006 14868 53058
rect 14812 53004 14868 53006
rect 12908 51772 12964 51828
rect 13468 51772 13524 51828
rect 13356 51602 13412 51604
rect 13356 51550 13358 51602
rect 13358 51550 13410 51602
rect 13410 51550 13412 51602
rect 13356 51548 13412 51550
rect 13916 51548 13972 51604
rect 14476 52162 14532 52164
rect 14476 52110 14478 52162
rect 14478 52110 14530 52162
rect 14530 52110 14532 52162
rect 14476 52108 14532 52110
rect 14364 51436 14420 51492
rect 14924 52220 14980 52276
rect 15260 52162 15316 52164
rect 15260 52110 15262 52162
rect 15262 52110 15314 52162
rect 15314 52110 15316 52162
rect 15260 52108 15316 52110
rect 15036 51490 15092 51492
rect 15036 51438 15038 51490
rect 15038 51438 15090 51490
rect 15090 51438 15092 51490
rect 15036 51436 15092 51438
rect 11900 46060 11956 46116
rect 12796 46060 12852 46116
rect 12796 45388 12852 45444
rect 12460 45330 12516 45332
rect 12460 45278 12462 45330
rect 12462 45278 12514 45330
rect 12514 45278 12516 45330
rect 12460 45276 12516 45278
rect 13244 49810 13300 49812
rect 13244 49758 13246 49810
rect 13246 49758 13298 49810
rect 13298 49758 13300 49810
rect 13244 49756 13300 49758
rect 13692 49644 13748 49700
rect 13356 48242 13412 48244
rect 13356 48190 13358 48242
rect 13358 48190 13410 48242
rect 13410 48190 13412 48242
rect 13356 48188 13412 48190
rect 13356 47852 13412 47908
rect 13692 48130 13748 48132
rect 13692 48078 13694 48130
rect 13694 48078 13746 48130
rect 13746 48078 13748 48130
rect 13692 48076 13748 48078
rect 13692 47852 13748 47908
rect 13356 47458 13412 47460
rect 13356 47406 13358 47458
rect 13358 47406 13410 47458
rect 13410 47406 13412 47458
rect 13356 47404 13412 47406
rect 13132 46844 13188 46900
rect 13580 47346 13636 47348
rect 13580 47294 13582 47346
rect 13582 47294 13634 47346
rect 13634 47294 13636 47346
rect 13580 47292 13636 47294
rect 13468 46956 13524 47012
rect 13132 46620 13188 46676
rect 13580 45948 13636 46004
rect 13580 45388 13636 45444
rect 13916 49698 13972 49700
rect 13916 49646 13918 49698
rect 13918 49646 13970 49698
rect 13970 49646 13972 49698
rect 13916 49644 13972 49646
rect 14364 49810 14420 49812
rect 14364 49758 14366 49810
rect 14366 49758 14418 49810
rect 14418 49758 14420 49810
rect 14364 49756 14420 49758
rect 14028 47458 14084 47460
rect 14028 47406 14030 47458
rect 14030 47406 14082 47458
rect 14082 47406 14084 47458
rect 14028 47404 14084 47406
rect 14028 46060 14084 46116
rect 14028 45164 14084 45220
rect 12348 42530 12404 42532
rect 12348 42478 12350 42530
rect 12350 42478 12402 42530
rect 12402 42478 12404 42530
rect 12348 42476 12404 42478
rect 11900 41804 11956 41860
rect 12124 42140 12180 42196
rect 12236 42028 12292 42084
rect 11004 37996 11060 38052
rect 13468 44380 13524 44436
rect 13468 43484 13524 43540
rect 12908 42476 12964 42532
rect 13468 42140 13524 42196
rect 13580 43260 13636 43316
rect 12348 40962 12404 40964
rect 12348 40910 12350 40962
rect 12350 40910 12402 40962
rect 12402 40910 12404 40962
rect 12348 40908 12404 40910
rect 12684 41074 12740 41076
rect 12684 41022 12686 41074
rect 12686 41022 12738 41074
rect 12738 41022 12740 41074
rect 12684 41020 12740 41022
rect 12572 40684 12628 40740
rect 12796 40460 12852 40516
rect 9996 35980 10052 36036
rect 10556 35868 10612 35924
rect 9548 33516 9604 33572
rect 9212 32060 9268 32116
rect 7756 29986 7812 29988
rect 7756 29934 7758 29986
rect 7758 29934 7810 29986
rect 7810 29934 7812 29986
rect 7756 29932 7812 29934
rect 8092 29708 8148 29764
rect 7308 27356 7364 27412
rect 7980 27858 8036 27860
rect 7980 27806 7982 27858
rect 7982 27806 8034 27858
rect 8034 27806 8036 27858
rect 7980 27804 8036 27806
rect 8652 31890 8708 31892
rect 8652 31838 8654 31890
rect 8654 31838 8706 31890
rect 8706 31838 8708 31890
rect 8652 31836 8708 31838
rect 8428 30156 8484 30212
rect 7868 27298 7924 27300
rect 7868 27246 7870 27298
rect 7870 27246 7922 27298
rect 7922 27246 7924 27298
rect 7868 27244 7924 27246
rect 9884 33906 9940 33908
rect 9884 33854 9886 33906
rect 9886 33854 9938 33906
rect 9938 33854 9940 33906
rect 9884 33852 9940 33854
rect 10220 35308 10276 35364
rect 10444 35084 10500 35140
rect 11340 37378 11396 37380
rect 11340 37326 11342 37378
rect 11342 37326 11394 37378
rect 11394 37326 11396 37378
rect 11340 37324 11396 37326
rect 11004 37212 11060 37268
rect 10780 36258 10836 36260
rect 10780 36206 10782 36258
rect 10782 36206 10834 36258
rect 10834 36206 10836 36258
rect 10780 36204 10836 36206
rect 11004 36092 11060 36148
rect 11004 35532 11060 35588
rect 10220 33516 10276 33572
rect 10780 34748 10836 34804
rect 11564 36370 11620 36372
rect 11564 36318 11566 36370
rect 11566 36318 11618 36370
rect 11618 36318 11620 36370
rect 11564 36316 11620 36318
rect 12796 39788 12852 39844
rect 12124 39004 12180 39060
rect 12796 39004 12852 39060
rect 13580 40684 13636 40740
rect 13356 40514 13412 40516
rect 13356 40462 13358 40514
rect 13358 40462 13410 40514
rect 13410 40462 13412 40514
rect 13356 40460 13412 40462
rect 13804 42530 13860 42532
rect 13804 42478 13806 42530
rect 13806 42478 13858 42530
rect 13858 42478 13860 42530
rect 13804 42476 13860 42478
rect 13916 41020 13972 41076
rect 13804 40402 13860 40404
rect 13804 40350 13806 40402
rect 13806 40350 13858 40402
rect 13858 40350 13860 40402
rect 13804 40348 13860 40350
rect 13916 40236 13972 40292
rect 14140 43036 14196 43092
rect 14812 48076 14868 48132
rect 16156 58716 16212 58772
rect 16156 58156 16212 58212
rect 16044 57036 16100 57092
rect 17164 59388 17220 59444
rect 17612 59330 17668 59332
rect 17612 59278 17614 59330
rect 17614 59278 17666 59330
rect 17666 59278 17668 59330
rect 17612 59276 17668 59278
rect 18060 59836 18116 59892
rect 19516 62354 19572 62356
rect 19516 62302 19518 62354
rect 19518 62302 19570 62354
rect 19570 62302 19572 62354
rect 19516 62300 19572 62302
rect 20412 62188 20468 62244
rect 20860 62242 20916 62244
rect 20860 62190 20862 62242
rect 20862 62190 20914 62242
rect 20914 62190 20916 62242
rect 20860 62188 20916 62190
rect 18844 60396 18900 60452
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 20188 60396 20244 60452
rect 18172 59724 18228 59780
rect 19852 59724 19908 59780
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 18060 59276 18116 59332
rect 18060 59106 18116 59108
rect 18060 59054 18062 59106
rect 18062 59054 18114 59106
rect 18114 59054 18116 59106
rect 18060 59052 18116 59054
rect 20300 58940 20356 58996
rect 21756 60620 21812 60676
rect 16492 58156 16548 58212
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19740 57820 19796 57876
rect 16604 57708 16660 57764
rect 16492 52444 16548 52500
rect 15932 52162 15988 52164
rect 15932 52110 15934 52162
rect 15934 52110 15986 52162
rect 15986 52110 15988 52162
rect 15932 52108 15988 52110
rect 19404 57650 19460 57652
rect 19404 57598 19406 57650
rect 19406 57598 19458 57650
rect 19458 57598 19460 57650
rect 19404 57596 19460 57598
rect 19068 57484 19124 57540
rect 20300 57820 20356 57876
rect 19852 56812 19908 56868
rect 16940 55020 16996 55076
rect 16716 54402 16772 54404
rect 16716 54350 16718 54402
rect 16718 54350 16770 54402
rect 16770 54350 16772 54402
rect 16716 54348 16772 54350
rect 15260 47516 15316 47572
rect 14700 47068 14756 47124
rect 14476 46674 14532 46676
rect 14476 46622 14478 46674
rect 14478 46622 14530 46674
rect 14530 46622 14532 46674
rect 14476 46620 14532 46622
rect 14476 45164 14532 45220
rect 14812 45666 14868 45668
rect 14812 45614 14814 45666
rect 14814 45614 14866 45666
rect 14866 45614 14868 45666
rect 14812 45612 14868 45614
rect 14812 45164 14868 45220
rect 15036 45052 15092 45108
rect 16268 49196 16324 49252
rect 16716 49084 16772 49140
rect 16492 47516 16548 47572
rect 16604 48076 16660 48132
rect 16380 47458 16436 47460
rect 16380 47406 16382 47458
rect 16382 47406 16434 47458
rect 16434 47406 16436 47458
rect 16380 47404 16436 47406
rect 15820 47068 15876 47124
rect 15932 46562 15988 46564
rect 15932 46510 15934 46562
rect 15934 46510 15986 46562
rect 15986 46510 15988 46562
rect 15932 46508 15988 46510
rect 15484 45778 15540 45780
rect 15484 45726 15486 45778
rect 15486 45726 15538 45778
rect 15538 45726 15540 45778
rect 15484 45724 15540 45726
rect 15372 45612 15428 45668
rect 15820 45890 15876 45892
rect 15820 45838 15822 45890
rect 15822 45838 15874 45890
rect 15874 45838 15876 45890
rect 15820 45836 15876 45838
rect 15820 45612 15876 45668
rect 15820 45106 15876 45108
rect 15820 45054 15822 45106
rect 15822 45054 15874 45106
rect 15874 45054 15876 45106
rect 15820 45052 15876 45054
rect 15372 44380 15428 44436
rect 15820 44380 15876 44436
rect 14700 42812 14756 42868
rect 14700 42028 14756 42084
rect 14140 41804 14196 41860
rect 14588 41858 14644 41860
rect 14588 41806 14590 41858
rect 14590 41806 14642 41858
rect 14642 41806 14644 41858
rect 14588 41804 14644 41806
rect 14252 40572 14308 40628
rect 14476 41692 14532 41748
rect 14364 40514 14420 40516
rect 14364 40462 14366 40514
rect 14366 40462 14418 40514
rect 14418 40462 14420 40514
rect 14364 40460 14420 40462
rect 14588 40962 14644 40964
rect 14588 40910 14590 40962
rect 14590 40910 14642 40962
rect 14642 40910 14644 40962
rect 14588 40908 14644 40910
rect 14252 40402 14308 40404
rect 14252 40350 14254 40402
rect 14254 40350 14306 40402
rect 14306 40350 14308 40402
rect 14252 40348 14308 40350
rect 14364 40236 14420 40292
rect 12236 38780 12292 38836
rect 12684 38892 12740 38948
rect 12460 38834 12516 38836
rect 12460 38782 12462 38834
rect 12462 38782 12514 38834
rect 12514 38782 12516 38834
rect 12460 38780 12516 38782
rect 12348 38556 12404 38612
rect 11900 37266 11956 37268
rect 11900 37214 11902 37266
rect 11902 37214 11954 37266
rect 11954 37214 11956 37266
rect 11900 37212 11956 37214
rect 12460 37378 12516 37380
rect 12460 37326 12462 37378
rect 12462 37326 12514 37378
rect 12514 37326 12516 37378
rect 12460 37324 12516 37326
rect 12796 38668 12852 38724
rect 13468 38668 13524 38724
rect 14252 39564 14308 39620
rect 14140 38892 14196 38948
rect 14028 37660 14084 37716
rect 15036 42700 15092 42756
rect 15484 43538 15540 43540
rect 15484 43486 15486 43538
rect 15486 43486 15538 43538
rect 15538 43486 15540 43538
rect 15484 43484 15540 43486
rect 16156 44434 16212 44436
rect 16156 44382 16158 44434
rect 16158 44382 16210 44434
rect 16210 44382 16212 44434
rect 16156 44380 16212 44382
rect 16380 43820 16436 43876
rect 16156 43426 16212 43428
rect 16156 43374 16158 43426
rect 16158 43374 16210 43426
rect 16210 43374 16212 43426
rect 16156 43372 16212 43374
rect 16156 42924 16212 42980
rect 15484 42700 15540 42756
rect 15148 42028 15204 42084
rect 15260 41746 15316 41748
rect 15260 41694 15262 41746
rect 15262 41694 15314 41746
rect 15314 41694 15316 41746
rect 15260 41692 15316 41694
rect 15596 42082 15652 42084
rect 15596 42030 15598 42082
rect 15598 42030 15650 42082
rect 15650 42030 15652 42082
rect 15596 42028 15652 42030
rect 15596 41804 15652 41860
rect 15372 41580 15428 41636
rect 14924 40572 14980 40628
rect 14812 40402 14868 40404
rect 14812 40350 14814 40402
rect 14814 40350 14866 40402
rect 14866 40350 14868 40402
rect 14812 40348 14868 40350
rect 14588 39900 14644 39956
rect 14812 39900 14868 39956
rect 15148 40572 15204 40628
rect 15820 42530 15876 42532
rect 15820 42478 15822 42530
rect 15822 42478 15874 42530
rect 15874 42478 15876 42530
rect 15820 42476 15876 42478
rect 15708 40908 15764 40964
rect 15148 39564 15204 39620
rect 14700 37938 14756 37940
rect 14700 37886 14702 37938
rect 14702 37886 14754 37938
rect 14754 37886 14756 37938
rect 14700 37884 14756 37886
rect 12236 36316 12292 36372
rect 12796 36482 12852 36484
rect 12796 36430 12798 36482
rect 12798 36430 12850 36482
rect 12850 36430 12852 36482
rect 12796 36428 12852 36430
rect 12684 36258 12740 36260
rect 12684 36206 12686 36258
rect 12686 36206 12738 36258
rect 12738 36206 12740 36258
rect 12684 36204 12740 36206
rect 11340 35420 11396 35476
rect 12572 35698 12628 35700
rect 12572 35646 12574 35698
rect 12574 35646 12626 35698
rect 12626 35646 12628 35698
rect 12572 35644 12628 35646
rect 12348 35308 12404 35364
rect 10332 32562 10388 32564
rect 10332 32510 10334 32562
rect 10334 32510 10386 32562
rect 10386 32510 10388 32562
rect 10332 32508 10388 32510
rect 9772 31836 9828 31892
rect 10444 32060 10500 32116
rect 8876 29932 8932 29988
rect 9660 29986 9716 29988
rect 9660 29934 9662 29986
rect 9662 29934 9714 29986
rect 9714 29934 9716 29986
rect 9660 29932 9716 29934
rect 9324 29820 9380 29876
rect 9100 29484 9156 29540
rect 8652 27580 8708 27636
rect 7420 27074 7476 27076
rect 7420 27022 7422 27074
rect 7422 27022 7474 27074
rect 7474 27022 7476 27074
rect 7420 27020 7476 27022
rect 9772 29538 9828 29540
rect 9772 29486 9774 29538
rect 9774 29486 9826 29538
rect 9826 29486 9828 29538
rect 9772 29484 9828 29486
rect 9548 29426 9604 29428
rect 9548 29374 9550 29426
rect 9550 29374 9602 29426
rect 9602 29374 9604 29426
rect 9548 29372 9604 29374
rect 9660 28588 9716 28644
rect 9548 28140 9604 28196
rect 9548 27804 9604 27860
rect 7084 26796 7140 26852
rect 7868 26796 7924 26852
rect 7644 25506 7700 25508
rect 7644 25454 7646 25506
rect 7646 25454 7698 25506
rect 7698 25454 7700 25506
rect 7644 25452 7700 25454
rect 8204 26124 8260 26180
rect 8428 25228 8484 25284
rect 9324 25394 9380 25396
rect 9324 25342 9326 25394
rect 9326 25342 9378 25394
rect 9378 25342 9380 25394
rect 9324 25340 9380 25342
rect 8876 25116 8932 25172
rect 9884 27804 9940 27860
rect 10108 30098 10164 30100
rect 10108 30046 10110 30098
rect 10110 30046 10162 30098
rect 10162 30046 10164 30098
rect 10108 30044 10164 30046
rect 10556 30044 10612 30100
rect 12460 33404 12516 33460
rect 11452 33180 11508 33236
rect 11564 32396 11620 32452
rect 11900 32786 11956 32788
rect 11900 32734 11902 32786
rect 11902 32734 11954 32786
rect 11954 32734 11956 32786
rect 11900 32732 11956 32734
rect 12236 32396 12292 32452
rect 12012 32172 12068 32228
rect 11340 30828 11396 30884
rect 10892 29820 10948 29876
rect 10780 29708 10836 29764
rect 10780 29372 10836 29428
rect 11116 29484 11172 29540
rect 11004 28140 11060 28196
rect 11004 27916 11060 27972
rect 10108 27580 10164 27636
rect 11004 27356 11060 27412
rect 10668 26796 10724 26852
rect 11564 29820 11620 29876
rect 11340 29596 11396 29652
rect 11452 29484 11508 29540
rect 13468 36482 13524 36484
rect 13468 36430 13470 36482
rect 13470 36430 13522 36482
rect 13522 36430 13524 36482
rect 13468 36428 13524 36430
rect 13580 35868 13636 35924
rect 13580 35586 13636 35588
rect 13580 35534 13582 35586
rect 13582 35534 13634 35586
rect 13634 35534 13636 35586
rect 13580 35532 13636 35534
rect 12796 35084 12852 35140
rect 12796 33292 12852 33348
rect 13020 33516 13076 33572
rect 12796 32732 12852 32788
rect 12796 31836 12852 31892
rect 13468 33180 13524 33236
rect 12908 30940 12964 30996
rect 12348 29596 12404 29652
rect 12124 29260 12180 29316
rect 12796 29260 12852 29316
rect 12348 29036 12404 29092
rect 11564 27244 11620 27300
rect 11228 26796 11284 26852
rect 12012 27132 12068 27188
rect 11788 26796 11844 26852
rect 10556 26178 10612 26180
rect 10556 26126 10558 26178
rect 10558 26126 10610 26178
rect 10610 26126 10612 26178
rect 10556 26124 10612 26126
rect 10444 25228 10500 25284
rect 13804 35532 13860 35588
rect 13916 33516 13972 33572
rect 15036 37772 15092 37828
rect 14924 37266 14980 37268
rect 14924 37214 14926 37266
rect 14926 37214 14978 37266
rect 14978 37214 14980 37266
rect 14924 37212 14980 37214
rect 16380 42866 16436 42868
rect 16380 42814 16382 42866
rect 16382 42814 16434 42866
rect 16434 42814 16436 42866
rect 16380 42812 16436 42814
rect 16492 42754 16548 42756
rect 16492 42702 16494 42754
rect 16494 42702 16546 42754
rect 16546 42702 16548 42754
rect 16492 42700 16548 42702
rect 16828 42028 16884 42084
rect 16716 41970 16772 41972
rect 16716 41918 16718 41970
rect 16718 41918 16770 41970
rect 16770 41918 16772 41970
rect 16716 41916 16772 41918
rect 15372 40290 15428 40292
rect 15372 40238 15374 40290
rect 15374 40238 15426 40290
rect 15426 40238 15428 40290
rect 15372 40236 15428 40238
rect 15932 39618 15988 39620
rect 15932 39566 15934 39618
rect 15934 39566 15986 39618
rect 15986 39566 15988 39618
rect 15932 39564 15988 39566
rect 16380 41804 16436 41860
rect 16492 41692 16548 41748
rect 16604 40178 16660 40180
rect 16604 40126 16606 40178
rect 16606 40126 16658 40178
rect 16658 40126 16660 40178
rect 16604 40124 16660 40126
rect 15260 38892 15316 38948
rect 15820 39004 15876 39060
rect 15372 38610 15428 38612
rect 15372 38558 15374 38610
rect 15374 38558 15426 38610
rect 15426 38558 15428 38610
rect 15372 38556 15428 38558
rect 15372 38332 15428 38388
rect 15708 37996 15764 38052
rect 15932 37548 15988 37604
rect 16492 38332 16548 38388
rect 16492 38108 16548 38164
rect 15148 37042 15204 37044
rect 15148 36990 15150 37042
rect 15150 36990 15202 37042
rect 15202 36990 15204 37042
rect 15148 36988 15204 36990
rect 15708 35644 15764 35700
rect 14364 35532 14420 35588
rect 14252 35084 14308 35140
rect 15148 34636 15204 34692
rect 15820 34636 15876 34692
rect 15484 33964 15540 34020
rect 15148 33516 15204 33572
rect 14588 33458 14644 33460
rect 14588 33406 14590 33458
rect 14590 33406 14642 33458
rect 14642 33406 14644 33458
rect 14588 33404 14644 33406
rect 14812 33346 14868 33348
rect 14812 33294 14814 33346
rect 14814 33294 14866 33346
rect 14866 33294 14868 33346
rect 14812 33292 14868 33294
rect 13580 31724 13636 31780
rect 13692 32284 13748 32340
rect 13916 32620 13972 32676
rect 14028 32396 14084 32452
rect 13132 29372 13188 29428
rect 13580 31276 13636 31332
rect 13468 29484 13524 29540
rect 13468 29202 13524 29204
rect 13468 29150 13470 29202
rect 13470 29150 13522 29202
rect 13522 29150 13524 29202
rect 13468 29148 13524 29150
rect 13580 29036 13636 29092
rect 15820 33404 15876 33460
rect 14588 32674 14644 32676
rect 14588 32622 14590 32674
rect 14590 32622 14642 32674
rect 14642 32622 14644 32674
rect 14588 32620 14644 32622
rect 14812 32338 14868 32340
rect 14812 32286 14814 32338
rect 14814 32286 14866 32338
rect 14866 32286 14868 32338
rect 14812 32284 14868 32286
rect 15372 32060 15428 32116
rect 14252 31890 14308 31892
rect 14252 31838 14254 31890
rect 14254 31838 14306 31890
rect 14306 31838 14308 31890
rect 14252 31836 14308 31838
rect 14140 31724 14196 31780
rect 13916 30994 13972 30996
rect 13916 30942 13918 30994
rect 13918 30942 13970 30994
rect 13970 30942 13972 30994
rect 13916 30940 13972 30942
rect 14476 31276 14532 31332
rect 12348 27244 12404 27300
rect 14028 28812 14084 28868
rect 13356 27692 13412 27748
rect 13132 27244 13188 27300
rect 12348 27020 12404 27076
rect 12236 26908 12292 26964
rect 14028 28588 14084 28644
rect 13580 27020 13636 27076
rect 13692 28530 13748 28532
rect 13692 28478 13694 28530
rect 13694 28478 13746 28530
rect 13746 28478 13748 28530
rect 13692 28476 13748 28478
rect 13244 26796 13300 26852
rect 14028 28418 14084 28420
rect 14028 28366 14030 28418
rect 14030 28366 14082 28418
rect 14082 28366 14084 28418
rect 14028 28364 14084 28366
rect 13916 28252 13972 28308
rect 14252 30156 14308 30212
rect 17836 53788 17892 53844
rect 17948 53452 18004 53508
rect 17500 52946 17556 52948
rect 17500 52894 17502 52946
rect 17502 52894 17554 52946
rect 17554 52894 17556 52946
rect 17500 52892 17556 52894
rect 17500 50876 17556 50932
rect 17388 48914 17444 48916
rect 17388 48862 17390 48914
rect 17390 48862 17442 48914
rect 17442 48862 17444 48914
rect 17388 48860 17444 48862
rect 17052 45890 17108 45892
rect 17052 45838 17054 45890
rect 17054 45838 17106 45890
rect 17106 45838 17108 45890
rect 17052 45836 17108 45838
rect 17612 47458 17668 47460
rect 17612 47406 17614 47458
rect 17614 47406 17666 47458
rect 17666 47406 17668 47458
rect 17612 47404 17668 47406
rect 17948 47068 18004 47124
rect 18284 54514 18340 54516
rect 18284 54462 18286 54514
rect 18286 54462 18338 54514
rect 18338 54462 18340 54514
rect 18284 54460 18340 54462
rect 19068 54460 19124 54516
rect 18732 53842 18788 53844
rect 18732 53790 18734 53842
rect 18734 53790 18786 53842
rect 18786 53790 18788 53842
rect 18732 53788 18788 53790
rect 20300 57650 20356 57652
rect 20300 57598 20302 57650
rect 20302 57598 20354 57650
rect 20354 57598 20356 57650
rect 20300 57596 20356 57598
rect 21084 58940 21140 58996
rect 20748 58268 20804 58324
rect 20748 57650 20804 57652
rect 20748 57598 20750 57650
rect 20750 57598 20802 57650
rect 20802 57598 20804 57650
rect 20748 57596 20804 57598
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20748 56866 20804 56868
rect 20748 56814 20750 56866
rect 20750 56814 20802 56866
rect 20802 56814 20804 56866
rect 20748 56812 20804 56814
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19628 54460 19684 54516
rect 20524 53788 20580 53844
rect 19852 53730 19908 53732
rect 19852 53678 19854 53730
rect 19854 53678 19906 53730
rect 19906 53678 19908 53730
rect 19852 53676 19908 53678
rect 19404 53564 19460 53620
rect 18844 53506 18900 53508
rect 18844 53454 18846 53506
rect 18846 53454 18898 53506
rect 18898 53454 18900 53506
rect 18844 53452 18900 53454
rect 19628 53506 19684 53508
rect 19628 53454 19630 53506
rect 19630 53454 19682 53506
rect 19682 53454 19684 53506
rect 19628 53452 19684 53454
rect 20076 53506 20132 53508
rect 20076 53454 20078 53506
rect 20078 53454 20130 53506
rect 20130 53454 20132 53506
rect 20076 53452 20132 53454
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19628 52556 19684 52612
rect 20300 52834 20356 52836
rect 20300 52782 20302 52834
rect 20302 52782 20354 52834
rect 20354 52782 20356 52834
rect 20300 52780 20356 52782
rect 19180 52162 19236 52164
rect 19180 52110 19182 52162
rect 19182 52110 19234 52162
rect 19234 52110 19236 52162
rect 19180 52108 19236 52110
rect 20636 53618 20692 53620
rect 20636 53566 20638 53618
rect 20638 53566 20690 53618
rect 20690 53566 20692 53618
rect 20636 53564 20692 53566
rect 20636 53228 20692 53284
rect 20636 52946 20692 52948
rect 20636 52894 20638 52946
rect 20638 52894 20690 52946
rect 20690 52894 20692 52946
rect 20636 52892 20692 52894
rect 20524 52780 20580 52836
rect 20524 52556 20580 52612
rect 20300 52108 20356 52164
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20748 52386 20804 52388
rect 20748 52334 20750 52386
rect 20750 52334 20802 52386
rect 20802 52334 20804 52386
rect 20748 52332 20804 52334
rect 19292 49922 19348 49924
rect 19292 49870 19294 49922
rect 19294 49870 19346 49922
rect 19346 49870 19348 49922
rect 19292 49868 19348 49870
rect 19180 49644 19236 49700
rect 19404 49756 19460 49812
rect 19068 49084 19124 49140
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20300 49868 20356 49924
rect 19740 49644 19796 49700
rect 18172 47458 18228 47460
rect 18172 47406 18174 47458
rect 18174 47406 18226 47458
rect 18226 47406 18228 47458
rect 18172 47404 18228 47406
rect 19068 47404 19124 47460
rect 18284 47180 18340 47236
rect 18620 47068 18676 47124
rect 18172 46114 18228 46116
rect 18172 46062 18174 46114
rect 18174 46062 18226 46114
rect 18226 46062 18228 46114
rect 18172 46060 18228 46062
rect 20188 48914 20244 48916
rect 20188 48862 20190 48914
rect 20190 48862 20242 48914
rect 20242 48862 20244 48914
rect 20188 48860 20244 48862
rect 20076 48748 20132 48804
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20524 49698 20580 49700
rect 20524 49646 20526 49698
rect 20526 49646 20578 49698
rect 20578 49646 20580 49698
rect 20524 49644 20580 49646
rect 20636 48914 20692 48916
rect 20636 48862 20638 48914
rect 20638 48862 20690 48914
rect 20690 48862 20692 48914
rect 20636 48860 20692 48862
rect 20412 48636 20468 48692
rect 20524 48748 20580 48804
rect 20972 48130 21028 48132
rect 20972 48078 20974 48130
rect 20974 48078 21026 48130
rect 21026 48078 21028 48130
rect 20972 48076 21028 48078
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19404 46674 19460 46676
rect 19404 46622 19406 46674
rect 19406 46622 19458 46674
rect 19458 46622 19460 46674
rect 19404 46620 19460 46622
rect 19740 46450 19796 46452
rect 19740 46398 19742 46450
rect 19742 46398 19794 46450
rect 19794 46398 19796 46450
rect 19740 46396 19796 46398
rect 19292 45948 19348 46004
rect 17836 43820 17892 43876
rect 18060 43708 18116 43764
rect 17164 43372 17220 43428
rect 17276 41692 17332 41748
rect 17388 40460 17444 40516
rect 16940 40236 16996 40292
rect 17276 40348 17332 40404
rect 16716 39004 16772 39060
rect 17052 37884 17108 37940
rect 16828 37660 16884 37716
rect 16604 37212 16660 37268
rect 16716 37436 16772 37492
rect 16044 35586 16100 35588
rect 16044 35534 16046 35586
rect 16046 35534 16098 35586
rect 16098 35534 16100 35586
rect 16044 35532 16100 35534
rect 16268 34636 16324 34692
rect 18732 44940 18788 44996
rect 20188 46172 20244 46228
rect 22652 61292 22708 61348
rect 22652 60786 22708 60788
rect 22652 60734 22654 60786
rect 22654 60734 22706 60786
rect 22706 60734 22708 60786
rect 22652 60732 22708 60734
rect 23212 60674 23268 60676
rect 23212 60622 23214 60674
rect 23214 60622 23266 60674
rect 23266 60622 23268 60674
rect 23212 60620 23268 60622
rect 23660 63868 23716 63924
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 39004 66444 39060 66500
rect 40796 66498 40852 66500
rect 40796 66446 40798 66498
rect 40798 66446 40850 66498
rect 40850 66446 40852 66498
rect 40796 66444 40852 66446
rect 33852 65436 33908 65492
rect 30268 64876 30324 64932
rect 25452 64428 25508 64484
rect 27804 64652 27860 64708
rect 26684 64204 26740 64260
rect 26348 63644 26404 63700
rect 24780 63196 24836 63252
rect 26236 63250 26292 63252
rect 26236 63198 26238 63250
rect 26238 63198 26290 63250
rect 26290 63198 26292 63250
rect 26236 63196 26292 63198
rect 26124 62860 26180 62916
rect 25900 62076 25956 62132
rect 23548 60620 23604 60676
rect 23996 59836 24052 59892
rect 21308 55468 21364 55524
rect 21196 53788 21252 53844
rect 21308 53228 21364 53284
rect 26684 63138 26740 63140
rect 26684 63086 26686 63138
rect 26686 63086 26738 63138
rect 26738 63086 26740 63138
rect 26684 63084 26740 63086
rect 26460 63026 26516 63028
rect 26460 62974 26462 63026
rect 26462 62974 26514 63026
rect 26514 62974 26516 63026
rect 26460 62972 26516 62974
rect 27468 64204 27524 64260
rect 28140 64204 28196 64260
rect 27244 63644 27300 63700
rect 27132 63138 27188 63140
rect 27132 63086 27134 63138
rect 27134 63086 27186 63138
rect 27186 63086 27188 63138
rect 27132 63084 27188 63086
rect 27020 62914 27076 62916
rect 27020 62862 27022 62914
rect 27022 62862 27074 62914
rect 27074 62862 27076 62914
rect 27020 62860 27076 62862
rect 27244 62972 27300 63028
rect 27580 62860 27636 62916
rect 27244 62300 27300 62356
rect 28252 63644 28308 63700
rect 29148 64652 29204 64708
rect 28364 62300 28420 62356
rect 28476 62860 28532 62916
rect 27692 62076 27748 62132
rect 25116 61068 25172 61124
rect 24668 59500 24724 59556
rect 25564 61346 25620 61348
rect 25564 61294 25566 61346
rect 25566 61294 25618 61346
rect 25618 61294 25620 61346
rect 25564 61292 25620 61294
rect 25452 61010 25508 61012
rect 25452 60958 25454 61010
rect 25454 60958 25506 61010
rect 25506 60958 25508 61010
rect 25452 60956 25508 60958
rect 25452 60732 25508 60788
rect 26012 61010 26068 61012
rect 26012 60958 26014 61010
rect 26014 60958 26066 61010
rect 26066 60958 26068 61010
rect 26012 60956 26068 60958
rect 25900 60786 25956 60788
rect 25900 60734 25902 60786
rect 25902 60734 25954 60786
rect 25954 60734 25956 60786
rect 25900 60732 25956 60734
rect 25676 60620 25732 60676
rect 25116 59052 25172 59108
rect 24668 57820 24724 57876
rect 25676 58434 25732 58436
rect 25676 58382 25678 58434
rect 25678 58382 25730 58434
rect 25730 58382 25732 58434
rect 25676 58380 25732 58382
rect 28140 61180 28196 61236
rect 27132 60786 27188 60788
rect 27132 60734 27134 60786
rect 27134 60734 27186 60786
rect 27186 60734 27188 60786
rect 27132 60732 27188 60734
rect 26572 59890 26628 59892
rect 26572 59838 26574 59890
rect 26574 59838 26626 59890
rect 26626 59838 26628 59890
rect 26572 59836 26628 59838
rect 27804 60898 27860 60900
rect 27804 60846 27806 60898
rect 27806 60846 27858 60898
rect 27858 60846 27860 60898
rect 27804 60844 27860 60846
rect 27244 60508 27300 60564
rect 27916 60786 27972 60788
rect 27916 60734 27918 60786
rect 27918 60734 27970 60786
rect 27970 60734 27972 60786
rect 27916 60732 27972 60734
rect 27692 60620 27748 60676
rect 28028 60508 28084 60564
rect 27468 59948 27524 60004
rect 26684 58434 26740 58436
rect 26684 58382 26686 58434
rect 26686 58382 26738 58434
rect 26738 58382 26740 58434
rect 26684 58380 26740 58382
rect 26012 58268 26068 58324
rect 22988 56140 23044 56196
rect 23660 56140 23716 56196
rect 23660 55804 23716 55860
rect 22316 53842 22372 53844
rect 22316 53790 22318 53842
rect 22318 53790 22370 53842
rect 22370 53790 22372 53842
rect 22316 53788 22372 53790
rect 26236 58156 26292 58212
rect 25676 57036 25732 57092
rect 24108 55916 24164 55972
rect 23324 54012 23380 54068
rect 24444 55804 24500 55860
rect 25228 55468 25284 55524
rect 24780 54012 24836 54068
rect 23100 53618 23156 53620
rect 23100 53566 23102 53618
rect 23102 53566 23154 53618
rect 23154 53566 23156 53618
rect 23100 53564 23156 53566
rect 23548 53564 23604 53620
rect 23212 53506 23268 53508
rect 23212 53454 23214 53506
rect 23214 53454 23266 53506
rect 23266 53454 23268 53506
rect 23212 53452 23268 53454
rect 23100 52892 23156 52948
rect 23884 53452 23940 53508
rect 24332 53618 24388 53620
rect 24332 53566 24334 53618
rect 24334 53566 24386 53618
rect 24386 53566 24388 53618
rect 24332 53564 24388 53566
rect 24220 52946 24276 52948
rect 24220 52894 24222 52946
rect 24222 52894 24274 52946
rect 24274 52894 24276 52946
rect 24220 52892 24276 52894
rect 23100 52332 23156 52388
rect 24668 53170 24724 53172
rect 24668 53118 24670 53170
rect 24670 53118 24722 53170
rect 24722 53118 24724 53170
rect 24668 53116 24724 53118
rect 25340 53170 25396 53172
rect 25340 53118 25342 53170
rect 25342 53118 25394 53170
rect 25394 53118 25396 53170
rect 25340 53116 25396 53118
rect 22428 51436 22484 51492
rect 23772 51436 23828 51492
rect 21980 49980 22036 50036
rect 21420 49810 21476 49812
rect 21420 49758 21422 49810
rect 21422 49758 21474 49810
rect 21474 49758 21476 49810
rect 21420 49756 21476 49758
rect 21420 48914 21476 48916
rect 21420 48862 21422 48914
rect 21422 48862 21474 48914
rect 21474 48862 21476 48914
rect 21420 48860 21476 48862
rect 21308 48802 21364 48804
rect 21308 48750 21310 48802
rect 21310 48750 21362 48802
rect 21362 48750 21364 48802
rect 21308 48748 21364 48750
rect 21532 48636 21588 48692
rect 22540 49138 22596 49140
rect 22540 49086 22542 49138
rect 22542 49086 22594 49138
rect 22594 49086 22596 49138
rect 22540 49084 22596 49086
rect 22988 49084 23044 49140
rect 23660 48748 23716 48804
rect 21980 48076 22036 48132
rect 21532 47628 21588 47684
rect 23436 48076 23492 48132
rect 22652 47682 22708 47684
rect 22652 47630 22654 47682
rect 22654 47630 22706 47682
rect 22706 47630 22708 47682
rect 22652 47628 22708 47630
rect 23100 47570 23156 47572
rect 23100 47518 23102 47570
rect 23102 47518 23154 47570
rect 23154 47518 23156 47570
rect 23100 47516 23156 47518
rect 22988 46284 23044 46340
rect 21084 46172 21140 46228
rect 20748 45666 20804 45668
rect 20748 45614 20750 45666
rect 20750 45614 20802 45666
rect 20802 45614 20804 45666
rect 20748 45612 20804 45614
rect 21420 45666 21476 45668
rect 21420 45614 21422 45666
rect 21422 45614 21474 45666
rect 21474 45614 21476 45666
rect 21420 45612 21476 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 22316 45330 22372 45332
rect 22316 45278 22318 45330
rect 22318 45278 22370 45330
rect 22370 45278 22372 45330
rect 22316 45276 22372 45278
rect 21644 45164 21700 45220
rect 20972 44994 21028 44996
rect 20972 44942 20974 44994
rect 20974 44942 21026 44994
rect 21026 44942 21028 44994
rect 20972 44940 21028 44942
rect 18620 43596 18676 43652
rect 21644 44268 21700 44324
rect 22204 45218 22260 45220
rect 22204 45166 22206 45218
rect 22206 45166 22258 45218
rect 22258 45166 22260 45218
rect 22204 45164 22260 45166
rect 23324 45276 23380 45332
rect 21756 45052 21812 45108
rect 22428 45106 22484 45108
rect 22428 45054 22430 45106
rect 22430 45054 22482 45106
rect 22482 45054 22484 45106
rect 22428 45052 22484 45054
rect 22204 44828 22260 44884
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19068 43538 19124 43540
rect 19068 43486 19070 43538
rect 19070 43486 19122 43538
rect 19122 43486 19124 43538
rect 19068 43484 19124 43486
rect 20188 43708 20244 43764
rect 19740 43426 19796 43428
rect 19740 43374 19742 43426
rect 19742 43374 19794 43426
rect 19794 43374 19796 43426
rect 19740 43372 19796 43374
rect 18396 42924 18452 42980
rect 21196 43596 21252 43652
rect 20860 43484 20916 43540
rect 20300 42924 20356 42980
rect 18060 41468 18116 41524
rect 17724 39730 17780 39732
rect 17724 39678 17726 39730
rect 17726 39678 17778 39730
rect 17778 39678 17780 39730
rect 17724 39676 17780 39678
rect 17948 40348 18004 40404
rect 18284 40460 18340 40516
rect 17612 38050 17668 38052
rect 17612 37998 17614 38050
rect 17614 37998 17666 38050
rect 17666 37998 17668 38050
rect 17612 37996 17668 37998
rect 17500 37660 17556 37716
rect 17948 38162 18004 38164
rect 17948 38110 17950 38162
rect 17950 38110 18002 38162
rect 18002 38110 18004 38162
rect 17948 38108 18004 38110
rect 17724 37212 17780 37268
rect 18284 36482 18340 36484
rect 18284 36430 18286 36482
rect 18286 36430 18338 36482
rect 18338 36430 18340 36482
rect 18284 36428 18340 36430
rect 18396 41244 18452 41300
rect 18396 37660 18452 37716
rect 17388 35644 17444 35700
rect 17052 35420 17108 35476
rect 16716 33404 16772 33460
rect 16716 33234 16772 33236
rect 16716 33182 16718 33234
rect 16718 33182 16770 33234
rect 16770 33182 16772 33234
rect 16716 33180 16772 33182
rect 16828 32732 16884 32788
rect 15036 31554 15092 31556
rect 15036 31502 15038 31554
rect 15038 31502 15090 31554
rect 15090 31502 15092 31554
rect 15036 31500 15092 31502
rect 15484 31500 15540 31556
rect 15148 29426 15204 29428
rect 15148 29374 15150 29426
rect 15150 29374 15202 29426
rect 15202 29374 15204 29426
rect 15148 29372 15204 29374
rect 15708 30882 15764 30884
rect 15708 30830 15710 30882
rect 15710 30830 15762 30882
rect 15762 30830 15764 30882
rect 15708 30828 15764 30830
rect 15820 29932 15876 29988
rect 15484 29372 15540 29428
rect 15596 29260 15652 29316
rect 14812 29036 14868 29092
rect 15372 29148 15428 29204
rect 14924 28754 14980 28756
rect 14924 28702 14926 28754
rect 14926 28702 14978 28754
rect 14978 28702 14980 28754
rect 14924 28700 14980 28702
rect 14364 28140 14420 28196
rect 13916 27186 13972 27188
rect 13916 27134 13918 27186
rect 13918 27134 13970 27186
rect 13970 27134 13972 27186
rect 13916 27132 13972 27134
rect 9660 25116 9716 25172
rect 10220 25116 10276 25172
rect 12796 25282 12852 25284
rect 12796 25230 12798 25282
rect 12798 25230 12850 25282
rect 12850 25230 12852 25282
rect 12796 25228 12852 25230
rect 12460 24780 12516 24836
rect 10892 24610 10948 24612
rect 10892 24558 10894 24610
rect 10894 24558 10946 24610
rect 10946 24558 10948 24610
rect 10892 24556 10948 24558
rect 13916 25340 13972 25396
rect 14364 26962 14420 26964
rect 14364 26910 14366 26962
rect 14366 26910 14418 26962
rect 14418 26910 14420 26962
rect 14364 26908 14420 26910
rect 14812 28588 14868 28644
rect 15820 28754 15876 28756
rect 15820 28702 15822 28754
rect 15822 28702 15874 28754
rect 15874 28702 15876 28754
rect 15820 28700 15876 28702
rect 15708 28364 15764 28420
rect 15260 27970 15316 27972
rect 15260 27918 15262 27970
rect 15262 27918 15314 27970
rect 15314 27918 15316 27970
rect 15260 27916 15316 27918
rect 14700 27804 14756 27860
rect 15708 27692 15764 27748
rect 15148 27132 15204 27188
rect 14700 27074 14756 27076
rect 14700 27022 14702 27074
rect 14702 27022 14754 27074
rect 14754 27022 14756 27074
rect 14700 27020 14756 27022
rect 15260 26908 15316 26964
rect 15820 27580 15876 27636
rect 15708 26908 15764 26964
rect 15932 27020 15988 27076
rect 14588 26460 14644 26516
rect 13580 25116 13636 25172
rect 13804 24668 13860 24724
rect 14924 26460 14980 26516
rect 15596 26514 15652 26516
rect 15596 26462 15598 26514
rect 15598 26462 15650 26514
rect 15650 26462 15652 26514
rect 15596 26460 15652 26462
rect 17948 34636 18004 34692
rect 17612 32786 17668 32788
rect 17612 32734 17614 32786
rect 17614 32734 17666 32786
rect 17666 32734 17668 32786
rect 17612 32732 17668 32734
rect 18172 32732 18228 32788
rect 17388 31836 17444 31892
rect 16492 30098 16548 30100
rect 16492 30046 16494 30098
rect 16494 30046 16546 30098
rect 16546 30046 16548 30098
rect 16492 30044 16548 30046
rect 17052 30098 17108 30100
rect 17052 30046 17054 30098
rect 17054 30046 17106 30098
rect 17106 30046 17108 30098
rect 17052 30044 17108 30046
rect 18284 31724 18340 31780
rect 16604 29986 16660 29988
rect 16604 29934 16606 29986
rect 16606 29934 16658 29986
rect 16658 29934 16660 29986
rect 16604 29932 16660 29934
rect 16380 29036 16436 29092
rect 16380 28812 16436 28868
rect 16828 29260 16884 29316
rect 17388 29260 17444 29316
rect 17836 29986 17892 29988
rect 17836 29934 17838 29986
rect 17838 29934 17890 29986
rect 17890 29934 17892 29986
rect 17836 29932 17892 29934
rect 17612 28812 17668 28868
rect 18172 28866 18228 28868
rect 18172 28814 18174 28866
rect 18174 28814 18226 28866
rect 18226 28814 18228 28866
rect 18172 28812 18228 28814
rect 17500 28530 17556 28532
rect 17500 28478 17502 28530
rect 17502 28478 17554 28530
rect 17554 28478 17556 28530
rect 17500 28476 17556 28478
rect 17052 28418 17108 28420
rect 17052 28366 17054 28418
rect 17054 28366 17106 28418
rect 17106 28366 17108 28418
rect 17052 28364 17108 28366
rect 15932 26514 15988 26516
rect 15932 26462 15934 26514
rect 15934 26462 15986 26514
rect 15986 26462 15988 26514
rect 15932 26460 15988 26462
rect 16604 26348 16660 26404
rect 14476 25004 14532 25060
rect 15036 25116 15092 25172
rect 15148 25004 15204 25060
rect 14252 24780 14308 24836
rect 14364 24610 14420 24612
rect 14364 24558 14366 24610
rect 14366 24558 14418 24610
rect 14418 24558 14420 24610
rect 14364 24556 14420 24558
rect 14588 24556 14644 24612
rect 15596 24610 15652 24612
rect 15596 24558 15598 24610
rect 15598 24558 15650 24610
rect 15650 24558 15652 24610
rect 15596 24556 15652 24558
rect 15820 25116 15876 25172
rect 15820 23660 15876 23716
rect 16604 25506 16660 25508
rect 16604 25454 16606 25506
rect 16606 25454 16658 25506
rect 16658 25454 16660 25506
rect 16604 25452 16660 25454
rect 16156 24946 16212 24948
rect 16156 24894 16158 24946
rect 16158 24894 16210 24946
rect 16210 24894 16212 24946
rect 16156 24892 16212 24894
rect 16828 26290 16884 26292
rect 16828 26238 16830 26290
rect 16830 26238 16882 26290
rect 16882 26238 16884 26290
rect 16828 26236 16884 26238
rect 17164 28028 17220 28084
rect 17612 27580 17668 27636
rect 17052 26348 17108 26404
rect 17388 26402 17444 26404
rect 17388 26350 17390 26402
rect 17390 26350 17442 26402
rect 17442 26350 17444 26402
rect 17388 26348 17444 26350
rect 16828 25340 16884 25396
rect 17388 25452 17444 25508
rect 18172 28588 18228 28644
rect 18284 28364 18340 28420
rect 18172 28082 18228 28084
rect 18172 28030 18174 28082
rect 18174 28030 18226 28082
rect 18226 28030 18228 28082
rect 18172 28028 18228 28030
rect 18060 26402 18116 26404
rect 18060 26350 18062 26402
rect 18062 26350 18114 26402
rect 18114 26350 18116 26402
rect 18060 26348 18116 26350
rect 17724 26290 17780 26292
rect 17724 26238 17726 26290
rect 17726 26238 17778 26290
rect 17778 26238 17780 26290
rect 17724 26236 17780 26238
rect 17724 25676 17780 25732
rect 16492 24668 16548 24724
rect 16380 24556 16436 24612
rect 19180 42028 19236 42084
rect 18732 41244 18788 41300
rect 19516 41356 19572 41412
rect 19180 41020 19236 41076
rect 19404 40908 19460 40964
rect 19404 40348 19460 40404
rect 18732 39676 18788 39732
rect 18844 40124 18900 40180
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19964 42140 20020 42196
rect 19964 41858 20020 41860
rect 19964 41806 19966 41858
rect 19966 41806 20018 41858
rect 20018 41806 20020 41858
rect 19964 41804 20020 41806
rect 20300 41916 20356 41972
rect 20188 41074 20244 41076
rect 20188 41022 20190 41074
rect 20190 41022 20242 41074
rect 20242 41022 20244 41074
rect 20188 41020 20244 41022
rect 19964 40908 20020 40964
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20748 42140 20804 42196
rect 20748 41692 20804 41748
rect 20636 41580 20692 41636
rect 20524 41244 20580 41300
rect 20300 40402 20356 40404
rect 20300 40350 20302 40402
rect 20302 40350 20354 40402
rect 20354 40350 20356 40402
rect 20300 40348 20356 40350
rect 20188 39618 20244 39620
rect 20188 39566 20190 39618
rect 20190 39566 20242 39618
rect 20242 39566 20244 39618
rect 20188 39564 20244 39566
rect 19628 39452 19684 39508
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19628 39058 19684 39060
rect 19628 39006 19630 39058
rect 19630 39006 19682 39058
rect 19682 39006 19684 39058
rect 19628 39004 19684 39006
rect 20412 40236 20468 40292
rect 20860 41580 20916 41636
rect 20636 39788 20692 39844
rect 20748 41356 20804 41412
rect 20300 38892 20356 38948
rect 19740 38668 19796 38724
rect 21084 42476 21140 42532
rect 22092 44322 22148 44324
rect 22092 44270 22094 44322
rect 22094 44270 22146 44322
rect 22146 44270 22148 44322
rect 22092 44268 22148 44270
rect 23100 44828 23156 44884
rect 23772 47964 23828 48020
rect 23660 47458 23716 47460
rect 23660 47406 23662 47458
rect 23662 47406 23714 47458
rect 23714 47406 23716 47458
rect 23660 47404 23716 47406
rect 25116 49084 25172 49140
rect 24444 48748 24500 48804
rect 24332 47516 24388 47572
rect 23660 47180 23716 47236
rect 24668 48018 24724 48020
rect 24668 47966 24670 48018
rect 24670 47966 24722 48018
rect 24722 47966 24724 48018
rect 24668 47964 24724 47966
rect 24556 47458 24612 47460
rect 24556 47406 24558 47458
rect 24558 47406 24610 47458
rect 24610 47406 24612 47458
rect 24556 47404 24612 47406
rect 24892 47180 24948 47236
rect 24332 47068 24388 47124
rect 23548 46674 23604 46676
rect 23548 46622 23550 46674
rect 23550 46622 23602 46674
rect 23602 46622 23604 46674
rect 23548 46620 23604 46622
rect 23660 46284 23716 46340
rect 23324 44156 23380 44212
rect 23212 43932 23268 43988
rect 22092 43484 22148 43540
rect 22316 43426 22372 43428
rect 22316 43374 22318 43426
rect 22318 43374 22370 43426
rect 22370 43374 22372 43426
rect 22316 43372 22372 43374
rect 21308 42642 21364 42644
rect 21308 42590 21310 42642
rect 21310 42590 21362 42642
rect 21362 42590 21364 42642
rect 21308 42588 21364 42590
rect 21532 42476 21588 42532
rect 21308 41468 21364 41524
rect 21196 41356 21252 41412
rect 21308 40514 21364 40516
rect 21308 40462 21310 40514
rect 21310 40462 21362 40514
rect 21362 40462 21364 40514
rect 21308 40460 21364 40462
rect 18844 38108 18900 38164
rect 18508 37436 18564 37492
rect 18620 37548 18676 37604
rect 18508 35698 18564 35700
rect 18508 35646 18510 35698
rect 18510 35646 18562 35698
rect 18562 35646 18564 35698
rect 18508 35644 18564 35646
rect 18844 35644 18900 35700
rect 18620 33180 18676 33236
rect 18844 32674 18900 32676
rect 18844 32622 18846 32674
rect 18846 32622 18898 32674
rect 18898 32622 18900 32674
rect 18844 32620 18900 32622
rect 18508 32562 18564 32564
rect 18508 32510 18510 32562
rect 18510 32510 18562 32562
rect 18562 32510 18564 32562
rect 18508 32508 18564 32510
rect 18620 31890 18676 31892
rect 18620 31838 18622 31890
rect 18622 31838 18674 31890
rect 18674 31838 18676 31890
rect 18620 31836 18676 31838
rect 19404 38332 19460 38388
rect 19628 38220 19684 38276
rect 20188 38050 20244 38052
rect 20188 37998 20190 38050
rect 20190 37998 20242 38050
rect 20242 37998 20244 38050
rect 20188 37996 20244 37998
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20636 37772 20692 37828
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19964 35644 20020 35700
rect 19180 34018 19236 34020
rect 19180 33966 19182 34018
rect 19182 33966 19234 34018
rect 19234 33966 19236 34018
rect 19180 33964 19236 33966
rect 19068 33068 19124 33124
rect 18844 29036 18900 29092
rect 18620 28476 18676 28532
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20300 37266 20356 37268
rect 20300 37214 20302 37266
rect 20302 37214 20354 37266
rect 20354 37214 20356 37266
rect 20300 37212 20356 37214
rect 20412 37154 20468 37156
rect 20412 37102 20414 37154
rect 20414 37102 20466 37154
rect 20466 37102 20468 37154
rect 20412 37100 20468 37102
rect 20300 36428 20356 36484
rect 20636 37042 20692 37044
rect 20636 36990 20638 37042
rect 20638 36990 20690 37042
rect 20690 36990 20692 37042
rect 20636 36988 20692 36990
rect 20748 36258 20804 36260
rect 20748 36206 20750 36258
rect 20750 36206 20802 36258
rect 20802 36206 20804 36258
rect 20748 36204 20804 36206
rect 21084 39788 21140 39844
rect 21196 39564 21252 39620
rect 21308 39506 21364 39508
rect 21308 39454 21310 39506
rect 21310 39454 21362 39506
rect 21362 39454 21364 39506
rect 21308 39452 21364 39454
rect 21308 38834 21364 38836
rect 21308 38782 21310 38834
rect 21310 38782 21362 38834
rect 21362 38782 21364 38834
rect 21308 38780 21364 38782
rect 22652 42028 22708 42084
rect 22316 41916 22372 41972
rect 21868 40402 21924 40404
rect 21868 40350 21870 40402
rect 21870 40350 21922 40402
rect 21922 40350 21924 40402
rect 21868 40348 21924 40350
rect 21532 38332 21588 38388
rect 21420 38220 21476 38276
rect 21308 38108 21364 38164
rect 20972 37884 21028 37940
rect 21644 37772 21700 37828
rect 21756 38780 21812 38836
rect 21868 38220 21924 38276
rect 22092 37938 22148 37940
rect 22092 37886 22094 37938
rect 22094 37886 22146 37938
rect 22146 37886 22148 37938
rect 22092 37884 22148 37886
rect 20972 37100 21028 37156
rect 21196 37212 21252 37268
rect 21308 36258 21364 36260
rect 21308 36206 21310 36258
rect 21310 36206 21362 36258
rect 21362 36206 21364 36258
rect 21308 36204 21364 36206
rect 20748 35756 20804 35812
rect 19404 32786 19460 32788
rect 19404 32734 19406 32786
rect 19406 32734 19458 32786
rect 19458 32734 19460 32786
rect 19404 32732 19460 32734
rect 20076 33122 20132 33124
rect 20076 33070 20078 33122
rect 20078 33070 20130 33122
rect 20130 33070 20132 33122
rect 20076 33068 20132 33070
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 32508 19684 32564
rect 19964 32620 20020 32676
rect 19852 31948 19908 32004
rect 19404 31778 19460 31780
rect 19404 31726 19406 31778
rect 19406 31726 19458 31778
rect 19458 31726 19460 31778
rect 19404 31724 19460 31726
rect 20300 31724 20356 31780
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20300 30828 20356 30884
rect 19628 30210 19684 30212
rect 19628 30158 19630 30210
rect 19630 30158 19682 30210
rect 19682 30158 19684 30210
rect 19628 30156 19684 30158
rect 18956 28588 19012 28644
rect 18620 27580 18676 27636
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19628 28812 19684 28868
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19628 27858 19684 27860
rect 19628 27806 19630 27858
rect 19630 27806 19682 27858
rect 19682 27806 19684 27858
rect 19628 27804 19684 27806
rect 19292 27580 19348 27636
rect 19180 25564 19236 25620
rect 18284 25004 18340 25060
rect 18172 24892 18228 24948
rect 17612 24332 17668 24388
rect 16380 23884 16436 23940
rect 19180 24946 19236 24948
rect 19180 24894 19182 24946
rect 19182 24894 19234 24946
rect 19234 24894 19236 24946
rect 19180 24892 19236 24894
rect 22540 41244 22596 41300
rect 22428 38556 22484 38612
rect 23660 43932 23716 43988
rect 23660 42082 23716 42084
rect 23660 42030 23662 42082
rect 23662 42030 23714 42082
rect 23714 42030 23716 42082
rect 23660 42028 23716 42030
rect 23660 41804 23716 41860
rect 23324 41580 23380 41636
rect 23436 41468 23492 41524
rect 23772 41356 23828 41412
rect 22204 36876 22260 36932
rect 22988 40402 23044 40404
rect 22988 40350 22990 40402
rect 22990 40350 23042 40402
rect 23042 40350 23044 40402
rect 22988 40348 23044 40350
rect 22652 39730 22708 39732
rect 22652 39678 22654 39730
rect 22654 39678 22706 39730
rect 22706 39678 22708 39730
rect 22652 39676 22708 39678
rect 23436 41186 23492 41188
rect 23436 41134 23438 41186
rect 23438 41134 23490 41186
rect 23490 41134 23492 41186
rect 23436 41132 23492 41134
rect 23436 40684 23492 40740
rect 23436 39676 23492 39732
rect 23772 40402 23828 40404
rect 23772 40350 23774 40402
rect 23774 40350 23826 40402
rect 23826 40350 23828 40402
rect 23772 40348 23828 40350
rect 25452 47068 25508 47124
rect 24556 46898 24612 46900
rect 24556 46846 24558 46898
rect 24558 46846 24610 46898
rect 24610 46846 24612 46898
rect 24556 46844 24612 46846
rect 25228 46620 25284 46676
rect 24780 45052 24836 45108
rect 24444 44268 24500 44324
rect 24108 44210 24164 44212
rect 24108 44158 24110 44210
rect 24110 44158 24162 44210
rect 24162 44158 24164 44210
rect 24108 44156 24164 44158
rect 25340 45052 25396 45108
rect 24668 44156 24724 44212
rect 25564 44210 25620 44212
rect 25564 44158 25566 44210
rect 25566 44158 25618 44210
rect 25618 44158 25620 44210
rect 25564 44156 25620 44158
rect 23996 41916 24052 41972
rect 25116 41804 25172 41860
rect 26460 57372 26516 57428
rect 26684 56866 26740 56868
rect 26684 56814 26686 56866
rect 26686 56814 26738 56866
rect 26738 56814 26740 56866
rect 26684 56812 26740 56814
rect 28364 60226 28420 60228
rect 28364 60174 28366 60226
rect 28366 60174 28418 60226
rect 28418 60174 28420 60226
rect 28364 60172 28420 60174
rect 27692 57762 27748 57764
rect 27692 57710 27694 57762
rect 27694 57710 27746 57762
rect 27746 57710 27748 57762
rect 27692 57708 27748 57710
rect 28252 57650 28308 57652
rect 28252 57598 28254 57650
rect 28254 57598 28306 57650
rect 28306 57598 28308 57650
rect 28252 57596 28308 57598
rect 27692 56812 27748 56868
rect 25788 48748 25844 48804
rect 27020 55020 27076 55076
rect 26684 54626 26740 54628
rect 26684 54574 26686 54626
rect 26686 54574 26738 54626
rect 26738 54574 26740 54626
rect 26684 54572 26740 54574
rect 26236 50482 26292 50484
rect 26236 50430 26238 50482
rect 26238 50430 26290 50482
rect 26290 50430 26292 50482
rect 26236 50428 26292 50430
rect 28924 62860 28980 62916
rect 29484 64706 29540 64708
rect 29484 64654 29486 64706
rect 29486 64654 29538 64706
rect 29538 64654 29540 64706
rect 29484 64652 29540 64654
rect 30380 64706 30436 64708
rect 30380 64654 30382 64706
rect 30382 64654 30434 64706
rect 30434 64654 30436 64706
rect 30380 64652 30436 64654
rect 30940 64594 30996 64596
rect 30940 64542 30942 64594
rect 30942 64542 30994 64594
rect 30994 64542 30996 64594
rect 30940 64540 30996 64542
rect 30156 63138 30212 63140
rect 30156 63086 30158 63138
rect 30158 63086 30210 63138
rect 30210 63086 30212 63138
rect 30156 63084 30212 63086
rect 29484 62860 29540 62916
rect 29484 62300 29540 62356
rect 30940 63084 30996 63140
rect 31724 63810 31780 63812
rect 31724 63758 31726 63810
rect 31726 63758 31778 63810
rect 31778 63758 31780 63810
rect 31724 63756 31780 63758
rect 31948 63532 32004 63588
rect 31276 63362 31332 63364
rect 31276 63310 31278 63362
rect 31278 63310 31330 63362
rect 31330 63310 31332 63362
rect 31276 63308 31332 63310
rect 31948 63308 32004 63364
rect 31276 63084 31332 63140
rect 32956 64594 33012 64596
rect 32956 64542 32958 64594
rect 32958 64542 33010 64594
rect 33010 64542 33012 64594
rect 32956 64540 33012 64542
rect 32284 63868 32340 63924
rect 32508 63922 32564 63924
rect 32508 63870 32510 63922
rect 32510 63870 32562 63922
rect 32562 63870 32564 63922
rect 32508 63868 32564 63870
rect 32844 63532 32900 63588
rect 33292 64482 33348 64484
rect 33292 64430 33294 64482
rect 33294 64430 33346 64482
rect 33346 64430 33348 64482
rect 33292 64428 33348 64430
rect 33180 63868 33236 63924
rect 33068 63308 33124 63364
rect 29596 61068 29652 61124
rect 28924 60786 28980 60788
rect 28924 60734 28926 60786
rect 28926 60734 28978 60786
rect 28978 60734 28980 60786
rect 28924 60732 28980 60734
rect 28700 60674 28756 60676
rect 28700 60622 28702 60674
rect 28702 60622 28754 60674
rect 28754 60622 28756 60674
rect 28700 60620 28756 60622
rect 29260 60172 29316 60228
rect 29372 60002 29428 60004
rect 29372 59950 29374 60002
rect 29374 59950 29426 60002
rect 29426 59950 29428 60002
rect 29372 59948 29428 59950
rect 30044 60674 30100 60676
rect 30044 60622 30046 60674
rect 30046 60622 30098 60674
rect 30098 60622 30100 60674
rect 30044 60620 30100 60622
rect 30492 60674 30548 60676
rect 30492 60622 30494 60674
rect 30494 60622 30546 60674
rect 30546 60622 30548 60674
rect 30492 60620 30548 60622
rect 30828 60620 30884 60676
rect 31052 61292 31108 61348
rect 29932 60562 29988 60564
rect 29932 60510 29934 60562
rect 29934 60510 29986 60562
rect 29986 60510 29988 60562
rect 29932 60508 29988 60510
rect 30380 59836 30436 59892
rect 30380 59500 30436 59556
rect 32956 62188 33012 62244
rect 34860 65436 34916 65492
rect 35532 65490 35588 65492
rect 35532 65438 35534 65490
rect 35534 65438 35586 65490
rect 35586 65438 35588 65490
rect 35532 65436 35588 65438
rect 34972 65378 35028 65380
rect 34972 65326 34974 65378
rect 34974 65326 35026 65378
rect 35026 65326 35028 65378
rect 34972 65324 35028 65326
rect 35644 65324 35700 65380
rect 34636 64428 34692 64484
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 37436 65212 37492 65268
rect 38556 65324 38612 65380
rect 36652 64652 36708 64708
rect 37100 64706 37156 64708
rect 37100 64654 37102 64706
rect 37102 64654 37154 64706
rect 37154 64654 37156 64706
rect 37100 64652 37156 64654
rect 38556 64706 38612 64708
rect 38556 64654 38558 64706
rect 38558 64654 38610 64706
rect 38610 64654 38612 64706
rect 38556 64652 38612 64654
rect 39228 64092 39284 64148
rect 45052 66444 45108 66500
rect 43036 66162 43092 66164
rect 43036 66110 43038 66162
rect 43038 66110 43090 66162
rect 43090 66110 43092 66162
rect 43036 66108 43092 66110
rect 46172 66108 46228 66164
rect 41020 65436 41076 65492
rect 42700 65436 42756 65492
rect 41132 65378 41188 65380
rect 41132 65326 41134 65378
rect 41134 65326 41186 65378
rect 41186 65326 41188 65378
rect 41132 65324 41188 65326
rect 40124 65212 40180 65268
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 37884 62748 37940 62804
rect 37436 62412 37492 62468
rect 32396 61346 32452 61348
rect 32396 61294 32398 61346
rect 32398 61294 32450 61346
rect 32450 61294 32452 61346
rect 32396 61292 32452 61294
rect 31276 60620 31332 60676
rect 31052 59724 31108 59780
rect 31164 60002 31220 60004
rect 31164 59950 31166 60002
rect 31166 59950 31218 60002
rect 31218 59950 31220 60002
rect 31164 59948 31220 59950
rect 29820 58322 29876 58324
rect 29820 58270 29822 58322
rect 29822 58270 29874 58322
rect 29874 58270 29876 58322
rect 29820 58268 29876 58270
rect 30492 58322 30548 58324
rect 30492 58270 30494 58322
rect 30494 58270 30546 58322
rect 30546 58270 30548 58322
rect 30492 58268 30548 58270
rect 30044 57260 30100 57316
rect 30156 57596 30212 57652
rect 27580 54514 27636 54516
rect 27580 54462 27582 54514
rect 27582 54462 27634 54514
rect 27634 54462 27636 54514
rect 27580 54460 27636 54462
rect 27916 55074 27972 55076
rect 27916 55022 27918 55074
rect 27918 55022 27970 55074
rect 27970 55022 27972 55074
rect 27916 55020 27972 55022
rect 28140 53842 28196 53844
rect 28140 53790 28142 53842
rect 28142 53790 28194 53842
rect 28194 53790 28196 53842
rect 28140 53788 28196 53790
rect 28476 54402 28532 54404
rect 28476 54350 28478 54402
rect 28478 54350 28530 54402
rect 28530 54350 28532 54402
rect 28476 54348 28532 54350
rect 29148 54402 29204 54404
rect 29148 54350 29150 54402
rect 29150 54350 29202 54402
rect 29202 54350 29204 54402
rect 29148 54348 29204 54350
rect 29372 55020 29428 55076
rect 30604 57260 30660 57316
rect 30940 57650 30996 57652
rect 30940 57598 30942 57650
rect 30942 57598 30994 57650
rect 30994 57598 30996 57650
rect 30940 57596 30996 57598
rect 30828 55020 30884 55076
rect 30380 54684 30436 54740
rect 29372 53954 29428 53956
rect 29372 53902 29374 53954
rect 29374 53902 29426 53954
rect 29426 53902 29428 53954
rect 29372 53900 29428 53902
rect 28924 53788 28980 53844
rect 28028 51212 28084 51268
rect 27356 49420 27412 49476
rect 26124 48188 26180 48244
rect 27468 48242 27524 48244
rect 27468 48190 27470 48242
rect 27470 48190 27522 48242
rect 27522 48190 27524 48242
rect 27468 48188 27524 48190
rect 26012 46508 26068 46564
rect 26236 46060 26292 46116
rect 26236 45106 26292 45108
rect 26236 45054 26238 45106
rect 26238 45054 26290 45106
rect 26290 45054 26292 45106
rect 26236 45052 26292 45054
rect 25900 43708 25956 43764
rect 26012 42754 26068 42756
rect 26012 42702 26014 42754
rect 26014 42702 26066 42754
rect 26066 42702 26068 42754
rect 26012 42700 26068 42702
rect 25116 41356 25172 41412
rect 24780 41244 24836 41300
rect 24332 41132 24388 41188
rect 24892 41132 24948 41188
rect 25564 41244 25620 41300
rect 24444 40796 24500 40852
rect 24108 40514 24164 40516
rect 24108 40462 24110 40514
rect 24110 40462 24162 40514
rect 24162 40462 24164 40514
rect 24108 40460 24164 40462
rect 23996 40348 24052 40404
rect 23660 38892 23716 38948
rect 24220 39340 24276 39396
rect 22652 38220 22708 38276
rect 23212 38556 23268 38612
rect 22876 37154 22932 37156
rect 22876 37102 22878 37154
rect 22878 37102 22930 37154
rect 22930 37102 22932 37154
rect 22876 37100 22932 37102
rect 22876 36876 22932 36932
rect 21644 35644 21700 35700
rect 22540 35644 22596 35700
rect 21644 35474 21700 35476
rect 21644 35422 21646 35474
rect 21646 35422 21698 35474
rect 21698 35422 21700 35474
rect 21644 35420 21700 35422
rect 21420 34076 21476 34132
rect 21308 34018 21364 34020
rect 21308 33966 21310 34018
rect 21310 33966 21362 34018
rect 21362 33966 21364 34018
rect 21308 33964 21364 33966
rect 21420 33068 21476 33124
rect 20636 32172 20692 32228
rect 20524 30156 20580 30212
rect 21084 31948 21140 32004
rect 20972 30044 21028 30100
rect 21196 30882 21252 30884
rect 21196 30830 21198 30882
rect 21198 30830 21250 30882
rect 21250 30830 21252 30882
rect 21196 30828 21252 30830
rect 22540 33404 22596 33460
rect 22092 33234 22148 33236
rect 22092 33182 22094 33234
rect 22094 33182 22146 33234
rect 22146 33182 22148 33234
rect 22092 33180 22148 33182
rect 21980 31164 22036 31220
rect 22540 31218 22596 31220
rect 22540 31166 22542 31218
rect 22542 31166 22594 31218
rect 22594 31166 22596 31218
rect 22540 31164 22596 31166
rect 22092 31106 22148 31108
rect 22092 31054 22094 31106
rect 22094 31054 22146 31106
rect 22146 31054 22148 31106
rect 22092 31052 22148 31054
rect 22092 30716 22148 30772
rect 22204 30380 22260 30436
rect 21532 30044 21588 30100
rect 21868 30044 21924 30100
rect 21532 29538 21588 29540
rect 21532 29486 21534 29538
rect 21534 29486 21586 29538
rect 21586 29486 21588 29538
rect 21532 29484 21588 29486
rect 21084 29148 21140 29204
rect 21644 28924 21700 28980
rect 22316 30044 22372 30100
rect 22204 29932 22260 29988
rect 22764 36482 22820 36484
rect 22764 36430 22766 36482
rect 22766 36430 22818 36482
rect 22818 36430 22820 36482
rect 22764 36428 22820 36430
rect 23100 37884 23156 37940
rect 22988 35644 23044 35700
rect 22764 33516 22820 33572
rect 22876 30994 22932 30996
rect 22876 30942 22878 30994
rect 22878 30942 22930 30994
rect 22930 30942 22932 30994
rect 22876 30940 22932 30942
rect 23884 38722 23940 38724
rect 23884 38670 23886 38722
rect 23886 38670 23938 38722
rect 23938 38670 23940 38722
rect 23884 38668 23940 38670
rect 23324 36428 23380 36484
rect 23324 35308 23380 35364
rect 23996 38556 24052 38612
rect 24220 38610 24276 38612
rect 24220 38558 24222 38610
rect 24222 38558 24274 38610
rect 24274 38558 24276 38610
rect 24220 38556 24276 38558
rect 24108 37996 24164 38052
rect 23996 37938 24052 37940
rect 23996 37886 23998 37938
rect 23998 37886 24050 37938
rect 24050 37886 24052 37938
rect 23996 37884 24052 37886
rect 24220 37884 24276 37940
rect 26012 41132 26068 41188
rect 25004 39676 25060 39732
rect 26124 39730 26180 39732
rect 26124 39678 26126 39730
rect 26126 39678 26178 39730
rect 26178 39678 26180 39730
rect 26124 39676 26180 39678
rect 25564 39618 25620 39620
rect 25564 39566 25566 39618
rect 25566 39566 25618 39618
rect 25618 39566 25620 39618
rect 25564 39564 25620 39566
rect 24780 39116 24836 39172
rect 24444 38892 24500 38948
rect 23660 36876 23716 36932
rect 23884 37100 23940 37156
rect 24332 36316 24388 36372
rect 24220 35922 24276 35924
rect 24220 35870 24222 35922
rect 24222 35870 24274 35922
rect 24274 35870 24276 35922
rect 24220 35868 24276 35870
rect 23548 33516 23604 33572
rect 24556 38780 24612 38836
rect 26236 38892 26292 38948
rect 25676 38834 25732 38836
rect 25676 38782 25678 38834
rect 25678 38782 25730 38834
rect 25730 38782 25732 38834
rect 25676 38780 25732 38782
rect 26012 38780 26068 38836
rect 24556 37884 24612 37940
rect 24892 38108 24948 38164
rect 24556 37266 24612 37268
rect 24556 37214 24558 37266
rect 24558 37214 24610 37266
rect 24610 37214 24612 37266
rect 24556 37212 24612 37214
rect 25340 37996 25396 38052
rect 25340 37490 25396 37492
rect 25340 37438 25342 37490
rect 25342 37438 25394 37490
rect 25394 37438 25396 37490
rect 25340 37436 25396 37438
rect 24892 37212 24948 37268
rect 25228 37154 25284 37156
rect 25228 37102 25230 37154
rect 25230 37102 25282 37154
rect 25282 37102 25284 37154
rect 25228 37100 25284 37102
rect 23884 33068 23940 33124
rect 25340 35868 25396 35924
rect 25452 35532 25508 35588
rect 26124 38556 26180 38612
rect 26012 37826 26068 37828
rect 26012 37774 26014 37826
rect 26014 37774 26066 37826
rect 26066 37774 26068 37826
rect 26012 37772 26068 37774
rect 26124 37378 26180 37380
rect 26124 37326 26126 37378
rect 26126 37326 26178 37378
rect 26178 37326 26180 37378
rect 26124 37324 26180 37326
rect 26012 35868 26068 35924
rect 25676 35308 25732 35364
rect 25116 33404 25172 33460
rect 24668 33122 24724 33124
rect 24668 33070 24670 33122
rect 24670 33070 24722 33122
rect 24722 33070 24724 33122
rect 24668 33068 24724 33070
rect 25788 33234 25844 33236
rect 25788 33182 25790 33234
rect 25790 33182 25842 33234
rect 25842 33182 25844 33234
rect 25788 33180 25844 33182
rect 24108 31836 24164 31892
rect 23100 30380 23156 30436
rect 22876 29986 22932 29988
rect 22876 29934 22878 29986
rect 22878 29934 22930 29986
rect 22930 29934 22932 29986
rect 22876 29932 22932 29934
rect 22092 29538 22148 29540
rect 22092 29486 22094 29538
rect 22094 29486 22146 29538
rect 22146 29486 22148 29538
rect 22092 29484 22148 29486
rect 22428 29538 22484 29540
rect 22428 29486 22430 29538
rect 22430 29486 22482 29538
rect 22482 29486 22484 29538
rect 22428 29484 22484 29486
rect 22876 29148 22932 29204
rect 22876 27858 22932 27860
rect 22876 27806 22878 27858
rect 22878 27806 22930 27858
rect 22930 27806 22932 27858
rect 22876 27804 22932 27806
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19964 25618 20020 25620
rect 19964 25566 19966 25618
rect 19966 25566 20018 25618
rect 20018 25566 20020 25618
rect 19964 25564 20020 25566
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 18620 24332 18676 24388
rect 16604 23714 16660 23716
rect 16604 23662 16606 23714
rect 16606 23662 16658 23714
rect 16658 23662 16660 23714
rect 16604 23660 16660 23662
rect 18284 23660 18340 23716
rect 18844 23996 18900 24052
rect 16716 22988 16772 23044
rect 17500 23042 17556 23044
rect 17500 22990 17502 23042
rect 17502 22990 17554 23042
rect 17554 22990 17556 23042
rect 17500 22988 17556 22990
rect 14812 20188 14868 20244
rect 15932 20690 15988 20692
rect 15932 20638 15934 20690
rect 15934 20638 15986 20690
rect 15986 20638 15988 20690
rect 15932 20636 15988 20638
rect 15260 20188 15316 20244
rect 18620 21810 18676 21812
rect 18620 21758 18622 21810
rect 18622 21758 18674 21810
rect 18674 21758 18676 21810
rect 18620 21756 18676 21758
rect 18172 20076 18228 20132
rect 19404 24050 19460 24052
rect 19404 23998 19406 24050
rect 19406 23998 19458 24050
rect 19458 23998 19460 24050
rect 19404 23996 19460 23998
rect 18956 23938 19012 23940
rect 18956 23886 18958 23938
rect 18958 23886 19010 23938
rect 19010 23886 19012 23938
rect 18956 23884 19012 23886
rect 19852 23660 19908 23716
rect 22876 26908 22932 26964
rect 21420 25116 21476 25172
rect 20412 23996 20468 24052
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18956 23324 19012 23380
rect 19628 23378 19684 23380
rect 19628 23326 19630 23378
rect 19630 23326 19682 23378
rect 19682 23326 19684 23378
rect 19628 23324 19684 23326
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19292 21810 19348 21812
rect 19292 21758 19294 21810
rect 19294 21758 19346 21810
rect 19346 21758 19348 21810
rect 19292 21756 19348 21758
rect 19964 21810 20020 21812
rect 19964 21758 19966 21810
rect 19966 21758 20018 21810
rect 20018 21758 20020 21810
rect 19964 21756 20020 21758
rect 18956 21698 19012 21700
rect 18956 21646 18958 21698
rect 18958 21646 19010 21698
rect 19010 21646 19012 21698
rect 18956 21644 19012 21646
rect 18060 20018 18116 20020
rect 18060 19966 18062 20018
rect 18062 19966 18114 20018
rect 18114 19966 18116 20018
rect 18060 19964 18116 19966
rect 18732 20860 18788 20916
rect 18508 20690 18564 20692
rect 18508 20638 18510 20690
rect 18510 20638 18562 20690
rect 18562 20638 18564 20690
rect 18508 20636 18564 20638
rect 18396 20524 18452 20580
rect 18620 20076 18676 20132
rect 17164 18956 17220 19012
rect 17836 18956 17892 19012
rect 15036 18396 15092 18452
rect 17388 18284 17444 18340
rect 14700 17388 14756 17444
rect 17500 17442 17556 17444
rect 17500 17390 17502 17442
rect 17502 17390 17554 17442
rect 17554 17390 17556 17442
rect 17500 17388 17556 17390
rect 17388 17276 17444 17332
rect 18508 19010 18564 19012
rect 18508 18958 18510 19010
rect 18510 18958 18562 19010
rect 18562 18958 18564 19010
rect 18508 18956 18564 18958
rect 18060 18450 18116 18452
rect 18060 18398 18062 18450
rect 18062 18398 18114 18450
rect 18114 18398 18116 18450
rect 18060 18396 18116 18398
rect 18284 18450 18340 18452
rect 18284 18398 18286 18450
rect 18286 18398 18338 18450
rect 18338 18398 18340 18450
rect 18284 18396 18340 18398
rect 17948 18284 18004 18340
rect 17724 17164 17780 17220
rect 16828 17052 16884 17108
rect 16716 16940 16772 16996
rect 12908 16268 12964 16324
rect 14028 16156 14084 16212
rect 15932 16716 15988 16772
rect 15932 16156 15988 16212
rect 18060 17052 18116 17108
rect 17612 16882 17668 16884
rect 17612 16830 17614 16882
rect 17614 16830 17666 16882
rect 17666 16830 17668 16882
rect 17612 16828 17668 16830
rect 14700 13916 14756 13972
rect 16828 13634 16884 13636
rect 16828 13582 16830 13634
rect 16830 13582 16882 13634
rect 16882 13582 16884 13634
rect 16828 13580 16884 13582
rect 17500 13468 17556 13524
rect 17836 13186 17892 13188
rect 17836 13134 17838 13186
rect 17838 13134 17890 13186
rect 17890 13134 17892 13186
rect 17836 13132 17892 13134
rect 17948 12962 18004 12964
rect 17948 12910 17950 12962
rect 17950 12910 18002 12962
rect 18002 12910 18004 12962
rect 17948 12908 18004 12910
rect 17836 12738 17892 12740
rect 17836 12686 17838 12738
rect 17838 12686 17890 12738
rect 17890 12686 17892 12738
rect 17836 12684 17892 12686
rect 5852 11676 5908 11732
rect 14476 11676 14532 11732
rect 17724 11676 17780 11732
rect 17276 11506 17332 11508
rect 17276 11454 17278 11506
rect 17278 11454 17330 11506
rect 17330 11454 17332 11506
rect 17276 11452 17332 11454
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 15820 11116 15876 11172
rect 17276 9772 17332 9828
rect 15820 9548 15876 9604
rect 18284 17442 18340 17444
rect 18284 17390 18286 17442
rect 18286 17390 18338 17442
rect 18338 17390 18340 17442
rect 18284 17388 18340 17390
rect 18396 17276 18452 17332
rect 18284 17164 18340 17220
rect 18508 17052 18564 17108
rect 18732 17106 18788 17108
rect 18732 17054 18734 17106
rect 18734 17054 18786 17106
rect 18786 17054 18788 17106
rect 18732 17052 18788 17054
rect 19068 19292 19124 19348
rect 19068 18450 19124 18452
rect 19068 18398 19070 18450
rect 19070 18398 19122 18450
rect 19122 18398 19124 18450
rect 19068 18396 19124 18398
rect 18956 17666 19012 17668
rect 18956 17614 18958 17666
rect 18958 17614 19010 17666
rect 19010 17614 19012 17666
rect 18956 17612 19012 17614
rect 19404 20914 19460 20916
rect 19404 20862 19406 20914
rect 19406 20862 19458 20914
rect 19458 20862 19460 20914
rect 19404 20860 19460 20862
rect 20076 21644 20132 21700
rect 20748 23714 20804 23716
rect 20748 23662 20750 23714
rect 20750 23662 20802 23714
rect 20802 23662 20804 23714
rect 20748 23660 20804 23662
rect 20748 23212 20804 23268
rect 20300 20860 20356 20916
rect 20524 20802 20580 20804
rect 20524 20750 20526 20802
rect 20526 20750 20578 20802
rect 20578 20750 20580 20802
rect 20524 20748 20580 20750
rect 20748 20690 20804 20692
rect 20748 20638 20750 20690
rect 20750 20638 20802 20690
rect 20802 20638 20804 20690
rect 20748 20636 20804 20638
rect 19628 20524 19684 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19404 20018 19460 20020
rect 19404 19966 19406 20018
rect 19406 19966 19458 20018
rect 19458 19966 19460 20018
rect 19404 19964 19460 19966
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19852 18060 19908 18116
rect 21532 17724 21588 17780
rect 22876 26572 22932 26628
rect 22316 26178 22372 26180
rect 22316 26126 22318 26178
rect 22318 26126 22370 26178
rect 22370 26126 22372 26178
rect 22316 26124 22372 26126
rect 22764 26124 22820 26180
rect 21756 25228 21812 25284
rect 22204 25116 22260 25172
rect 22540 25282 22596 25284
rect 22540 25230 22542 25282
rect 22542 25230 22594 25282
rect 22594 25230 22596 25282
rect 22540 25228 22596 25230
rect 22204 23938 22260 23940
rect 22204 23886 22206 23938
rect 22206 23886 22258 23938
rect 22258 23886 22260 23938
rect 22204 23884 22260 23886
rect 21980 23324 22036 23380
rect 22428 23548 22484 23604
rect 22652 24610 22708 24612
rect 22652 24558 22654 24610
rect 22654 24558 22706 24610
rect 22706 24558 22708 24610
rect 22652 24556 22708 24558
rect 23212 29650 23268 29652
rect 23212 29598 23214 29650
rect 23214 29598 23266 29650
rect 23266 29598 23268 29650
rect 23212 29596 23268 29598
rect 23436 30994 23492 30996
rect 23436 30942 23438 30994
rect 23438 30942 23490 30994
rect 23490 30942 23492 30994
rect 23436 30940 23492 30942
rect 23996 30994 24052 30996
rect 23996 30942 23998 30994
rect 23998 30942 24050 30994
rect 24050 30942 24052 30994
rect 23996 30940 24052 30942
rect 23996 30156 24052 30212
rect 24220 30098 24276 30100
rect 24220 30046 24222 30098
rect 24222 30046 24274 30098
rect 24274 30046 24276 30098
rect 24220 30044 24276 30046
rect 24444 29986 24500 29988
rect 24444 29934 24446 29986
rect 24446 29934 24498 29986
rect 24498 29934 24500 29986
rect 24444 29932 24500 29934
rect 23660 29538 23716 29540
rect 23660 29486 23662 29538
rect 23662 29486 23714 29538
rect 23714 29486 23716 29538
rect 23660 29484 23716 29486
rect 24780 29372 24836 29428
rect 23996 26908 24052 26964
rect 23212 25788 23268 25844
rect 23324 26124 23380 26180
rect 23772 26124 23828 26180
rect 22988 24332 23044 24388
rect 23100 23548 23156 23604
rect 22876 23324 22932 23380
rect 21756 21586 21812 21588
rect 21756 21534 21758 21586
rect 21758 21534 21810 21586
rect 21810 21534 21812 21586
rect 21756 21532 21812 21534
rect 21868 20690 21924 20692
rect 21868 20638 21870 20690
rect 21870 20638 21922 20690
rect 21922 20638 21924 20690
rect 21868 20636 21924 20638
rect 21756 20578 21812 20580
rect 21756 20526 21758 20578
rect 21758 20526 21810 20578
rect 21810 20526 21812 20578
rect 21756 20524 21812 20526
rect 22652 22764 22708 22820
rect 22652 20748 22708 20804
rect 22988 23154 23044 23156
rect 22988 23102 22990 23154
rect 22990 23102 23042 23154
rect 23042 23102 23044 23154
rect 22988 23100 23044 23102
rect 21980 19852 22036 19908
rect 22876 19852 22932 19908
rect 19180 17388 19236 17444
rect 18508 15932 18564 15988
rect 18508 14530 18564 14532
rect 18508 14478 18510 14530
rect 18510 14478 18562 14530
rect 18562 14478 18564 14530
rect 18508 14476 18564 14478
rect 18284 13356 18340 13412
rect 18284 13132 18340 13188
rect 18284 12012 18340 12068
rect 21196 17388 21252 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16882 19684 16884
rect 19628 16830 19630 16882
rect 19630 16830 19682 16882
rect 19682 16830 19684 16882
rect 19628 16828 19684 16830
rect 22316 17778 22372 17780
rect 22316 17726 22318 17778
rect 22318 17726 22370 17778
rect 22370 17726 22372 17778
rect 22316 17724 22372 17726
rect 22428 17612 22484 17668
rect 21756 16156 21812 16212
rect 19292 15986 19348 15988
rect 19292 15934 19294 15986
rect 19294 15934 19346 15986
rect 19346 15934 19348 15986
rect 19292 15932 19348 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 22428 16210 22484 16212
rect 22428 16158 22430 16210
rect 22430 16158 22482 16210
rect 22482 16158 22484 16210
rect 22428 16156 22484 16158
rect 22764 16156 22820 16212
rect 23212 19180 23268 19236
rect 23100 18396 23156 18452
rect 23436 24556 23492 24612
rect 24556 26850 24612 26852
rect 24556 26798 24558 26850
rect 24558 26798 24610 26850
rect 24610 26798 24612 26850
rect 24556 26796 24612 26798
rect 24108 26178 24164 26180
rect 24108 26126 24110 26178
rect 24110 26126 24162 26178
rect 24162 26126 24164 26178
rect 24108 26124 24164 26126
rect 24108 25730 24164 25732
rect 24108 25678 24110 25730
rect 24110 25678 24162 25730
rect 24162 25678 24164 25730
rect 24108 25676 24164 25678
rect 24220 25506 24276 25508
rect 24220 25454 24222 25506
rect 24222 25454 24274 25506
rect 24274 25454 24276 25506
rect 24220 25452 24276 25454
rect 24108 25394 24164 25396
rect 24108 25342 24110 25394
rect 24110 25342 24162 25394
rect 24162 25342 24164 25394
rect 24108 25340 24164 25342
rect 24556 25788 24612 25844
rect 25900 30156 25956 30212
rect 25452 29932 25508 29988
rect 25228 29372 25284 29428
rect 25564 29650 25620 29652
rect 25564 29598 25566 29650
rect 25566 29598 25618 29650
rect 25618 29598 25620 29650
rect 25564 29596 25620 29598
rect 25564 29148 25620 29204
rect 25452 28588 25508 28644
rect 25788 27692 25844 27748
rect 26460 46956 26516 47012
rect 27244 47180 27300 47236
rect 26460 46060 26516 46116
rect 27468 46956 27524 47012
rect 27132 42754 27188 42756
rect 27132 42702 27134 42754
rect 27134 42702 27186 42754
rect 27186 42702 27188 42754
rect 27132 42700 27188 42702
rect 27244 42082 27300 42084
rect 27244 42030 27246 42082
rect 27246 42030 27298 42082
rect 27298 42030 27300 42082
rect 27244 42028 27300 42030
rect 26908 41132 26964 41188
rect 26460 41074 26516 41076
rect 26460 41022 26462 41074
rect 26462 41022 26514 41074
rect 26514 41022 26516 41074
rect 26460 41020 26516 41022
rect 26572 40796 26628 40852
rect 26460 39618 26516 39620
rect 26460 39566 26462 39618
rect 26462 39566 26514 39618
rect 26514 39566 26516 39618
rect 26460 39564 26516 39566
rect 27692 48188 27748 48244
rect 27916 47964 27972 48020
rect 29036 53452 29092 53508
rect 28252 50876 28308 50932
rect 28588 51154 28644 51156
rect 28588 51102 28590 51154
rect 28590 51102 28642 51154
rect 28642 51102 28644 51154
rect 28588 51100 28644 51102
rect 29260 51100 29316 51156
rect 29372 50764 29428 50820
rect 28812 49980 28868 50036
rect 28700 49810 28756 49812
rect 28700 49758 28702 49810
rect 28702 49758 28754 49810
rect 28754 49758 28756 49810
rect 28700 49756 28756 49758
rect 28364 48354 28420 48356
rect 28364 48302 28366 48354
rect 28366 48302 28418 48354
rect 28418 48302 28420 48354
rect 28364 48300 28420 48302
rect 28252 48242 28308 48244
rect 28252 48190 28254 48242
rect 28254 48190 28306 48242
rect 28306 48190 28308 48242
rect 28252 48188 28308 48190
rect 28364 48018 28420 48020
rect 28364 47966 28366 48018
rect 28366 47966 28418 48018
rect 28418 47966 28420 48018
rect 28364 47964 28420 47966
rect 27692 47180 27748 47236
rect 27916 45052 27972 45108
rect 27804 42812 27860 42868
rect 27916 42140 27972 42196
rect 28028 41916 28084 41972
rect 27580 41244 27636 41300
rect 27356 40908 27412 40964
rect 27804 41356 27860 41412
rect 27468 40572 27524 40628
rect 27580 40348 27636 40404
rect 26908 39116 26964 39172
rect 26684 39004 26740 39060
rect 26572 38892 26628 38948
rect 27804 40684 27860 40740
rect 27468 39394 27524 39396
rect 27468 39342 27470 39394
rect 27470 39342 27522 39394
rect 27522 39342 27524 39394
rect 27468 39340 27524 39342
rect 26908 38722 26964 38724
rect 26908 38670 26910 38722
rect 26910 38670 26962 38722
rect 26962 38670 26964 38722
rect 26908 38668 26964 38670
rect 27020 38162 27076 38164
rect 27020 38110 27022 38162
rect 27022 38110 27074 38162
rect 27074 38110 27076 38162
rect 27020 38108 27076 38110
rect 26572 37996 26628 38052
rect 26796 37212 26852 37268
rect 27132 37324 27188 37380
rect 27356 38556 27412 38612
rect 28140 41356 28196 41412
rect 28140 40908 28196 40964
rect 28028 40684 28084 40740
rect 27916 39340 27972 39396
rect 27692 39058 27748 39060
rect 27692 39006 27694 39058
rect 27694 39006 27746 39058
rect 27746 39006 27748 39058
rect 27692 39004 27748 39006
rect 28028 38834 28084 38836
rect 28028 38782 28030 38834
rect 28030 38782 28082 38834
rect 28082 38782 28084 38834
rect 28028 38780 28084 38782
rect 27468 38050 27524 38052
rect 27468 37998 27470 38050
rect 27470 37998 27522 38050
rect 27522 37998 27524 38050
rect 27468 37996 27524 37998
rect 27580 37884 27636 37940
rect 28140 37938 28196 37940
rect 28140 37886 28142 37938
rect 28142 37886 28194 37938
rect 28194 37886 28196 37938
rect 28140 37884 28196 37886
rect 27580 37436 27636 37492
rect 27020 36428 27076 36484
rect 26908 36316 26964 36372
rect 28476 47570 28532 47572
rect 28476 47518 28478 47570
rect 28478 47518 28530 47570
rect 28530 47518 28532 47570
rect 28476 47516 28532 47518
rect 28700 46786 28756 46788
rect 28700 46734 28702 46786
rect 28702 46734 28754 46786
rect 28754 46734 28756 46786
rect 28700 46732 28756 46734
rect 30940 54572 30996 54628
rect 30380 54012 30436 54068
rect 30044 53506 30100 53508
rect 30044 53454 30046 53506
rect 30046 53454 30098 53506
rect 30098 53454 30100 53506
rect 30044 53452 30100 53454
rect 30604 53452 30660 53508
rect 30716 53676 30772 53732
rect 30716 52780 30772 52836
rect 30940 52220 30996 52276
rect 29708 50876 29764 50932
rect 29820 50652 29876 50708
rect 29596 50540 29652 50596
rect 30716 50652 30772 50708
rect 30156 50594 30212 50596
rect 30156 50542 30158 50594
rect 30158 50542 30210 50594
rect 30210 50542 30212 50594
rect 30156 50540 30212 50542
rect 30604 50482 30660 50484
rect 30604 50430 30606 50482
rect 30606 50430 30658 50482
rect 30658 50430 30660 50482
rect 30604 50428 30660 50430
rect 30940 50764 30996 50820
rect 30492 50034 30548 50036
rect 30492 49982 30494 50034
rect 30494 49982 30546 50034
rect 30546 49982 30548 50034
rect 30492 49980 30548 49982
rect 29820 49810 29876 49812
rect 29820 49758 29822 49810
rect 29822 49758 29874 49810
rect 29874 49758 29876 49810
rect 29820 49756 29876 49758
rect 30492 49084 30548 49140
rect 29372 48300 29428 48356
rect 29820 46786 29876 46788
rect 29820 46734 29822 46786
rect 29822 46734 29874 46786
rect 29874 46734 29876 46786
rect 29820 46732 29876 46734
rect 29820 45948 29876 46004
rect 30156 46172 30212 46228
rect 28476 45106 28532 45108
rect 28476 45054 28478 45106
rect 28478 45054 28530 45106
rect 28530 45054 28532 45106
rect 28476 45052 28532 45054
rect 29148 45052 29204 45108
rect 28364 43484 28420 43540
rect 30156 44940 30212 44996
rect 29148 42754 29204 42756
rect 29148 42702 29150 42754
rect 29150 42702 29202 42754
rect 29202 42702 29204 42754
rect 29148 42700 29204 42702
rect 28588 42476 28644 42532
rect 29820 43650 29876 43652
rect 29820 43598 29822 43650
rect 29822 43598 29874 43650
rect 29874 43598 29876 43650
rect 29820 43596 29876 43598
rect 29932 43538 29988 43540
rect 29932 43486 29934 43538
rect 29934 43486 29986 43538
rect 29986 43486 29988 43538
rect 29932 43484 29988 43486
rect 30156 43484 30212 43540
rect 29708 42812 29764 42868
rect 28364 42140 28420 42196
rect 28588 42028 28644 42084
rect 28588 41692 28644 41748
rect 29484 41970 29540 41972
rect 29484 41918 29486 41970
rect 29486 41918 29538 41970
rect 29538 41918 29540 41970
rect 29484 41916 29540 41918
rect 28924 40572 28980 40628
rect 28588 39900 28644 39956
rect 29372 40348 29428 40404
rect 29260 38556 29316 38612
rect 28588 38050 28644 38052
rect 28588 37998 28590 38050
rect 28590 37998 28642 38050
rect 28642 37998 28644 38050
rect 28588 37996 28644 37998
rect 28364 37826 28420 37828
rect 28364 37774 28366 37826
rect 28366 37774 28418 37826
rect 28418 37774 28420 37826
rect 28364 37772 28420 37774
rect 29148 37996 29204 38052
rect 29260 37938 29316 37940
rect 29260 37886 29262 37938
rect 29262 37886 29314 37938
rect 29314 37886 29316 37938
rect 29260 37884 29316 37886
rect 29260 37212 29316 37268
rect 27356 35532 27412 35588
rect 28364 35026 28420 35028
rect 28364 34974 28366 35026
rect 28366 34974 28418 35026
rect 28418 34974 28420 35026
rect 28364 34972 28420 34974
rect 29148 34972 29204 35028
rect 27916 34300 27972 34356
rect 28364 33628 28420 33684
rect 28140 33346 28196 33348
rect 28140 33294 28142 33346
rect 28142 33294 28194 33346
rect 28194 33294 28196 33346
rect 28140 33292 28196 33294
rect 27468 33180 27524 33236
rect 27804 33068 27860 33124
rect 30044 42028 30100 42084
rect 29708 40572 29764 40628
rect 30604 41356 30660 41412
rect 30268 40460 30324 40516
rect 32060 60508 32116 60564
rect 32396 59890 32452 59892
rect 32396 59838 32398 59890
rect 32398 59838 32450 59890
rect 32450 59838 32452 59890
rect 32396 59836 32452 59838
rect 31388 59052 31444 59108
rect 32284 59106 32340 59108
rect 32284 59054 32286 59106
rect 32286 59054 32338 59106
rect 32338 59054 32340 59106
rect 32284 59052 32340 59054
rect 31612 57260 31668 57316
rect 35868 62300 35924 62356
rect 33180 60284 33236 60340
rect 33292 60508 33348 60564
rect 33404 60284 33460 60340
rect 33628 60002 33684 60004
rect 33628 59950 33630 60002
rect 33630 59950 33682 60002
rect 33682 59950 33684 60002
rect 33628 59948 33684 59950
rect 32396 57650 32452 57652
rect 32396 57598 32398 57650
rect 32398 57598 32450 57650
rect 32450 57598 32452 57650
rect 32396 57596 32452 57598
rect 33180 57596 33236 57652
rect 32284 57036 32340 57092
rect 32396 56924 32452 56980
rect 32508 56194 32564 56196
rect 32508 56142 32510 56194
rect 32510 56142 32562 56194
rect 32562 56142 32564 56194
rect 32508 56140 32564 56142
rect 31612 55132 31668 55188
rect 31500 55074 31556 55076
rect 31500 55022 31502 55074
rect 31502 55022 31554 55074
rect 31554 55022 31556 55074
rect 31500 55020 31556 55022
rect 31388 54684 31444 54740
rect 32284 55186 32340 55188
rect 32284 55134 32286 55186
rect 32286 55134 32338 55186
rect 32338 55134 32340 55186
rect 32284 55132 32340 55134
rect 33068 55132 33124 55188
rect 31948 54626 32004 54628
rect 31948 54574 31950 54626
rect 31950 54574 32002 54626
rect 32002 54574 32004 54626
rect 31948 54572 32004 54574
rect 31276 53900 31332 53956
rect 31276 53170 31332 53172
rect 31276 53118 31278 53170
rect 31278 53118 31330 53170
rect 31330 53118 31332 53170
rect 31276 53116 31332 53118
rect 32396 54236 32452 54292
rect 32172 53116 32228 53172
rect 31948 52834 32004 52836
rect 31948 52782 31950 52834
rect 31950 52782 32002 52834
rect 32002 52782 32004 52834
rect 31948 52780 32004 52782
rect 32508 52444 32564 52500
rect 31836 52108 31892 52164
rect 31948 52220 32004 52276
rect 32396 52274 32452 52276
rect 32396 52222 32398 52274
rect 32398 52222 32450 52274
rect 32450 52222 32452 52274
rect 32396 52220 32452 52222
rect 32284 52162 32340 52164
rect 32284 52110 32286 52162
rect 32286 52110 32338 52162
rect 32338 52110 32340 52162
rect 32284 52108 32340 52110
rect 32284 50876 32340 50932
rect 31164 49698 31220 49700
rect 31164 49646 31166 49698
rect 31166 49646 31218 49698
rect 31218 49646 31220 49698
rect 31164 49644 31220 49646
rect 31164 46172 31220 46228
rect 31052 46002 31108 46004
rect 31052 45950 31054 46002
rect 31054 45950 31106 46002
rect 31106 45950 31108 46002
rect 31052 45948 31108 45950
rect 31164 44268 31220 44324
rect 32508 49868 32564 49924
rect 32732 49756 32788 49812
rect 32060 46844 32116 46900
rect 31388 44156 31444 44212
rect 31276 43596 31332 43652
rect 31276 42866 31332 42868
rect 31276 42814 31278 42866
rect 31278 42814 31330 42866
rect 31330 42814 31332 42866
rect 31276 42812 31332 42814
rect 30940 42476 30996 42532
rect 31164 40460 31220 40516
rect 30044 39004 30100 39060
rect 30828 39340 30884 39396
rect 29932 38722 29988 38724
rect 29932 38670 29934 38722
rect 29934 38670 29986 38722
rect 29986 38670 29988 38722
rect 29932 38668 29988 38670
rect 30604 37938 30660 37940
rect 30604 37886 30606 37938
rect 30606 37886 30658 37938
rect 30658 37886 30660 37938
rect 30604 37884 30660 37886
rect 30268 37212 30324 37268
rect 30156 36092 30212 36148
rect 29596 35196 29652 35252
rect 29708 35644 29764 35700
rect 29932 34860 29988 34916
rect 29820 34802 29876 34804
rect 29820 34750 29822 34802
rect 29822 34750 29874 34802
rect 29874 34750 29876 34802
rect 29820 34748 29876 34750
rect 29596 34690 29652 34692
rect 29596 34638 29598 34690
rect 29598 34638 29650 34690
rect 29650 34638 29652 34690
rect 29596 34636 29652 34638
rect 28812 33628 28868 33684
rect 28924 33292 28980 33348
rect 28700 33068 28756 33124
rect 29372 33068 29428 33124
rect 26796 31890 26852 31892
rect 26796 31838 26798 31890
rect 26798 31838 26850 31890
rect 26850 31838 26852 31890
rect 26796 31836 26852 31838
rect 28812 31612 28868 31668
rect 28140 30156 28196 30212
rect 26460 29260 26516 29316
rect 26908 29650 26964 29652
rect 26908 29598 26910 29650
rect 26910 29598 26962 29650
rect 26962 29598 26964 29650
rect 26908 29596 26964 29598
rect 26348 29036 26404 29092
rect 27804 29650 27860 29652
rect 27804 29598 27806 29650
rect 27806 29598 27858 29650
rect 27858 29598 27860 29650
rect 27804 29596 27860 29598
rect 28028 29650 28084 29652
rect 28028 29598 28030 29650
rect 28030 29598 28082 29650
rect 28082 29598 28084 29650
rect 28028 29596 28084 29598
rect 27692 29538 27748 29540
rect 27692 29486 27694 29538
rect 27694 29486 27746 29538
rect 27746 29486 27748 29538
rect 27692 29484 27748 29486
rect 27580 29372 27636 29428
rect 27692 29314 27748 29316
rect 27692 29262 27694 29314
rect 27694 29262 27746 29314
rect 27746 29262 27748 29314
rect 27692 29260 27748 29262
rect 29708 30828 29764 30884
rect 29596 30268 29652 30324
rect 29036 29596 29092 29652
rect 28476 29538 28532 29540
rect 28476 29486 28478 29538
rect 28478 29486 28530 29538
rect 28530 29486 28532 29538
rect 28476 29484 28532 29486
rect 28140 29260 28196 29316
rect 26908 28924 26964 28980
rect 28364 28812 28420 28868
rect 28252 28082 28308 28084
rect 28252 28030 28254 28082
rect 28254 28030 28306 28082
rect 28306 28030 28308 28082
rect 28252 28028 28308 28030
rect 24668 25564 24724 25620
rect 24780 26796 24836 26852
rect 24668 25394 24724 25396
rect 24668 25342 24670 25394
rect 24670 25342 24722 25394
rect 24722 25342 24724 25394
rect 24668 25340 24724 25342
rect 26348 27020 26404 27076
rect 26796 27074 26852 27076
rect 26796 27022 26798 27074
rect 26798 27022 26850 27074
rect 26850 27022 26852 27074
rect 26796 27020 26852 27022
rect 28028 27074 28084 27076
rect 28028 27022 28030 27074
rect 28030 27022 28082 27074
rect 28082 27022 28084 27074
rect 28028 27020 28084 27022
rect 24444 25228 24500 25284
rect 24332 23826 24388 23828
rect 24332 23774 24334 23826
rect 24334 23774 24386 23826
rect 24386 23774 24388 23826
rect 24332 23772 24388 23774
rect 23436 23378 23492 23380
rect 23436 23326 23438 23378
rect 23438 23326 23490 23378
rect 23490 23326 23492 23378
rect 23436 23324 23492 23326
rect 23996 23324 24052 23380
rect 23884 22258 23940 22260
rect 23884 22206 23886 22258
rect 23886 22206 23938 22258
rect 23938 22206 23940 22258
rect 23884 22204 23940 22206
rect 24892 23548 24948 23604
rect 24220 23154 24276 23156
rect 24220 23102 24222 23154
rect 24222 23102 24274 23154
rect 24274 23102 24276 23154
rect 24220 23100 24276 23102
rect 24444 23100 24500 23156
rect 24108 22204 24164 22260
rect 23996 21532 24052 21588
rect 24892 21532 24948 21588
rect 23660 19234 23716 19236
rect 23660 19182 23662 19234
rect 23662 19182 23714 19234
rect 23714 19182 23716 19234
rect 23660 19180 23716 19182
rect 24332 19234 24388 19236
rect 24332 19182 24334 19234
rect 24334 19182 24386 19234
rect 24386 19182 24388 19234
rect 24332 19180 24388 19182
rect 25340 26796 25396 26852
rect 25116 26514 25172 26516
rect 25116 26462 25118 26514
rect 25118 26462 25170 26514
rect 25170 26462 25172 26514
rect 25116 26460 25172 26462
rect 25452 26684 25508 26740
rect 25900 26460 25956 26516
rect 26236 26348 26292 26404
rect 26124 26290 26180 26292
rect 26124 26238 26126 26290
rect 26126 26238 26178 26290
rect 26178 26238 26180 26290
rect 26124 26236 26180 26238
rect 26572 26850 26628 26852
rect 26572 26798 26574 26850
rect 26574 26798 26626 26850
rect 26626 26798 26628 26850
rect 26572 26796 26628 26798
rect 27020 26460 27076 26516
rect 25564 25676 25620 25732
rect 26124 26012 26180 26068
rect 25900 25676 25956 25732
rect 26012 25900 26068 25956
rect 25228 24556 25284 24612
rect 25340 23772 25396 23828
rect 25228 23154 25284 23156
rect 25228 23102 25230 23154
rect 25230 23102 25282 23154
rect 25282 23102 25284 23154
rect 25228 23100 25284 23102
rect 25228 22204 25284 22260
rect 26348 26012 26404 26068
rect 26572 26290 26628 26292
rect 26572 26238 26574 26290
rect 26574 26238 26626 26290
rect 26626 26238 26628 26290
rect 26572 26236 26628 26238
rect 26572 25900 26628 25956
rect 26908 26124 26964 26180
rect 26124 25618 26180 25620
rect 26124 25566 26126 25618
rect 26126 25566 26178 25618
rect 26178 25566 26180 25618
rect 26124 25564 26180 25566
rect 26348 25564 26404 25620
rect 25900 25340 25956 25396
rect 25564 24946 25620 24948
rect 25564 24894 25566 24946
rect 25566 24894 25618 24946
rect 25618 24894 25620 24946
rect 25564 24892 25620 24894
rect 25788 24556 25844 24612
rect 25900 23772 25956 23828
rect 26348 24444 26404 24500
rect 25340 21810 25396 21812
rect 25340 21758 25342 21810
rect 25342 21758 25394 21810
rect 25394 21758 25396 21810
rect 25340 21756 25396 21758
rect 26684 25788 26740 25844
rect 26908 25564 26964 25620
rect 27356 26514 27412 26516
rect 27356 26462 27358 26514
rect 27358 26462 27410 26514
rect 27410 26462 27412 26514
rect 27356 26460 27412 26462
rect 28700 27020 28756 27076
rect 30828 39004 30884 39060
rect 30828 38610 30884 38612
rect 30828 38558 30830 38610
rect 30830 38558 30882 38610
rect 30882 38558 30884 38610
rect 30828 38556 30884 38558
rect 31276 37436 31332 37492
rect 30492 35698 30548 35700
rect 30492 35646 30494 35698
rect 30494 35646 30546 35698
rect 30546 35646 30548 35698
rect 30492 35644 30548 35646
rect 30268 34914 30324 34916
rect 30268 34862 30270 34914
rect 30270 34862 30322 34914
rect 30322 34862 30324 34914
rect 30268 34860 30324 34862
rect 30268 34636 30324 34692
rect 30268 34076 30324 34132
rect 30380 33180 30436 33236
rect 30940 34972 30996 35028
rect 30716 34748 30772 34804
rect 31164 36258 31220 36260
rect 31164 36206 31166 36258
rect 31166 36206 31218 36258
rect 31218 36206 31220 36258
rect 31164 36204 31220 36206
rect 31948 46172 32004 46228
rect 31836 45218 31892 45220
rect 31836 45166 31838 45218
rect 31838 45166 31890 45218
rect 31890 45166 31892 45218
rect 31836 45164 31892 45166
rect 32060 45724 32116 45780
rect 31836 44268 31892 44324
rect 32172 44156 32228 44212
rect 32172 41916 32228 41972
rect 31612 39340 31668 39396
rect 32956 49138 33012 49140
rect 32956 49086 32958 49138
rect 32958 49086 33010 49138
rect 33010 49086 33012 49138
rect 32956 49084 33012 49086
rect 33292 52444 33348 52500
rect 33180 52332 33236 52388
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 36764 62188 36820 62244
rect 34524 61180 34580 61236
rect 34412 61068 34468 61124
rect 33852 60844 33908 60900
rect 34748 60844 34804 60900
rect 34748 60508 34804 60564
rect 34972 61068 35028 61124
rect 34860 59164 34916 59220
rect 35196 61180 35252 61236
rect 35420 60898 35476 60900
rect 35420 60846 35422 60898
rect 35422 60846 35474 60898
rect 35474 60846 35476 60898
rect 35420 60844 35476 60846
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 36092 61180 36148 61236
rect 35868 61068 35924 61124
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 36988 60508 37044 60564
rect 38220 62412 38276 62468
rect 33740 57596 33796 57652
rect 35532 57708 35588 57764
rect 34972 57372 35028 57428
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 33740 56978 33796 56980
rect 33740 56926 33742 56978
rect 33742 56926 33794 56978
rect 33794 56926 33796 56978
rect 33740 56924 33796 56926
rect 35196 56700 35252 56756
rect 33628 55356 33684 55412
rect 33516 52444 33572 52500
rect 36204 57708 36260 57764
rect 35644 56194 35700 56196
rect 35644 56142 35646 56194
rect 35646 56142 35698 56194
rect 35698 56142 35700 56194
rect 35644 56140 35700 56142
rect 36092 56754 36148 56756
rect 36092 56702 36094 56754
rect 36094 56702 36146 56754
rect 36146 56702 36148 56754
rect 36092 56700 36148 56702
rect 36428 56812 36484 56868
rect 36204 56140 36260 56196
rect 35980 56028 36036 56084
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35196 55522 35252 55524
rect 35196 55470 35198 55522
rect 35198 55470 35250 55522
rect 35250 55470 35252 55522
rect 35196 55468 35252 55470
rect 35980 55468 36036 55524
rect 34860 55410 34916 55412
rect 34860 55358 34862 55410
rect 34862 55358 34914 55410
rect 34914 55358 34916 55410
rect 34860 55356 34916 55358
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 37100 59218 37156 59220
rect 37100 59166 37102 59218
rect 37102 59166 37154 59218
rect 37154 59166 37156 59218
rect 37100 59164 37156 59166
rect 39452 62466 39508 62468
rect 39452 62414 39454 62466
rect 39454 62414 39506 62466
rect 39506 62414 39508 62466
rect 39452 62412 39508 62414
rect 37324 61010 37380 61012
rect 37324 60958 37326 61010
rect 37326 60958 37378 61010
rect 37378 60958 37380 61010
rect 37324 60956 37380 60958
rect 37548 60844 37604 60900
rect 37772 61292 37828 61348
rect 38332 61346 38388 61348
rect 38332 61294 38334 61346
rect 38334 61294 38386 61346
rect 38386 61294 38388 61346
rect 38332 61292 38388 61294
rect 37772 60844 37828 60900
rect 37884 60956 37940 61012
rect 38668 61068 38724 61124
rect 39116 60898 39172 60900
rect 39116 60846 39118 60898
rect 39118 60846 39170 60898
rect 39170 60846 39172 60898
rect 39116 60844 39172 60846
rect 38108 60060 38164 60116
rect 37772 58492 37828 58548
rect 37660 57708 37716 57764
rect 37772 57372 37828 57428
rect 36876 57036 36932 57092
rect 34524 53730 34580 53732
rect 34524 53678 34526 53730
rect 34526 53678 34578 53730
rect 34578 53678 34580 53730
rect 34524 53676 34580 53678
rect 35980 53116 36036 53172
rect 35644 53004 35700 53060
rect 34412 52946 34468 52948
rect 34412 52894 34414 52946
rect 34414 52894 34466 52946
rect 34466 52894 34468 52946
rect 34412 52892 34468 52894
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 33740 52220 33796 52276
rect 35644 52332 35700 52388
rect 33852 52108 33908 52164
rect 33404 49810 33460 49812
rect 33404 49758 33406 49810
rect 33406 49758 33458 49810
rect 33458 49758 33460 49810
rect 33404 49756 33460 49758
rect 32508 46898 32564 46900
rect 32508 46846 32510 46898
rect 32510 46846 32562 46898
rect 32562 46846 32564 46898
rect 32508 46844 32564 46846
rect 33180 45778 33236 45780
rect 33180 45726 33182 45778
rect 33182 45726 33234 45778
rect 33234 45726 33236 45778
rect 33180 45724 33236 45726
rect 32620 44322 32676 44324
rect 32620 44270 32622 44322
rect 32622 44270 32674 44322
rect 32674 44270 32676 44322
rect 32620 44268 32676 44270
rect 33292 44268 33348 44324
rect 33068 44210 33124 44212
rect 33068 44158 33070 44210
rect 33070 44158 33122 44210
rect 33122 44158 33124 44210
rect 33068 44156 33124 44158
rect 33740 49138 33796 49140
rect 33740 49086 33742 49138
rect 33742 49086 33794 49138
rect 33794 49086 33796 49138
rect 33740 49084 33796 49086
rect 33628 44156 33684 44212
rect 33628 43932 33684 43988
rect 32620 43036 32676 43092
rect 33516 43036 33572 43092
rect 35980 52946 36036 52948
rect 35980 52894 35982 52946
rect 35982 52894 36034 52946
rect 36034 52894 36036 52946
rect 35980 52892 36036 52894
rect 36204 53788 36260 53844
rect 36428 53676 36484 53732
rect 36316 53116 36372 53172
rect 36652 53058 36708 53060
rect 36652 53006 36654 53058
rect 36654 53006 36706 53058
rect 36706 53006 36708 53058
rect 36652 53004 36708 53006
rect 36764 52946 36820 52948
rect 36764 52894 36766 52946
rect 36766 52894 36818 52946
rect 36818 52894 36820 52946
rect 36764 52892 36820 52894
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 34188 49756 34244 49812
rect 36764 51212 36820 51268
rect 36092 51100 36148 51156
rect 35084 49810 35140 49812
rect 35084 49758 35086 49810
rect 35086 49758 35138 49810
rect 35138 49758 35140 49810
rect 35084 49756 35140 49758
rect 34860 49420 34916 49476
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35084 48972 35140 49028
rect 34636 47570 34692 47572
rect 34636 47518 34638 47570
rect 34638 47518 34690 47570
rect 34690 47518 34692 47570
rect 34636 47516 34692 47518
rect 34972 47516 35028 47572
rect 34748 46786 34804 46788
rect 34748 46734 34750 46786
rect 34750 46734 34802 46786
rect 34802 46734 34804 46786
rect 34748 46732 34804 46734
rect 34412 45276 34468 45332
rect 34076 45164 34132 45220
rect 33964 44940 34020 44996
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35420 47682 35476 47684
rect 35420 47630 35422 47682
rect 35422 47630 35474 47682
rect 35474 47630 35476 47682
rect 35420 47628 35476 47630
rect 35868 46620 35924 46676
rect 35756 46396 35812 46452
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35420 44994 35476 44996
rect 35420 44942 35422 44994
rect 35422 44942 35474 44994
rect 35474 44942 35476 44994
rect 35420 44940 35476 44942
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35644 44434 35700 44436
rect 35644 44382 35646 44434
rect 35646 44382 35698 44434
rect 35698 44382 35700 44434
rect 35644 44380 35700 44382
rect 34076 44210 34132 44212
rect 34076 44158 34078 44210
rect 34078 44158 34130 44210
rect 34130 44158 34132 44210
rect 34076 44156 34132 44158
rect 34636 44098 34692 44100
rect 34636 44046 34638 44098
rect 34638 44046 34690 44098
rect 34690 44046 34692 44098
rect 34636 44044 34692 44046
rect 34860 44098 34916 44100
rect 34860 44046 34862 44098
rect 34862 44046 34914 44098
rect 34914 44046 34916 44098
rect 34860 44044 34916 44046
rect 33628 42364 33684 42420
rect 35084 43708 35140 43764
rect 36652 47628 36708 47684
rect 36428 47404 36484 47460
rect 36092 47292 36148 47348
rect 36652 46674 36708 46676
rect 36652 46622 36654 46674
rect 36654 46622 36706 46674
rect 36706 46622 36708 46674
rect 36652 46620 36708 46622
rect 36316 46450 36372 46452
rect 36316 46398 36318 46450
rect 36318 46398 36370 46450
rect 36370 46398 36372 46450
rect 36316 46396 36372 46398
rect 36204 45276 36260 45332
rect 36652 45330 36708 45332
rect 36652 45278 36654 45330
rect 36654 45278 36706 45330
rect 36706 45278 36708 45330
rect 36652 45276 36708 45278
rect 37100 56866 37156 56868
rect 37100 56814 37102 56866
rect 37102 56814 37154 56866
rect 37154 56814 37156 56866
rect 37100 56812 37156 56814
rect 37324 56700 37380 56756
rect 37100 56140 37156 56196
rect 37212 56082 37268 56084
rect 37212 56030 37214 56082
rect 37214 56030 37266 56082
rect 37266 56030 37268 56082
rect 37212 56028 37268 56030
rect 37996 56866 38052 56868
rect 37996 56814 37998 56866
rect 37998 56814 38050 56866
rect 38050 56814 38052 56866
rect 37996 56812 38052 56814
rect 37100 53842 37156 53844
rect 37100 53790 37102 53842
rect 37102 53790 37154 53842
rect 37154 53790 37156 53842
rect 37100 53788 37156 53790
rect 37996 53788 38052 53844
rect 37324 53116 37380 53172
rect 37772 51266 37828 51268
rect 37772 51214 37774 51266
rect 37774 51214 37826 51266
rect 37826 51214 37828 51266
rect 37772 51212 37828 51214
rect 39452 59612 39508 59668
rect 39228 59052 39284 59108
rect 38556 58492 38612 58548
rect 39900 61292 39956 61348
rect 40012 60732 40068 60788
rect 39900 60508 39956 60564
rect 40012 59778 40068 59780
rect 40012 59726 40014 59778
rect 40014 59726 40066 59778
rect 40066 59726 40068 59778
rect 40012 59724 40068 59726
rect 38220 56700 38276 56756
rect 39004 56082 39060 56084
rect 39004 56030 39006 56082
rect 39006 56030 39058 56082
rect 39058 56030 39060 56082
rect 39004 56028 39060 56030
rect 38332 55186 38388 55188
rect 38332 55134 38334 55186
rect 38334 55134 38386 55186
rect 38386 55134 38388 55186
rect 38332 55132 38388 55134
rect 39564 55132 39620 55188
rect 39452 54626 39508 54628
rect 39452 54574 39454 54626
rect 39454 54574 39506 54626
rect 39506 54574 39508 54626
rect 39452 54572 39508 54574
rect 39564 53618 39620 53620
rect 39564 53566 39566 53618
rect 39566 53566 39618 53618
rect 39618 53566 39620 53618
rect 39564 53564 39620 53566
rect 38556 53004 38612 53060
rect 38556 51212 38612 51268
rect 37772 49922 37828 49924
rect 37772 49870 37774 49922
rect 37774 49870 37826 49922
rect 37826 49870 37828 49922
rect 37772 49868 37828 49870
rect 37436 47628 37492 47684
rect 38108 47516 38164 47572
rect 37100 47180 37156 47236
rect 37660 47180 37716 47236
rect 37548 46844 37604 46900
rect 38556 49868 38612 49924
rect 39340 49980 39396 50036
rect 39900 54572 39956 54628
rect 41580 64146 41636 64148
rect 41580 64094 41582 64146
rect 41582 64094 41634 64146
rect 41634 64094 41636 64146
rect 41580 64092 41636 64094
rect 41020 63026 41076 63028
rect 41020 62974 41022 63026
rect 41022 62974 41074 63026
rect 41074 62974 41076 63026
rect 41020 62972 41076 62974
rect 42028 65324 42084 65380
rect 41804 62972 41860 63028
rect 41916 62860 41972 62916
rect 41244 62354 41300 62356
rect 41244 62302 41246 62354
rect 41246 62302 41298 62354
rect 41298 62302 41300 62354
rect 41244 62300 41300 62302
rect 41020 62242 41076 62244
rect 41020 62190 41022 62242
rect 41022 62190 41074 62242
rect 41074 62190 41076 62242
rect 41020 62188 41076 62190
rect 42028 61404 42084 61460
rect 40460 60620 40516 60676
rect 41468 60562 41524 60564
rect 41468 60510 41470 60562
rect 41470 60510 41522 60562
rect 41522 60510 41524 60562
rect 41468 60508 41524 60510
rect 40348 58940 40404 58996
rect 40684 59500 40740 59556
rect 41244 59218 41300 59220
rect 41244 59166 41246 59218
rect 41246 59166 41298 59218
rect 41298 59166 41300 59218
rect 41244 59164 41300 59166
rect 41916 60674 41972 60676
rect 41916 60622 41918 60674
rect 41918 60622 41970 60674
rect 41970 60622 41972 60674
rect 41916 60620 41972 60622
rect 41804 60508 41860 60564
rect 41020 59106 41076 59108
rect 41020 59054 41022 59106
rect 41022 59054 41074 59106
rect 41074 59054 41076 59106
rect 41020 59052 41076 59054
rect 41692 59724 41748 59780
rect 40796 58940 40852 58996
rect 41020 58492 41076 58548
rect 40460 55020 40516 55076
rect 40124 53900 40180 53956
rect 40796 54572 40852 54628
rect 41916 59612 41972 59668
rect 43372 63922 43428 63924
rect 43372 63870 43374 63922
rect 43374 63870 43426 63922
rect 43426 63870 43428 63922
rect 43372 63868 43428 63870
rect 44380 65324 44436 65380
rect 44940 64204 44996 64260
rect 44828 63980 44884 64036
rect 42252 62188 42308 62244
rect 42924 62914 42980 62916
rect 42924 62862 42926 62914
rect 42926 62862 42978 62914
rect 42978 62862 42980 62914
rect 42924 62860 42980 62862
rect 43820 63922 43876 63924
rect 43820 63870 43822 63922
rect 43822 63870 43874 63922
rect 43874 63870 43876 63922
rect 43820 63868 43876 63870
rect 43484 63138 43540 63140
rect 43484 63086 43486 63138
rect 43486 63086 43538 63138
rect 43538 63086 43540 63138
rect 43484 63084 43540 63086
rect 42700 62300 42756 62356
rect 43484 62354 43540 62356
rect 43484 62302 43486 62354
rect 43486 62302 43538 62354
rect 43538 62302 43540 62354
rect 43484 62300 43540 62302
rect 43596 62188 43652 62244
rect 43708 61458 43764 61460
rect 43708 61406 43710 61458
rect 43710 61406 43762 61458
rect 43762 61406 43764 61458
rect 43708 61404 43764 61406
rect 42476 60508 42532 60564
rect 42364 59330 42420 59332
rect 42364 59278 42366 59330
rect 42366 59278 42418 59330
rect 42418 59278 42420 59330
rect 42364 59276 42420 59278
rect 41804 58546 41860 58548
rect 41804 58494 41806 58546
rect 41806 58494 41858 58546
rect 41858 58494 41860 58546
rect 41804 58492 41860 58494
rect 42812 59612 42868 59668
rect 43036 59330 43092 59332
rect 43036 59278 43038 59330
rect 43038 59278 43090 59330
rect 43090 59278 43092 59330
rect 43036 59276 43092 59278
rect 42364 58492 42420 58548
rect 43260 59218 43316 59220
rect 43260 59166 43262 59218
rect 43262 59166 43314 59218
rect 43314 59166 43316 59218
rect 43260 59164 43316 59166
rect 44044 63138 44100 63140
rect 44044 63086 44046 63138
rect 44046 63086 44098 63138
rect 44098 63086 44100 63138
rect 44044 63084 44100 63086
rect 44156 63026 44212 63028
rect 44156 62974 44158 63026
rect 44158 62974 44210 63026
rect 44210 62974 44212 63026
rect 44156 62972 44212 62974
rect 43932 62354 43988 62356
rect 43932 62302 43934 62354
rect 43934 62302 43986 62354
rect 43986 62302 43988 62354
rect 43932 62300 43988 62302
rect 45164 63868 45220 63924
rect 45612 64092 45668 64148
rect 44940 63138 44996 63140
rect 44940 63086 44942 63138
rect 44942 63086 44994 63138
rect 44994 63086 44996 63138
rect 44940 63084 44996 63086
rect 45052 63026 45108 63028
rect 45052 62974 45054 63026
rect 45054 62974 45106 63026
rect 45106 62974 45108 63026
rect 45052 62972 45108 62974
rect 45276 62914 45332 62916
rect 45276 62862 45278 62914
rect 45278 62862 45330 62914
rect 45330 62862 45332 62914
rect 45276 62860 45332 62862
rect 44940 62354 44996 62356
rect 44940 62302 44942 62354
rect 44942 62302 44994 62354
rect 44994 62302 44996 62354
rect 44940 62300 44996 62302
rect 46060 63138 46116 63140
rect 46060 63086 46062 63138
rect 46062 63086 46114 63138
rect 46114 63086 46116 63138
rect 46060 63084 46116 63086
rect 46508 65324 46564 65380
rect 46508 64092 46564 64148
rect 46396 63922 46452 63924
rect 46396 63870 46398 63922
rect 46398 63870 46450 63922
rect 46450 63870 46452 63922
rect 46396 63868 46452 63870
rect 46732 64146 46788 64148
rect 46732 64094 46734 64146
rect 46734 64094 46786 64146
rect 46786 64094 46788 64146
rect 46732 64092 46788 64094
rect 46844 64034 46900 64036
rect 46844 63982 46846 64034
rect 46846 63982 46898 64034
rect 46898 63982 46900 64034
rect 46844 63980 46900 63982
rect 45612 62578 45668 62580
rect 45612 62526 45614 62578
rect 45614 62526 45666 62578
rect 45666 62526 45668 62578
rect 45612 62524 45668 62526
rect 44156 61404 44212 61460
rect 45724 62354 45780 62356
rect 45724 62302 45726 62354
rect 45726 62302 45778 62354
rect 45778 62302 45780 62354
rect 45724 62300 45780 62302
rect 46508 62524 46564 62580
rect 47292 63084 47348 63140
rect 47180 62914 47236 62916
rect 47180 62862 47182 62914
rect 47182 62862 47234 62914
rect 47234 62862 47236 62914
rect 47180 62860 47236 62862
rect 48412 66498 48468 66500
rect 48412 66446 48414 66498
rect 48414 66446 48466 66498
rect 48466 66446 48468 66498
rect 48412 66444 48468 66446
rect 49084 66444 49140 66500
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 52220 66498 52276 66500
rect 52220 66446 52222 66498
rect 52222 66446 52274 66498
rect 52274 66446 52276 66498
rect 52220 66444 52276 66446
rect 53116 66444 53172 66500
rect 51100 65548 51156 65604
rect 47740 65378 47796 65380
rect 47740 65326 47742 65378
rect 47742 65326 47794 65378
rect 47794 65326 47796 65378
rect 47740 65324 47796 65326
rect 47516 64316 47572 64372
rect 44940 60620 44996 60676
rect 44268 60226 44324 60228
rect 44268 60174 44270 60226
rect 44270 60174 44322 60226
rect 44322 60174 44324 60226
rect 44268 60172 44324 60174
rect 44156 59612 44212 59668
rect 43820 59164 43876 59220
rect 45276 59218 45332 59220
rect 45276 59166 45278 59218
rect 45278 59166 45330 59218
rect 45330 59166 45332 59218
rect 45276 59164 45332 59166
rect 43260 58716 43316 58772
rect 41692 58268 41748 58324
rect 43148 58380 43204 58436
rect 42588 57538 42644 57540
rect 42588 57486 42590 57538
rect 42590 57486 42642 57538
rect 42642 57486 42644 57538
rect 42588 57484 42644 57486
rect 44828 58380 44884 58436
rect 45724 58828 45780 58884
rect 45276 58492 45332 58548
rect 43148 57538 43204 57540
rect 43148 57486 43150 57538
rect 43150 57486 43202 57538
rect 43202 57486 43204 57538
rect 43148 57484 43204 57486
rect 43596 57596 43652 57652
rect 42252 56866 42308 56868
rect 42252 56814 42254 56866
rect 42254 56814 42306 56866
rect 42306 56814 42308 56866
rect 42252 56812 42308 56814
rect 42924 56700 42980 56756
rect 41692 55916 41748 55972
rect 41580 55410 41636 55412
rect 41580 55358 41582 55410
rect 41582 55358 41634 55410
rect 41634 55358 41636 55410
rect 41580 55356 41636 55358
rect 41468 55020 41524 55076
rect 41020 54012 41076 54068
rect 40124 53506 40180 53508
rect 40124 53454 40126 53506
rect 40126 53454 40178 53506
rect 40178 53454 40180 53506
rect 40124 53452 40180 53454
rect 39676 49308 39732 49364
rect 42924 55916 42980 55972
rect 43260 56754 43316 56756
rect 43260 56702 43262 56754
rect 43262 56702 43314 56754
rect 43314 56702 43316 56754
rect 43260 56700 43316 56702
rect 44492 57650 44548 57652
rect 44492 57598 44494 57650
rect 44494 57598 44546 57650
rect 44546 57598 44548 57650
rect 44492 57596 44548 57598
rect 45500 55970 45556 55972
rect 45500 55918 45502 55970
rect 45502 55918 45554 55970
rect 45554 55918 45556 55970
rect 45500 55916 45556 55918
rect 42140 55410 42196 55412
rect 42140 55358 42142 55410
rect 42142 55358 42194 55410
rect 42194 55358 42196 55410
rect 42140 55356 42196 55358
rect 41804 54738 41860 54740
rect 41804 54686 41806 54738
rect 41806 54686 41858 54738
rect 41858 54686 41860 54738
rect 41804 54684 41860 54686
rect 44268 55244 44324 55300
rect 42364 55020 42420 55076
rect 44940 55298 44996 55300
rect 44940 55246 44942 55298
rect 44942 55246 44994 55298
rect 44994 55246 44996 55298
rect 44940 55244 44996 55246
rect 47068 59388 47124 59444
rect 46956 58546 47012 58548
rect 46956 58494 46958 58546
rect 46958 58494 47010 58546
rect 47010 58494 47012 58546
rect 46956 58492 47012 58494
rect 47068 57372 47124 57428
rect 47740 63532 47796 63588
rect 47740 63084 47796 63140
rect 48860 62524 48916 62580
rect 49532 64204 49588 64260
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 52332 65436 52388 65492
rect 49532 63922 49588 63924
rect 49532 63870 49534 63922
rect 49534 63870 49586 63922
rect 49586 63870 49588 63922
rect 49532 63868 49588 63870
rect 49980 63196 50036 63252
rect 49644 63084 49700 63140
rect 48860 61852 48916 61908
rect 48860 60172 48916 60228
rect 50092 62188 50148 62244
rect 49084 61010 49140 61012
rect 49084 60958 49086 61010
rect 49086 60958 49138 61010
rect 49138 60958 49140 61010
rect 49084 60956 49140 60958
rect 48300 59388 48356 59444
rect 48188 59330 48244 59332
rect 48188 59278 48190 59330
rect 48190 59278 48242 59330
rect 48242 59278 48244 59330
rect 48188 59276 48244 59278
rect 49756 60956 49812 61012
rect 48860 58716 48916 58772
rect 49532 60620 49588 60676
rect 50652 63532 50708 63588
rect 50764 63138 50820 63140
rect 50764 63086 50766 63138
rect 50766 63086 50818 63138
rect 50818 63086 50820 63138
rect 50764 63084 50820 63086
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 51772 65324 51828 65380
rect 50988 61852 51044 61908
rect 51100 63196 51156 63252
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50428 60956 50484 61012
rect 50988 61010 51044 61012
rect 50988 60958 50990 61010
rect 50990 60958 51042 61010
rect 51042 60958 51044 61010
rect 50988 60956 51044 60958
rect 50204 60844 50260 60900
rect 49756 60674 49812 60676
rect 49756 60622 49758 60674
rect 49758 60622 49810 60674
rect 49810 60622 49812 60674
rect 49756 60620 49812 60622
rect 49532 59276 49588 59332
rect 48188 57372 48244 57428
rect 47628 56252 47684 56308
rect 46396 55916 46452 55972
rect 42476 54738 42532 54740
rect 42476 54686 42478 54738
rect 42478 54686 42530 54738
rect 42530 54686 42532 54738
rect 42476 54684 42532 54686
rect 40908 53618 40964 53620
rect 40908 53566 40910 53618
rect 40910 53566 40962 53618
rect 40962 53566 40964 53618
rect 40908 53564 40964 53566
rect 42028 53788 42084 53844
rect 42476 54012 42532 54068
rect 41356 53506 41412 53508
rect 41356 53454 41358 53506
rect 41358 53454 41410 53506
rect 41410 53454 41412 53506
rect 41356 53452 41412 53454
rect 41020 53004 41076 53060
rect 38444 47458 38500 47460
rect 38444 47406 38446 47458
rect 38446 47406 38498 47458
rect 38498 47406 38500 47458
rect 38444 47404 38500 47406
rect 39004 47292 39060 47348
rect 38556 47234 38612 47236
rect 38556 47182 38558 47234
rect 38558 47182 38610 47234
rect 38610 47182 38612 47234
rect 38556 47180 38612 47182
rect 38332 46844 38388 46900
rect 37436 46620 37492 46676
rect 37100 46396 37156 46452
rect 33628 42194 33684 42196
rect 33628 42142 33630 42194
rect 33630 42142 33682 42194
rect 33682 42142 33684 42194
rect 33628 42140 33684 42142
rect 33740 42028 33796 42084
rect 33852 43484 33908 43540
rect 33404 41746 33460 41748
rect 33404 41694 33406 41746
rect 33406 41694 33458 41746
rect 33458 41694 33460 41746
rect 33404 41692 33460 41694
rect 32508 41298 32564 41300
rect 32508 41246 32510 41298
rect 32510 41246 32562 41298
rect 32562 41246 32564 41298
rect 32508 41244 32564 41246
rect 33180 41186 33236 41188
rect 33180 41134 33182 41186
rect 33182 41134 33234 41186
rect 33234 41134 33236 41186
rect 33180 41132 33236 41134
rect 32060 39004 32116 39060
rect 31500 37884 31556 37940
rect 31948 38444 32004 38500
rect 31500 37100 31556 37156
rect 31052 34748 31108 34804
rect 31164 35532 31220 35588
rect 30940 34076 30996 34132
rect 30828 31890 30884 31892
rect 30828 31838 30830 31890
rect 30830 31838 30882 31890
rect 30882 31838 30884 31890
rect 30828 31836 30884 31838
rect 30604 31612 30660 31668
rect 31500 35196 31556 35252
rect 31612 34972 31668 35028
rect 31836 34130 31892 34132
rect 31836 34078 31838 34130
rect 31838 34078 31890 34130
rect 31890 34078 31892 34130
rect 31836 34076 31892 34078
rect 31836 33852 31892 33908
rect 31836 32620 31892 32676
rect 31276 31836 31332 31892
rect 30044 30268 30100 30324
rect 31276 30156 31332 30212
rect 30492 30098 30548 30100
rect 30492 30046 30494 30098
rect 30494 30046 30546 30098
rect 30546 30046 30548 30098
rect 30492 30044 30548 30046
rect 29932 29596 29988 29652
rect 29484 29484 29540 29540
rect 29708 29314 29764 29316
rect 29708 29262 29710 29314
rect 29710 29262 29762 29314
rect 29762 29262 29764 29314
rect 29708 29260 29764 29262
rect 29708 28588 29764 28644
rect 31164 30098 31220 30100
rect 31164 30046 31166 30098
rect 31166 30046 31218 30098
rect 31218 30046 31220 30098
rect 31164 30044 31220 30046
rect 30604 29596 30660 29652
rect 30716 29036 30772 29092
rect 30604 28812 30660 28868
rect 30380 28700 30436 28756
rect 30268 28642 30324 28644
rect 30268 28590 30270 28642
rect 30270 28590 30322 28642
rect 30322 28590 30324 28642
rect 30268 28588 30324 28590
rect 32620 36988 32676 37044
rect 32060 36204 32116 36260
rect 32172 32732 32228 32788
rect 33068 37772 33124 37828
rect 33068 37212 33124 37268
rect 33404 37266 33460 37268
rect 33404 37214 33406 37266
rect 33406 37214 33458 37266
rect 33458 37214 33460 37266
rect 33404 37212 33460 37214
rect 33404 36876 33460 36932
rect 33292 36594 33348 36596
rect 33292 36542 33294 36594
rect 33294 36542 33346 36594
rect 33346 36542 33348 36594
rect 33292 36540 33348 36542
rect 32284 32620 32340 32676
rect 32284 32060 32340 32116
rect 32508 31836 32564 31892
rect 33292 35308 33348 35364
rect 33180 32786 33236 32788
rect 33180 32734 33182 32786
rect 33182 32734 33234 32786
rect 33234 32734 33236 32786
rect 33180 32732 33236 32734
rect 32956 31778 33012 31780
rect 32956 31726 32958 31778
rect 32958 31726 33010 31778
rect 33010 31726 33012 31778
rect 32956 31724 33012 31726
rect 31612 29596 31668 29652
rect 31276 29538 31332 29540
rect 31276 29486 31278 29538
rect 31278 29486 31330 29538
rect 31330 29486 31332 29538
rect 31276 29484 31332 29486
rect 30940 29260 30996 29316
rect 31388 29036 31444 29092
rect 31164 28642 31220 28644
rect 31164 28590 31166 28642
rect 31166 28590 31218 28642
rect 31218 28590 31220 28642
rect 31164 28588 31220 28590
rect 30380 27916 30436 27972
rect 27804 26460 27860 26516
rect 28476 26514 28532 26516
rect 28476 26462 28478 26514
rect 28478 26462 28530 26514
rect 28530 26462 28532 26514
rect 28476 26460 28532 26462
rect 27468 26348 27524 26404
rect 28812 26402 28868 26404
rect 28812 26350 28814 26402
rect 28814 26350 28866 26402
rect 28866 26350 28868 26402
rect 28812 26348 28868 26350
rect 28252 26290 28308 26292
rect 28252 26238 28254 26290
rect 28254 26238 28306 26290
rect 28306 26238 28308 26290
rect 28252 26236 28308 26238
rect 28588 26290 28644 26292
rect 28588 26238 28590 26290
rect 28590 26238 28642 26290
rect 28642 26238 28644 26290
rect 28588 26236 28644 26238
rect 27804 25676 27860 25732
rect 27692 25618 27748 25620
rect 27692 25566 27694 25618
rect 27694 25566 27746 25618
rect 27746 25566 27748 25618
rect 27692 25564 27748 25566
rect 27916 25564 27972 25620
rect 27244 25452 27300 25508
rect 28588 25618 28644 25620
rect 28588 25566 28590 25618
rect 28590 25566 28642 25618
rect 28642 25566 28644 25618
rect 28588 25564 28644 25566
rect 27132 25340 27188 25396
rect 27356 24892 27412 24948
rect 28028 25228 28084 25284
rect 27692 24892 27748 24948
rect 27020 24444 27076 24500
rect 26796 23212 26852 23268
rect 26908 23548 26964 23604
rect 27580 23378 27636 23380
rect 27580 23326 27582 23378
rect 27582 23326 27634 23378
rect 27634 23326 27636 23378
rect 27580 23324 27636 23326
rect 27356 23212 27412 23268
rect 29148 26290 29204 26292
rect 29148 26238 29150 26290
rect 29150 26238 29202 26290
rect 29202 26238 29204 26290
rect 29148 26236 29204 26238
rect 30156 27692 30212 27748
rect 31052 27970 31108 27972
rect 31052 27918 31054 27970
rect 31054 27918 31106 27970
rect 31106 27918 31108 27970
rect 31052 27916 31108 27918
rect 31948 29314 32004 29316
rect 31948 29262 31950 29314
rect 31950 29262 32002 29314
rect 32002 29262 32004 29314
rect 31948 29260 32004 29262
rect 32060 27970 32116 27972
rect 32060 27918 32062 27970
rect 32062 27918 32114 27970
rect 32114 27918 32116 27970
rect 32060 27916 32116 27918
rect 31500 27858 31556 27860
rect 31500 27806 31502 27858
rect 31502 27806 31554 27858
rect 31554 27806 31556 27858
rect 31500 27804 31556 27806
rect 32508 27858 32564 27860
rect 32508 27806 32510 27858
rect 32510 27806 32562 27858
rect 32562 27806 32564 27858
rect 32508 27804 32564 27806
rect 33404 27804 33460 27860
rect 29596 26460 29652 26516
rect 29372 26236 29428 26292
rect 30268 26066 30324 26068
rect 30268 26014 30270 26066
rect 30270 26014 30322 26066
rect 30322 26014 30324 26066
rect 30268 26012 30324 26014
rect 29708 25228 29764 25284
rect 29484 25004 29540 25060
rect 28252 23884 28308 23940
rect 29036 24892 29092 24948
rect 29148 24780 29204 24836
rect 33292 26124 33348 26180
rect 32396 25900 32452 25956
rect 33180 25730 33236 25732
rect 33180 25678 33182 25730
rect 33182 25678 33234 25730
rect 33234 25678 33236 25730
rect 33180 25676 33236 25678
rect 32620 25452 32676 25508
rect 29932 25004 29988 25060
rect 33180 25282 33236 25284
rect 33180 25230 33182 25282
rect 33182 25230 33234 25282
rect 33234 25230 33236 25282
rect 33180 25228 33236 25230
rect 29820 24780 29876 24836
rect 28812 23212 28868 23268
rect 28924 24332 28980 24388
rect 27804 22204 27860 22260
rect 28476 21756 28532 21812
rect 26796 20130 26852 20132
rect 26796 20078 26798 20130
rect 26798 20078 26850 20130
rect 26850 20078 26852 20130
rect 26796 20076 26852 20078
rect 26572 20018 26628 20020
rect 26572 19966 26574 20018
rect 26574 19966 26626 20018
rect 26626 19966 26628 20018
rect 26572 19964 26628 19966
rect 26236 19346 26292 19348
rect 26236 19294 26238 19346
rect 26238 19294 26290 19346
rect 26290 19294 26292 19346
rect 26236 19292 26292 19294
rect 25004 19180 25060 19236
rect 27132 20076 27188 20132
rect 27580 20524 27636 20580
rect 27468 20130 27524 20132
rect 27468 20078 27470 20130
rect 27470 20078 27522 20130
rect 27522 20078 27524 20130
rect 27468 20076 27524 20078
rect 27356 19964 27412 20020
rect 31276 24556 31332 24612
rect 30716 23324 30772 23380
rect 28924 20412 28980 20468
rect 29372 20860 29428 20916
rect 30156 20914 30212 20916
rect 30156 20862 30158 20914
rect 30158 20862 30210 20914
rect 30210 20862 30212 20914
rect 30156 20860 30212 20862
rect 30716 20802 30772 20804
rect 30716 20750 30718 20802
rect 30718 20750 30770 20802
rect 30770 20750 30772 20802
rect 30716 20748 30772 20750
rect 27132 19852 27188 19908
rect 27692 19852 27748 19908
rect 26796 19292 26852 19348
rect 24220 18508 24276 18564
rect 23772 18338 23828 18340
rect 23772 18286 23774 18338
rect 23774 18286 23826 18338
rect 23826 18286 23828 18338
rect 23772 18284 23828 18286
rect 24444 18284 24500 18340
rect 24444 18060 24500 18116
rect 25004 18172 25060 18228
rect 22988 15874 23044 15876
rect 22988 15822 22990 15874
rect 22990 15822 23042 15874
rect 23042 15822 23044 15874
rect 22988 15820 23044 15822
rect 24668 16156 24724 16212
rect 22204 14476 22260 14532
rect 18732 14028 18788 14084
rect 18844 13746 18900 13748
rect 18844 13694 18846 13746
rect 18846 13694 18898 13746
rect 18898 13694 18900 13746
rect 18844 13692 18900 13694
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20748 13970 20804 13972
rect 20748 13918 20750 13970
rect 20750 13918 20802 13970
rect 20802 13918 20804 13970
rect 20748 13916 20804 13918
rect 21308 13916 21364 13972
rect 21084 13804 21140 13860
rect 18732 13580 18788 13636
rect 19516 13468 19572 13524
rect 18732 12908 18788 12964
rect 18284 11452 18340 11508
rect 18508 12460 18564 12516
rect 17836 9996 17892 10052
rect 18396 10722 18452 10724
rect 18396 10670 18398 10722
rect 18398 10670 18450 10722
rect 18450 10670 18452 10722
rect 18396 10668 18452 10670
rect 17948 9772 18004 9828
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 15484 6690 15540 6692
rect 15484 6638 15486 6690
rect 15486 6638 15538 6690
rect 15538 6638 15540 6690
rect 15484 6636 15540 6638
rect 18172 9212 18228 9268
rect 18284 8988 18340 9044
rect 18732 11788 18788 11844
rect 18732 11452 18788 11508
rect 18844 11170 18900 11172
rect 18844 11118 18846 11170
rect 18846 11118 18898 11170
rect 18898 11118 18900 11170
rect 18844 11116 18900 11118
rect 19180 11452 19236 11508
rect 19404 12738 19460 12740
rect 19404 12686 19406 12738
rect 19406 12686 19458 12738
rect 19458 12686 19460 12738
rect 19404 12684 19460 12686
rect 19852 13580 19908 13636
rect 19628 13356 19684 13412
rect 19516 11676 19572 11732
rect 20412 13580 20468 13636
rect 19852 12962 19908 12964
rect 19852 12910 19854 12962
rect 19854 12910 19906 12962
rect 19906 12910 19908 12962
rect 19852 12908 19908 12910
rect 22092 13804 22148 13860
rect 22204 13916 22260 13972
rect 21196 13580 21252 13636
rect 21756 13746 21812 13748
rect 21756 13694 21758 13746
rect 21758 13694 21810 13746
rect 21810 13694 21812 13746
rect 21756 13692 21812 13694
rect 22652 14418 22708 14420
rect 22652 14366 22654 14418
rect 22654 14366 22706 14418
rect 22706 14366 22708 14418
rect 22652 14364 22708 14366
rect 22652 13746 22708 13748
rect 22652 13694 22654 13746
rect 22654 13694 22706 13746
rect 22706 13694 22708 13746
rect 22652 13692 22708 13694
rect 23660 15820 23716 15876
rect 23324 14588 23380 14644
rect 22876 13916 22932 13972
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20188 12572 20244 12628
rect 20044 12516 20100 12518
rect 20860 12572 20916 12628
rect 22540 12850 22596 12852
rect 22540 12798 22542 12850
rect 22542 12798 22594 12850
rect 22594 12798 22596 12850
rect 22540 12796 22596 12798
rect 22428 12348 22484 12404
rect 21196 12066 21252 12068
rect 21196 12014 21198 12066
rect 21198 12014 21250 12066
rect 21250 12014 21252 12066
rect 21196 12012 21252 12014
rect 20188 11788 20244 11844
rect 22652 11564 22708 11620
rect 23212 13468 23268 13524
rect 23324 13746 23380 13748
rect 23324 13694 23326 13746
rect 23326 13694 23378 13746
rect 23378 13694 23380 13746
rect 23324 13692 23380 13694
rect 23548 13580 23604 13636
rect 24332 14252 24388 14308
rect 23772 12962 23828 12964
rect 23772 12910 23774 12962
rect 23774 12910 23826 12962
rect 23826 12910 23828 12962
rect 23772 12908 23828 12910
rect 21308 11452 21364 11508
rect 18844 10332 18900 10388
rect 18732 9826 18788 9828
rect 18732 9774 18734 9826
rect 18734 9774 18786 9826
rect 18786 9774 18788 9826
rect 18732 9772 18788 9774
rect 19180 9772 19236 9828
rect 20300 11004 20356 11060
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 21532 10668 21588 10724
rect 19292 9714 19348 9716
rect 19292 9662 19294 9714
rect 19294 9662 19346 9714
rect 19346 9662 19348 9714
rect 19292 9660 19348 9662
rect 18844 9602 18900 9604
rect 18844 9550 18846 9602
rect 18846 9550 18898 9602
rect 18898 9550 18900 9602
rect 18844 9548 18900 9550
rect 18732 9266 18788 9268
rect 18732 9214 18734 9266
rect 18734 9214 18786 9266
rect 18786 9214 18788 9266
rect 18732 9212 18788 9214
rect 18956 9212 19012 9268
rect 18956 9042 19012 9044
rect 18956 8990 18958 9042
rect 18958 8990 19010 9042
rect 19010 8990 19012 9042
rect 18956 8988 19012 8990
rect 18844 7868 18900 7924
rect 19292 7980 19348 8036
rect 19516 10050 19572 10052
rect 19516 9998 19518 10050
rect 19518 9998 19570 10050
rect 19570 9998 19572 10050
rect 19516 9996 19572 9998
rect 20076 10332 20132 10388
rect 19852 9660 19908 9716
rect 20412 9548 20468 9604
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19628 9212 19684 9268
rect 19404 7868 19460 7924
rect 19516 8988 19572 9044
rect 19068 7532 19124 7588
rect 17500 6636 17556 6692
rect 16156 6578 16212 6580
rect 16156 6526 16158 6578
rect 16158 6526 16210 6578
rect 16210 6526 16212 6578
rect 16156 6524 16212 6526
rect 17388 6524 17444 6580
rect 17500 6076 17556 6132
rect 17724 6748 17780 6804
rect 18620 6802 18676 6804
rect 18620 6750 18622 6802
rect 18622 6750 18674 6802
rect 18674 6750 18676 6802
rect 18620 6748 18676 6750
rect 18956 6578 19012 6580
rect 18956 6526 18958 6578
rect 18958 6526 19010 6578
rect 19010 6526 19012 6578
rect 18956 6524 19012 6526
rect 18396 6076 18452 6132
rect 19404 7474 19460 7476
rect 19404 7422 19406 7474
rect 19406 7422 19458 7474
rect 19458 7422 19460 7474
rect 19404 7420 19460 7422
rect 19292 7196 19348 7252
rect 19180 6466 19236 6468
rect 19180 6414 19182 6466
rect 19182 6414 19234 6466
rect 19234 6414 19236 6466
rect 19180 6412 19236 6414
rect 20300 7980 20356 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19628 7586 19684 7588
rect 19628 7534 19630 7586
rect 19630 7534 19682 7586
rect 19682 7534 19684 7586
rect 19628 7532 19684 7534
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19852 7196 19908 7252
rect 20188 6748 20244 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18396 5180 18452 5236
rect 21420 9602 21476 9604
rect 21420 9550 21422 9602
rect 21422 9550 21474 9602
rect 21474 9550 21476 9602
rect 21420 9548 21476 9550
rect 21644 10332 21700 10388
rect 24556 13468 24612 13524
rect 24108 12796 24164 12852
rect 23324 12402 23380 12404
rect 23324 12350 23326 12402
rect 23326 12350 23378 12402
rect 23378 12350 23380 12402
rect 23324 12348 23380 12350
rect 24780 12684 24836 12740
rect 22764 10332 22820 10388
rect 21756 9884 21812 9940
rect 22204 9938 22260 9940
rect 22204 9886 22206 9938
rect 22206 9886 22258 9938
rect 22258 9886 22260 9938
rect 22204 9884 22260 9886
rect 23436 9714 23492 9716
rect 23436 9662 23438 9714
rect 23438 9662 23490 9714
rect 23490 9662 23492 9714
rect 23436 9660 23492 9662
rect 22428 8428 22484 8484
rect 24556 10610 24612 10612
rect 24556 10558 24558 10610
rect 24558 10558 24610 10610
rect 24610 10558 24612 10610
rect 24556 10556 24612 10558
rect 24668 10108 24724 10164
rect 27132 18396 27188 18452
rect 25340 17388 25396 17444
rect 25228 16210 25284 16212
rect 25228 16158 25230 16210
rect 25230 16158 25282 16210
rect 25282 16158 25284 16210
rect 25228 16156 25284 16158
rect 27580 16994 27636 16996
rect 27580 16942 27582 16994
rect 27582 16942 27634 16994
rect 27634 16942 27636 16994
rect 27580 16940 27636 16942
rect 27916 18284 27972 18340
rect 27916 18060 27972 18116
rect 28252 19964 28308 20020
rect 28476 20076 28532 20132
rect 29148 19852 29204 19908
rect 30492 19964 30548 20020
rect 28476 18956 28532 19012
rect 29932 19010 29988 19012
rect 29932 18958 29934 19010
rect 29934 18958 29986 19010
rect 29986 18958 29988 19010
rect 29932 18956 29988 18958
rect 30156 19010 30212 19012
rect 30156 18958 30158 19010
rect 30158 18958 30210 19010
rect 30210 18958 30212 19010
rect 30156 18956 30212 18958
rect 29372 18620 29428 18676
rect 28588 18450 28644 18452
rect 28588 18398 28590 18450
rect 28590 18398 28642 18450
rect 28642 18398 28644 18450
rect 28588 18396 28644 18398
rect 28140 18338 28196 18340
rect 28140 18286 28142 18338
rect 28142 18286 28194 18338
rect 28194 18286 28196 18338
rect 28140 18284 28196 18286
rect 28700 18284 28756 18340
rect 28028 17388 28084 17444
rect 29148 18284 29204 18340
rect 29148 18060 29204 18116
rect 28700 17164 28756 17220
rect 28924 17612 28980 17668
rect 28364 17052 28420 17108
rect 28140 16994 28196 16996
rect 28140 16942 28142 16994
rect 28142 16942 28194 16994
rect 28194 16942 28196 16994
rect 28140 16940 28196 16942
rect 27468 15986 27524 15988
rect 27468 15934 27470 15986
rect 27470 15934 27522 15986
rect 27522 15934 27524 15986
rect 27468 15932 27524 15934
rect 25788 14588 25844 14644
rect 25228 12738 25284 12740
rect 25228 12686 25230 12738
rect 25230 12686 25282 12738
rect 25282 12686 25284 12738
rect 25228 12684 25284 12686
rect 25340 10610 25396 10612
rect 25340 10558 25342 10610
rect 25342 10558 25394 10610
rect 25394 10558 25396 10610
rect 25340 10556 25396 10558
rect 25004 9884 25060 9940
rect 25340 10332 25396 10388
rect 26460 14642 26516 14644
rect 26460 14590 26462 14642
rect 26462 14590 26514 14642
rect 26514 14590 26516 14642
rect 26460 14588 26516 14590
rect 26796 14418 26852 14420
rect 26796 14366 26798 14418
rect 26798 14366 26850 14418
rect 26850 14366 26852 14418
rect 26796 14364 26852 14366
rect 27580 14642 27636 14644
rect 27580 14590 27582 14642
rect 27582 14590 27634 14642
rect 27634 14590 27636 14642
rect 27580 14588 27636 14590
rect 27132 14306 27188 14308
rect 27132 14254 27134 14306
rect 27134 14254 27186 14306
rect 27186 14254 27188 14306
rect 27132 14252 27188 14254
rect 27020 12684 27076 12740
rect 26236 10834 26292 10836
rect 26236 10782 26238 10834
rect 26238 10782 26290 10834
rect 26290 10782 26292 10834
rect 26236 10780 26292 10782
rect 26572 9772 26628 9828
rect 21532 7420 21588 7476
rect 20748 7250 20804 7252
rect 20748 7198 20750 7250
rect 20750 7198 20802 7250
rect 20802 7198 20804 7250
rect 20748 7196 20804 7198
rect 20524 6972 20580 7028
rect 20636 6636 20692 6692
rect 20412 6412 20468 6468
rect 20300 6300 20356 6356
rect 21308 6972 21364 7028
rect 21420 7196 21476 7252
rect 21308 6636 21364 6692
rect 21196 5852 21252 5908
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22764 6972 22820 7028
rect 22204 6802 22260 6804
rect 22204 6750 22206 6802
rect 22206 6750 22258 6802
rect 22258 6750 22260 6802
rect 22204 6748 22260 6750
rect 23212 6748 23268 6804
rect 21980 6578 22036 6580
rect 21980 6526 21982 6578
rect 21982 6526 22034 6578
rect 22034 6526 22036 6578
rect 21980 6524 22036 6526
rect 21756 6466 21812 6468
rect 21756 6414 21758 6466
rect 21758 6414 21810 6466
rect 21810 6414 21812 6466
rect 21756 6412 21812 6414
rect 22204 6412 22260 6468
rect 21980 5906 22036 5908
rect 21980 5854 21982 5906
rect 21982 5854 22034 5906
rect 22034 5854 22036 5906
rect 21980 5852 22036 5854
rect 21756 5516 21812 5572
rect 21420 5234 21476 5236
rect 21420 5182 21422 5234
rect 21422 5182 21474 5234
rect 21474 5182 21476 5234
rect 21420 5180 21476 5182
rect 23548 6972 23604 7028
rect 23324 6524 23380 6580
rect 23660 6412 23716 6468
rect 24108 7474 24164 7476
rect 24108 7422 24110 7474
rect 24110 7422 24162 7474
rect 24162 7422 24164 7474
rect 24108 7420 24164 7422
rect 23772 7196 23828 7252
rect 23884 6860 23940 6916
rect 24108 6690 24164 6692
rect 24108 6638 24110 6690
rect 24110 6638 24162 6690
rect 24162 6638 24164 6690
rect 24108 6636 24164 6638
rect 23884 6466 23940 6468
rect 23884 6414 23886 6466
rect 23886 6414 23938 6466
rect 23938 6414 23940 6466
rect 23884 6412 23940 6414
rect 25452 8428 25508 8484
rect 24444 6860 24500 6916
rect 24332 6802 24388 6804
rect 24332 6750 24334 6802
rect 24334 6750 24386 6802
rect 24386 6750 24388 6802
rect 24332 6748 24388 6750
rect 24220 6300 24276 6356
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 26572 8428 26628 8484
rect 26348 7980 26404 8036
rect 27132 12348 27188 12404
rect 28252 16716 28308 16772
rect 28812 16770 28868 16772
rect 28812 16718 28814 16770
rect 28814 16718 28866 16770
rect 28866 16718 28868 16770
rect 28812 16716 28868 16718
rect 28140 15986 28196 15988
rect 28140 15934 28142 15986
rect 28142 15934 28194 15986
rect 28194 15934 28196 15986
rect 28140 15932 28196 15934
rect 28364 15986 28420 15988
rect 28364 15934 28366 15986
rect 28366 15934 28418 15986
rect 28418 15934 28420 15986
rect 28364 15932 28420 15934
rect 28476 14700 28532 14756
rect 30716 18956 30772 19012
rect 31836 24610 31892 24612
rect 31836 24558 31838 24610
rect 31838 24558 31890 24610
rect 31890 24558 31892 24610
rect 31836 24556 31892 24558
rect 31276 20524 31332 20580
rect 31612 20130 31668 20132
rect 31612 20078 31614 20130
rect 31614 20078 31666 20130
rect 31666 20078 31668 20130
rect 31612 20076 31668 20078
rect 31052 20018 31108 20020
rect 31052 19966 31054 20018
rect 31054 19966 31106 20018
rect 31106 19966 31108 20018
rect 31052 19964 31108 19966
rect 31388 20018 31444 20020
rect 31388 19966 31390 20018
rect 31390 19966 31442 20018
rect 31442 19966 31444 20018
rect 31388 19964 31444 19966
rect 30604 18620 30660 18676
rect 30492 17666 30548 17668
rect 30492 17614 30494 17666
rect 30494 17614 30546 17666
rect 30546 17614 30548 17666
rect 30492 17612 30548 17614
rect 30828 18060 30884 18116
rect 30828 17724 30884 17780
rect 29708 17052 29764 17108
rect 31500 19068 31556 19124
rect 30940 17052 30996 17108
rect 31052 18956 31108 19012
rect 29372 15986 29428 15988
rect 29372 15934 29374 15986
rect 29374 15934 29426 15986
rect 29426 15934 29428 15986
rect 29372 15932 29428 15934
rect 28924 13916 28980 13972
rect 28476 12572 28532 12628
rect 29372 13804 29428 13860
rect 27580 12348 27636 12404
rect 27244 11340 27300 11396
rect 26684 9548 26740 9604
rect 27020 9772 27076 9828
rect 27468 12012 27524 12068
rect 28364 12402 28420 12404
rect 28364 12350 28366 12402
rect 28366 12350 28418 12402
rect 28418 12350 28420 12402
rect 28364 12348 28420 12350
rect 27916 12066 27972 12068
rect 27916 12014 27918 12066
rect 27918 12014 27970 12066
rect 27970 12014 27972 12066
rect 27916 12012 27972 12014
rect 29484 13020 29540 13076
rect 29484 12348 29540 12404
rect 29372 11452 29428 11508
rect 28252 11394 28308 11396
rect 28252 11342 28254 11394
rect 28254 11342 28306 11394
rect 28306 11342 28308 11394
rect 28252 11340 28308 11342
rect 29260 11394 29316 11396
rect 29260 11342 29262 11394
rect 29262 11342 29314 11394
rect 29314 11342 29316 11394
rect 29260 11340 29316 11342
rect 27580 10668 27636 10724
rect 27356 10108 27412 10164
rect 27692 9660 27748 9716
rect 27580 9602 27636 9604
rect 27580 9550 27582 9602
rect 27582 9550 27634 9602
rect 27634 9550 27636 9602
rect 27580 9548 27636 9550
rect 26908 8258 26964 8260
rect 26908 8206 26910 8258
rect 26910 8206 26962 8258
rect 26962 8206 26964 8258
rect 26908 8204 26964 8206
rect 27356 8258 27412 8260
rect 27356 8206 27358 8258
rect 27358 8206 27410 8258
rect 27410 8206 27412 8258
rect 27356 8204 27412 8206
rect 28028 9826 28084 9828
rect 28028 9774 28030 9826
rect 28030 9774 28082 9826
rect 28082 9774 28084 9826
rect 28028 9772 28084 9774
rect 28588 9714 28644 9716
rect 28588 9662 28590 9714
rect 28590 9662 28642 9714
rect 28642 9662 28644 9714
rect 28588 9660 28644 9662
rect 30044 13916 30100 13972
rect 30156 13692 30212 13748
rect 29932 13020 29988 13076
rect 30492 13634 30548 13636
rect 30492 13582 30494 13634
rect 30494 13582 30546 13634
rect 30546 13582 30548 13634
rect 30492 13580 30548 13582
rect 30380 12796 30436 12852
rect 30156 12460 30212 12516
rect 30380 12348 30436 12404
rect 30156 12178 30212 12180
rect 30156 12126 30158 12178
rect 30158 12126 30210 12178
rect 30210 12126 30212 12178
rect 30156 12124 30212 12126
rect 29708 9884 29764 9940
rect 29932 9714 29988 9716
rect 29932 9662 29934 9714
rect 29934 9662 29986 9714
rect 29986 9662 29988 9714
rect 29932 9660 29988 9662
rect 30044 9602 30100 9604
rect 30044 9550 30046 9602
rect 30046 9550 30098 9602
rect 30098 9550 30100 9602
rect 30044 9548 30100 9550
rect 29708 9436 29764 9492
rect 29820 7980 29876 8036
rect 28028 7756 28084 7812
rect 25788 7250 25844 7252
rect 25788 7198 25790 7250
rect 25790 7198 25842 7250
rect 25842 7198 25844 7250
rect 25788 7196 25844 7198
rect 26796 7196 26852 7252
rect 27244 7474 27300 7476
rect 27244 7422 27246 7474
rect 27246 7422 27298 7474
rect 27298 7422 27300 7474
rect 27244 7420 27300 7422
rect 27020 7308 27076 7364
rect 27692 7362 27748 7364
rect 27692 7310 27694 7362
rect 27694 7310 27746 7362
rect 27746 7310 27748 7362
rect 27692 7308 27748 7310
rect 25228 6578 25284 6580
rect 25228 6526 25230 6578
rect 25230 6526 25282 6578
rect 25282 6526 25284 6578
rect 25228 6524 25284 6526
rect 25116 6188 25172 6244
rect 26236 6690 26292 6692
rect 26236 6638 26238 6690
rect 26238 6638 26290 6690
rect 26290 6638 26292 6690
rect 26236 6636 26292 6638
rect 27244 6636 27300 6692
rect 26572 6578 26628 6580
rect 26572 6526 26574 6578
rect 26574 6526 26626 6578
rect 26626 6526 26628 6578
rect 26572 6524 26628 6526
rect 30492 9938 30548 9940
rect 30492 9886 30494 9938
rect 30494 9886 30546 9938
rect 30546 9886 30548 9938
rect 30492 9884 30548 9886
rect 31388 18060 31444 18116
rect 31500 17164 31556 17220
rect 31724 16716 31780 16772
rect 31724 15202 31780 15204
rect 31724 15150 31726 15202
rect 31726 15150 31778 15202
rect 31778 15150 31780 15202
rect 31724 15148 31780 15150
rect 31500 12796 31556 12852
rect 31612 12348 31668 12404
rect 31948 22764 32004 22820
rect 31948 21644 32004 21700
rect 31948 20188 32004 20244
rect 32060 20130 32116 20132
rect 32060 20078 32062 20130
rect 32062 20078 32114 20130
rect 32114 20078 32116 20130
rect 32060 20076 32116 20078
rect 31948 19068 32004 19124
rect 32172 18396 32228 18452
rect 32284 18284 32340 18340
rect 32508 16770 32564 16772
rect 32508 16718 32510 16770
rect 32510 16718 32562 16770
rect 32562 16718 32564 16770
rect 32508 16716 32564 16718
rect 32060 16098 32116 16100
rect 32060 16046 32062 16098
rect 32062 16046 32114 16098
rect 32114 16046 32116 16098
rect 32060 16044 32116 16046
rect 32508 15820 32564 15876
rect 32396 15148 32452 15204
rect 32620 15708 32676 15764
rect 32060 13634 32116 13636
rect 32060 13582 32062 13634
rect 32062 13582 32114 13634
rect 32114 13582 32116 13634
rect 32060 13580 32116 13582
rect 33180 23324 33236 23380
rect 33180 22482 33236 22484
rect 33180 22430 33182 22482
rect 33182 22430 33234 22482
rect 33234 22430 33236 22482
rect 33180 22428 33236 22430
rect 33068 18732 33124 18788
rect 33740 41858 33796 41860
rect 33740 41806 33742 41858
rect 33742 41806 33794 41858
rect 33794 41806 33796 41858
rect 33740 41804 33796 41806
rect 33628 41298 33684 41300
rect 33628 41246 33630 41298
rect 33630 41246 33682 41298
rect 33682 41246 33684 41298
rect 33628 41244 33684 41246
rect 34076 42140 34132 42196
rect 33964 41692 34020 41748
rect 34076 41356 34132 41412
rect 33628 36988 33684 37044
rect 34524 41132 34580 41188
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35532 42082 35588 42084
rect 35532 42030 35534 42082
rect 35534 42030 35586 42082
rect 35586 42030 35588 42082
rect 35532 42028 35588 42030
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 36428 43260 36484 43316
rect 34076 38444 34132 38500
rect 33964 37884 34020 37940
rect 33852 34860 33908 34916
rect 33964 37548 34020 37604
rect 34300 37212 34356 37268
rect 34076 37154 34132 37156
rect 34076 37102 34078 37154
rect 34078 37102 34130 37154
rect 34130 37102 34132 37154
rect 34076 37100 34132 37102
rect 35084 40962 35140 40964
rect 35084 40910 35086 40962
rect 35086 40910 35138 40962
rect 35138 40910 35140 40962
rect 35084 40908 35140 40910
rect 34972 40460 35028 40516
rect 34636 37324 34692 37380
rect 34748 38668 34804 38724
rect 34412 36988 34468 37044
rect 34188 35586 34244 35588
rect 34188 35534 34190 35586
rect 34190 35534 34242 35586
rect 34242 35534 34244 35586
rect 34188 35532 34244 35534
rect 35644 40908 35700 40964
rect 35644 40514 35700 40516
rect 35644 40462 35646 40514
rect 35646 40462 35698 40514
rect 35698 40462 35700 40514
rect 35644 40460 35700 40462
rect 37548 45388 37604 45444
rect 37660 46620 37716 46676
rect 39900 46786 39956 46788
rect 39900 46734 39902 46786
rect 39902 46734 39954 46786
rect 39954 46734 39956 46786
rect 39900 46732 39956 46734
rect 38892 46674 38948 46676
rect 38892 46622 38894 46674
rect 38894 46622 38946 46674
rect 38946 46622 38948 46674
rect 38892 46620 38948 46622
rect 39564 46396 39620 46452
rect 37996 45612 38052 45668
rect 38332 45388 38388 45444
rect 37772 42924 37828 42980
rect 38108 43260 38164 43316
rect 36876 41804 36932 41860
rect 36652 41356 36708 41412
rect 36092 41186 36148 41188
rect 36092 41134 36094 41186
rect 36094 41134 36146 41186
rect 36146 41134 36148 41186
rect 36092 41132 36148 41134
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 39730 35252 39732
rect 35196 39678 35198 39730
rect 35198 39678 35250 39730
rect 35250 39678 35252 39730
rect 35196 39676 35252 39678
rect 37436 41186 37492 41188
rect 37436 41134 37438 41186
rect 37438 41134 37490 41186
rect 37490 41134 37492 41186
rect 37436 41132 37492 41134
rect 37100 39676 37156 39732
rect 38220 41916 38276 41972
rect 38108 41858 38164 41860
rect 38108 41806 38110 41858
rect 38110 41806 38162 41858
rect 38162 41806 38164 41858
rect 38108 41804 38164 41806
rect 37548 38946 37604 38948
rect 37548 38894 37550 38946
rect 37550 38894 37602 38946
rect 37602 38894 37604 38946
rect 37548 38892 37604 38894
rect 37100 38668 37156 38724
rect 35532 38556 35588 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 36316 38162 36372 38164
rect 36316 38110 36318 38162
rect 36318 38110 36370 38162
rect 36370 38110 36372 38162
rect 36316 38108 36372 38110
rect 37324 38108 37380 38164
rect 35308 38050 35364 38052
rect 35308 37998 35310 38050
rect 35310 37998 35362 38050
rect 35362 37998 35364 38050
rect 35308 37996 35364 37998
rect 35532 37548 35588 37604
rect 35756 37378 35812 37380
rect 35756 37326 35758 37378
rect 35758 37326 35810 37378
rect 35810 37326 35812 37378
rect 35756 37324 35812 37326
rect 35644 37212 35700 37268
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35756 36876 35812 36932
rect 35196 36540 35252 36596
rect 35420 36482 35476 36484
rect 35420 36430 35422 36482
rect 35422 36430 35474 36482
rect 35474 36430 35476 36482
rect 35420 36428 35476 36430
rect 35196 35756 35252 35812
rect 35532 35644 35588 35700
rect 34972 35532 35028 35588
rect 34972 35308 35028 35364
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34748 34972 34804 35028
rect 34972 34860 35028 34916
rect 33628 34076 33684 34132
rect 34524 33180 34580 33236
rect 34748 32732 34804 32788
rect 34860 33516 34916 33572
rect 33852 31836 33908 31892
rect 33740 30156 33796 30212
rect 34636 32060 34692 32116
rect 34524 31778 34580 31780
rect 34524 31726 34526 31778
rect 34526 31726 34578 31778
rect 34578 31726 34580 31778
rect 34524 31724 34580 31726
rect 34524 31500 34580 31556
rect 34860 32284 34916 32340
rect 34748 29650 34804 29652
rect 34748 29598 34750 29650
rect 34750 29598 34802 29650
rect 34802 29598 34804 29650
rect 34748 29596 34804 29598
rect 34524 27858 34580 27860
rect 34524 27806 34526 27858
rect 34526 27806 34578 27858
rect 34578 27806 34580 27858
rect 34524 27804 34580 27806
rect 35084 34748 35140 34804
rect 35084 33852 35140 33908
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 32732 35140 32788
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 31836 35252 31892
rect 35420 31778 35476 31780
rect 35420 31726 35422 31778
rect 35422 31726 35474 31778
rect 35474 31726 35476 31778
rect 35420 31724 35476 31726
rect 35196 31612 35252 31668
rect 35084 31500 35140 31556
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35756 35026 35812 35028
rect 35756 34974 35758 35026
rect 35758 34974 35810 35026
rect 35810 34974 35812 35026
rect 35756 34972 35812 34974
rect 35980 37938 36036 37940
rect 35980 37886 35982 37938
rect 35982 37886 36034 37938
rect 36034 37886 36036 37938
rect 35980 37884 36036 37886
rect 36204 37826 36260 37828
rect 36204 37774 36206 37826
rect 36206 37774 36258 37826
rect 36258 37774 36260 37826
rect 36204 37772 36260 37774
rect 36204 37212 36260 37268
rect 36092 36988 36148 37044
rect 35980 35698 36036 35700
rect 35980 35646 35982 35698
rect 35982 35646 36034 35698
rect 36034 35646 36036 35698
rect 35980 35644 36036 35646
rect 36204 36764 36260 36820
rect 36988 37996 37044 38052
rect 36652 37266 36708 37268
rect 36652 37214 36654 37266
rect 36654 37214 36706 37266
rect 36706 37214 36708 37266
rect 36652 37212 36708 37214
rect 36540 35868 36596 35924
rect 36316 35810 36372 35812
rect 36316 35758 36318 35810
rect 36318 35758 36370 35810
rect 36370 35758 36372 35810
rect 36316 35756 36372 35758
rect 36428 35532 36484 35588
rect 36652 35420 36708 35476
rect 36204 35308 36260 35364
rect 36204 34914 36260 34916
rect 36204 34862 36206 34914
rect 36206 34862 36258 34914
rect 36258 34862 36260 34914
rect 36204 34860 36260 34862
rect 36092 34130 36148 34132
rect 36092 34078 36094 34130
rect 36094 34078 36146 34130
rect 36146 34078 36148 34130
rect 36092 34076 36148 34078
rect 36092 33906 36148 33908
rect 36092 33854 36094 33906
rect 36094 33854 36146 33906
rect 36146 33854 36148 33906
rect 36092 33852 36148 33854
rect 36876 36706 36932 36708
rect 36876 36654 36878 36706
rect 36878 36654 36930 36706
rect 36930 36654 36932 36706
rect 36876 36652 36932 36654
rect 37100 37490 37156 37492
rect 37100 37438 37102 37490
rect 37102 37438 37154 37490
rect 37154 37438 37156 37490
rect 37100 37436 37156 37438
rect 37100 36764 37156 36820
rect 37212 36428 37268 36484
rect 36652 33964 36708 34020
rect 36988 35308 37044 35364
rect 37996 38892 38052 38948
rect 38108 39564 38164 39620
rect 37884 38108 37940 38164
rect 38892 45276 38948 45332
rect 44268 54012 44324 54068
rect 43148 53900 43204 53956
rect 44268 53676 44324 53732
rect 47964 56252 48020 56308
rect 46732 55356 46788 55412
rect 46060 54572 46116 54628
rect 46844 54572 46900 54628
rect 46956 55132 47012 55188
rect 45500 53564 45556 53620
rect 45836 53676 45892 53732
rect 43820 52780 43876 52836
rect 45500 52220 45556 52276
rect 43148 52050 43204 52052
rect 43148 51998 43150 52050
rect 43150 51998 43202 52050
rect 43202 51998 43204 52050
rect 43148 51996 43204 51998
rect 44156 52050 44212 52052
rect 44156 51998 44158 52050
rect 44158 51998 44210 52050
rect 44210 51998 44212 52050
rect 44156 51996 44212 51998
rect 42476 51548 42532 51604
rect 43260 51602 43316 51604
rect 43260 51550 43262 51602
rect 43262 51550 43314 51602
rect 43314 51550 43316 51602
rect 43260 51548 43316 51550
rect 41020 50764 41076 50820
rect 43260 51324 43316 51380
rect 41804 51212 41860 51268
rect 42252 51266 42308 51268
rect 42252 51214 42254 51266
rect 42254 51214 42306 51266
rect 42306 51214 42308 51266
rect 42252 51212 42308 51214
rect 41804 50818 41860 50820
rect 41804 50766 41806 50818
rect 41806 50766 41858 50818
rect 41858 50766 41860 50818
rect 41804 50764 41860 50766
rect 41468 50594 41524 50596
rect 41468 50542 41470 50594
rect 41470 50542 41522 50594
rect 41522 50542 41524 50594
rect 41468 50540 41524 50542
rect 41020 50034 41076 50036
rect 41020 49982 41022 50034
rect 41022 49982 41074 50034
rect 41074 49982 41076 50034
rect 41020 49980 41076 49982
rect 41468 49810 41524 49812
rect 41468 49758 41470 49810
rect 41470 49758 41522 49810
rect 41522 49758 41524 49810
rect 41468 49756 41524 49758
rect 42140 49980 42196 50036
rect 42812 50594 42868 50596
rect 42812 50542 42814 50594
rect 42814 50542 42866 50594
rect 42866 50542 42868 50594
rect 42812 50540 42868 50542
rect 42252 49756 42308 49812
rect 42140 49698 42196 49700
rect 42140 49646 42142 49698
rect 42142 49646 42194 49698
rect 42194 49646 42196 49698
rect 42140 49644 42196 49646
rect 41580 48130 41636 48132
rect 41580 48078 41582 48130
rect 41582 48078 41634 48130
rect 41634 48078 41636 48130
rect 41580 48076 41636 48078
rect 40908 46450 40964 46452
rect 40908 46398 40910 46450
rect 40910 46398 40962 46450
rect 40962 46398 40964 46450
rect 40908 46396 40964 46398
rect 41692 47516 41748 47572
rect 42364 48354 42420 48356
rect 42364 48302 42366 48354
rect 42366 48302 42418 48354
rect 42418 48302 42420 48354
rect 42364 48300 42420 48302
rect 42588 48076 42644 48132
rect 42140 47516 42196 47572
rect 40684 45276 40740 45332
rect 40236 44828 40292 44884
rect 38892 44268 38948 44324
rect 39116 44380 39172 44436
rect 38444 41916 38500 41972
rect 39004 42924 39060 42980
rect 38892 41916 38948 41972
rect 40796 44322 40852 44324
rect 40796 44270 40798 44322
rect 40798 44270 40850 44322
rect 40850 44270 40852 44322
rect 40796 44268 40852 44270
rect 42700 47852 42756 47908
rect 41916 45276 41972 45332
rect 41020 43538 41076 43540
rect 41020 43486 41022 43538
rect 41022 43486 41074 43538
rect 41074 43486 41076 43538
rect 41020 43484 41076 43486
rect 40348 43426 40404 43428
rect 40348 43374 40350 43426
rect 40350 43374 40402 43426
rect 40402 43374 40404 43426
rect 40348 43372 40404 43374
rect 40796 42924 40852 42980
rect 41468 43538 41524 43540
rect 41468 43486 41470 43538
rect 41470 43486 41522 43538
rect 41522 43486 41524 43538
rect 41468 43484 41524 43486
rect 39788 42588 39844 42644
rect 40572 42642 40628 42644
rect 40572 42590 40574 42642
rect 40574 42590 40626 42642
rect 40626 42590 40628 42642
rect 40572 42588 40628 42590
rect 41692 42642 41748 42644
rect 41692 42590 41694 42642
rect 41694 42590 41746 42642
rect 41746 42590 41748 42642
rect 41692 42588 41748 42590
rect 39340 42028 39396 42084
rect 39452 42364 39508 42420
rect 37548 36652 37604 36708
rect 37772 37548 37828 37604
rect 38332 36428 38388 36484
rect 37324 35922 37380 35924
rect 37324 35870 37326 35922
rect 37326 35870 37378 35922
rect 37378 35870 37380 35922
rect 37324 35868 37380 35870
rect 37436 35644 37492 35700
rect 37212 34690 37268 34692
rect 37212 34638 37214 34690
rect 37214 34638 37266 34690
rect 37266 34638 37268 34690
rect 37212 34636 37268 34638
rect 38332 35922 38388 35924
rect 38332 35870 38334 35922
rect 38334 35870 38386 35922
rect 38386 35870 38388 35922
rect 38332 35868 38388 35870
rect 37100 34130 37156 34132
rect 37100 34078 37102 34130
rect 37102 34078 37154 34130
rect 37154 34078 37156 34130
rect 37100 34076 37156 34078
rect 37996 35698 38052 35700
rect 37996 35646 37998 35698
rect 37998 35646 38050 35698
rect 38050 35646 38052 35698
rect 37996 35644 38052 35646
rect 37884 34860 37940 34916
rect 37660 34636 37716 34692
rect 37660 34018 37716 34020
rect 37660 33966 37662 34018
rect 37662 33966 37714 34018
rect 37714 33966 37716 34018
rect 37660 33964 37716 33966
rect 37548 33570 37604 33572
rect 37548 33518 37550 33570
rect 37550 33518 37602 33570
rect 37602 33518 37604 33570
rect 37548 33516 37604 33518
rect 37212 32562 37268 32564
rect 37212 32510 37214 32562
rect 37214 32510 37266 32562
rect 37266 32510 37268 32562
rect 37212 32508 37268 32510
rect 37100 32396 37156 32452
rect 37660 32450 37716 32452
rect 37660 32398 37662 32450
rect 37662 32398 37714 32450
rect 37714 32398 37716 32450
rect 37660 32396 37716 32398
rect 37212 32284 37268 32340
rect 38108 35532 38164 35588
rect 38220 35420 38276 35476
rect 38780 38162 38836 38164
rect 38780 38110 38782 38162
rect 38782 38110 38834 38162
rect 38834 38110 38836 38162
rect 38780 38108 38836 38110
rect 38668 37884 38724 37940
rect 38780 37324 38836 37380
rect 39228 37100 39284 37156
rect 39004 35922 39060 35924
rect 39004 35870 39006 35922
rect 39006 35870 39058 35922
rect 39058 35870 39060 35922
rect 39004 35868 39060 35870
rect 39116 35698 39172 35700
rect 39116 35646 39118 35698
rect 39118 35646 39170 35698
rect 39170 35646 39172 35698
rect 39116 35644 39172 35646
rect 38108 33516 38164 33572
rect 38556 35532 38612 35588
rect 38780 34972 38836 35028
rect 38668 34690 38724 34692
rect 38668 34638 38670 34690
rect 38670 34638 38722 34690
rect 38722 34638 38724 34690
rect 38668 34636 38724 34638
rect 40348 41692 40404 41748
rect 40348 41132 40404 41188
rect 41132 41020 41188 41076
rect 40236 40348 40292 40404
rect 41244 40402 41300 40404
rect 41244 40350 41246 40402
rect 41246 40350 41298 40402
rect 41298 40350 41300 40402
rect 41244 40348 41300 40350
rect 41468 40348 41524 40404
rect 41692 41692 41748 41748
rect 41692 40348 41748 40404
rect 39788 39452 39844 39508
rect 39676 38556 39732 38612
rect 39564 37378 39620 37380
rect 39564 37326 39566 37378
rect 39566 37326 39618 37378
rect 39618 37326 39620 37378
rect 39564 37324 39620 37326
rect 39676 37100 39732 37156
rect 39340 34972 39396 35028
rect 39116 34748 39172 34804
rect 37996 32562 38052 32564
rect 37996 32510 37998 32562
rect 37998 32510 38050 32562
rect 38050 32510 38052 32562
rect 37996 32508 38052 32510
rect 36988 31948 37044 32004
rect 36204 31500 36260 31556
rect 37772 31836 37828 31892
rect 37436 31778 37492 31780
rect 37436 31726 37438 31778
rect 37438 31726 37490 31778
rect 37490 31726 37492 31778
rect 37436 31724 37492 31726
rect 37884 31778 37940 31780
rect 37884 31726 37886 31778
rect 37886 31726 37938 31778
rect 37938 31726 37940 31778
rect 37884 31724 37940 31726
rect 37100 31500 37156 31556
rect 35084 30156 35140 30212
rect 37100 30210 37156 30212
rect 37100 30158 37102 30210
rect 37102 30158 37154 30210
rect 37154 30158 37156 30210
rect 37100 30156 37156 30158
rect 34972 28028 35028 28084
rect 35084 29148 35140 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 28588 35140 28644
rect 35308 28812 35364 28868
rect 37772 29820 37828 29876
rect 36876 29426 36932 29428
rect 36876 29374 36878 29426
rect 36878 29374 36930 29426
rect 36930 29374 36932 29426
rect 36876 29372 36932 29374
rect 36540 29260 36596 29316
rect 35980 28812 36036 28868
rect 34860 27580 34916 27636
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 36092 28588 36148 28644
rect 35420 26572 35476 26628
rect 34412 26514 34468 26516
rect 34412 26462 34414 26514
rect 34414 26462 34466 26514
rect 34466 26462 34468 26514
rect 34412 26460 34468 26462
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34188 25618 34244 25620
rect 34188 25566 34190 25618
rect 34190 25566 34242 25618
rect 34242 25566 34244 25618
rect 34188 25564 34244 25566
rect 33516 25004 33572 25060
rect 33740 25452 33796 25508
rect 33740 25228 33796 25284
rect 34076 25282 34132 25284
rect 34076 25230 34078 25282
rect 34078 25230 34130 25282
rect 34130 25230 34132 25282
rect 34076 25228 34132 25230
rect 34188 24780 34244 24836
rect 33628 23154 33684 23156
rect 33628 23102 33630 23154
rect 33630 23102 33682 23154
rect 33682 23102 33684 23154
rect 33628 23100 33684 23102
rect 34972 25564 35028 25620
rect 34636 25452 34692 25508
rect 35308 25340 35364 25396
rect 36204 25618 36260 25620
rect 36204 25566 36206 25618
rect 36206 25566 36258 25618
rect 36258 25566 36260 25618
rect 36204 25564 36260 25566
rect 35420 24722 35476 24724
rect 35420 24670 35422 24722
rect 35422 24670 35474 24722
rect 35474 24670 35476 24722
rect 35420 24668 35476 24670
rect 35308 24556 35364 24612
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36764 25340 36820 25396
rect 36092 25228 36148 25284
rect 36540 25116 36596 25172
rect 35980 24556 36036 24612
rect 34076 23154 34132 23156
rect 34076 23102 34078 23154
rect 34078 23102 34130 23154
rect 34130 23102 34132 23154
rect 34076 23100 34132 23102
rect 33516 22764 33572 22820
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35532 22540 35588 22596
rect 33516 22428 33572 22484
rect 33404 22092 33460 22148
rect 33180 17106 33236 17108
rect 33180 17054 33182 17106
rect 33182 17054 33234 17106
rect 33234 17054 33236 17106
rect 33180 17052 33236 17054
rect 33068 15708 33124 15764
rect 32620 14588 32676 14644
rect 32172 13020 32228 13076
rect 33068 13746 33124 13748
rect 33068 13694 33070 13746
rect 33070 13694 33122 13746
rect 33122 13694 33124 13746
rect 33068 13692 33124 13694
rect 32396 12796 32452 12852
rect 32508 12348 32564 12404
rect 31164 10722 31220 10724
rect 31164 10670 31166 10722
rect 31166 10670 31218 10722
rect 31218 10670 31220 10722
rect 31164 10668 31220 10670
rect 31836 11506 31892 11508
rect 31836 11454 31838 11506
rect 31838 11454 31890 11506
rect 31890 11454 31892 11506
rect 31836 11452 31892 11454
rect 31836 11116 31892 11172
rect 31724 10722 31780 10724
rect 31724 10670 31726 10722
rect 31726 10670 31778 10722
rect 31778 10670 31780 10722
rect 31724 10668 31780 10670
rect 31052 9996 31108 10052
rect 31164 9884 31220 9940
rect 31388 9772 31444 9828
rect 30604 9602 30660 9604
rect 30604 9550 30606 9602
rect 30606 9550 30658 9602
rect 30658 9550 30660 9602
rect 30604 9548 30660 9550
rect 33628 21810 33684 21812
rect 33628 21758 33630 21810
rect 33630 21758 33682 21810
rect 33682 21758 33684 21810
rect 33628 21756 33684 21758
rect 36428 22540 36484 22596
rect 36316 21756 36372 21812
rect 34524 21644 34580 21700
rect 33964 20802 34020 20804
rect 33964 20750 33966 20802
rect 33966 20750 34018 20802
rect 34018 20750 34020 20802
rect 33964 20748 34020 20750
rect 33740 20412 33796 20468
rect 34860 21586 34916 21588
rect 34860 21534 34862 21586
rect 34862 21534 34914 21586
rect 34914 21534 34916 21586
rect 34860 21532 34916 21534
rect 34300 19404 34356 19460
rect 34188 19346 34244 19348
rect 34188 19294 34190 19346
rect 34190 19294 34242 19346
rect 34242 19294 34244 19346
rect 34188 19292 34244 19294
rect 34636 19292 34692 19348
rect 34076 19180 34132 19236
rect 33852 18674 33908 18676
rect 33852 18622 33854 18674
rect 33854 18622 33906 18674
rect 33906 18622 33908 18674
rect 33852 18620 33908 18622
rect 33516 18396 33572 18452
rect 33628 18508 33684 18564
rect 33628 16098 33684 16100
rect 33628 16046 33630 16098
rect 33630 16046 33682 16098
rect 33682 16046 33684 16098
rect 33628 16044 33684 16046
rect 34972 19010 35028 19012
rect 34972 18958 34974 19010
rect 34974 18958 35026 19010
rect 35026 18958 35028 19010
rect 34972 18956 35028 18958
rect 35644 21586 35700 21588
rect 35644 21534 35646 21586
rect 35646 21534 35698 21586
rect 35698 21534 35700 21586
rect 35644 21532 35700 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35420 19234 35476 19236
rect 35420 19182 35422 19234
rect 35422 19182 35474 19234
rect 35474 19182 35476 19234
rect 35420 19180 35476 19182
rect 35084 18620 35140 18676
rect 34636 18508 34692 18564
rect 35980 18508 36036 18564
rect 35308 18284 35364 18340
rect 35532 18396 35588 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34300 15986 34356 15988
rect 34300 15934 34302 15986
rect 34302 15934 34354 15986
rect 34354 15934 34356 15986
rect 34300 15932 34356 15934
rect 33852 15820 33908 15876
rect 33740 15148 33796 15204
rect 32060 11618 32116 11620
rect 32060 11566 32062 11618
rect 32062 11566 32114 11618
rect 32114 11566 32116 11618
rect 32060 11564 32116 11566
rect 33068 13074 33124 13076
rect 33068 13022 33070 13074
rect 33070 13022 33122 13074
rect 33122 13022 33124 13074
rect 33068 13020 33124 13022
rect 33404 13020 33460 13076
rect 33292 12796 33348 12852
rect 32284 9938 32340 9940
rect 32284 9886 32286 9938
rect 32286 9886 32338 9938
rect 32338 9886 32340 9938
rect 32284 9884 32340 9886
rect 31836 9826 31892 9828
rect 31836 9774 31838 9826
rect 31838 9774 31890 9826
rect 31890 9774 31892 9826
rect 31836 9772 31892 9774
rect 28140 7420 28196 7476
rect 26012 6300 26068 6356
rect 30268 6524 30324 6580
rect 30492 6636 30548 6692
rect 28140 6188 28196 6244
rect 27580 6076 27636 6132
rect 25340 4338 25396 4340
rect 25340 4286 25342 4338
rect 25342 4286 25394 4338
rect 25394 4286 25396 4338
rect 25340 4284 25396 4286
rect 29372 5404 29428 5460
rect 28588 4562 28644 4564
rect 28588 4510 28590 4562
rect 28590 4510 28642 4562
rect 28642 4510 28644 4562
rect 28588 4508 28644 4510
rect 29708 5180 29764 5236
rect 30940 8316 30996 8372
rect 30716 8034 30772 8036
rect 30716 7982 30718 8034
rect 30718 7982 30770 8034
rect 30770 7982 30772 8034
rect 30716 7980 30772 7982
rect 33404 12684 33460 12740
rect 33404 12124 33460 12180
rect 33740 13692 33796 13748
rect 34076 14140 34132 14196
rect 35084 17388 35140 17444
rect 35532 16940 35588 16996
rect 36316 18732 36372 18788
rect 35980 17442 36036 17444
rect 35980 17390 35982 17442
rect 35982 17390 36034 17442
rect 36034 17390 36036 17442
rect 35980 17388 36036 17390
rect 36764 21810 36820 21812
rect 36764 21758 36766 21810
rect 36766 21758 36818 21810
rect 36818 21758 36820 21810
rect 36764 21756 36820 21758
rect 37324 28642 37380 28644
rect 37324 28590 37326 28642
rect 37326 28590 37378 28642
rect 37378 28590 37380 28642
rect 37324 28588 37380 28590
rect 37324 28364 37380 28420
rect 37100 27244 37156 27300
rect 36988 26908 37044 26964
rect 37100 26460 37156 26516
rect 37100 25282 37156 25284
rect 37100 25230 37102 25282
rect 37102 25230 37154 25282
rect 37154 25230 37156 25282
rect 37100 25228 37156 25230
rect 37884 29372 37940 29428
rect 37436 28140 37492 28196
rect 37772 27580 37828 27636
rect 38220 31836 38276 31892
rect 38108 28364 38164 28420
rect 37660 26572 37716 26628
rect 37324 25676 37380 25732
rect 37324 25394 37380 25396
rect 37324 25342 37326 25394
rect 37326 25342 37378 25394
rect 37378 25342 37380 25394
rect 37324 25340 37380 25342
rect 38108 28140 38164 28196
rect 38108 27692 38164 27748
rect 38220 27244 38276 27300
rect 38108 26908 38164 26964
rect 37996 26460 38052 26516
rect 38892 33346 38948 33348
rect 38892 33294 38894 33346
rect 38894 33294 38946 33346
rect 38946 33294 38948 33346
rect 38892 33292 38948 33294
rect 39340 34690 39396 34692
rect 39340 34638 39342 34690
rect 39342 34638 39394 34690
rect 39394 34638 39396 34690
rect 39340 34636 39396 34638
rect 39228 34130 39284 34132
rect 39228 34078 39230 34130
rect 39230 34078 39282 34130
rect 39282 34078 39284 34130
rect 39228 34076 39284 34078
rect 39676 34130 39732 34132
rect 39676 34078 39678 34130
rect 39678 34078 39730 34130
rect 39730 34078 39732 34130
rect 39676 34076 39732 34078
rect 41692 39452 41748 39508
rect 40236 38556 40292 38612
rect 40908 37154 40964 37156
rect 40908 37102 40910 37154
rect 40910 37102 40962 37154
rect 40962 37102 40964 37154
rect 40908 37100 40964 37102
rect 41244 37100 41300 37156
rect 41804 37212 41860 37268
rect 40124 35196 40180 35252
rect 40796 35026 40852 35028
rect 40796 34974 40798 35026
rect 40798 34974 40850 35026
rect 40850 34974 40852 35026
rect 40796 34972 40852 34974
rect 40124 34188 40180 34244
rect 40236 34412 40292 34468
rect 38444 31724 38500 31780
rect 39564 32284 39620 32340
rect 38668 29932 38724 29988
rect 39116 29148 39172 29204
rect 38780 28028 38836 28084
rect 38444 27970 38500 27972
rect 38444 27918 38446 27970
rect 38446 27918 38498 27970
rect 38498 27918 38500 27970
rect 38444 27916 38500 27918
rect 38668 27692 38724 27748
rect 38668 27244 38724 27300
rect 39004 27970 39060 27972
rect 39004 27918 39006 27970
rect 39006 27918 39058 27970
rect 39058 27918 39060 27970
rect 39004 27916 39060 27918
rect 39116 27580 39172 27636
rect 38892 27132 38948 27188
rect 38444 26460 38500 26516
rect 37548 25394 37604 25396
rect 37548 25342 37550 25394
rect 37550 25342 37602 25394
rect 37602 25342 37604 25394
rect 37548 25340 37604 25342
rect 37436 25228 37492 25284
rect 37996 25282 38052 25284
rect 37996 25230 37998 25282
rect 37998 25230 38050 25282
rect 38050 25230 38052 25282
rect 37996 25228 38052 25230
rect 38332 25394 38388 25396
rect 38332 25342 38334 25394
rect 38334 25342 38386 25394
rect 38386 25342 38388 25394
rect 38332 25340 38388 25342
rect 38444 24668 38500 24724
rect 39228 26514 39284 26516
rect 39228 26462 39230 26514
rect 39230 26462 39282 26514
rect 39282 26462 39284 26514
rect 39228 26460 39284 26462
rect 39452 26460 39508 26516
rect 39116 26066 39172 26068
rect 39116 26014 39118 26066
rect 39118 26014 39170 26066
rect 39170 26014 39172 26066
rect 39116 26012 39172 26014
rect 39452 26290 39508 26292
rect 39452 26238 39454 26290
rect 39454 26238 39506 26290
rect 39506 26238 39508 26290
rect 39452 26236 39508 26238
rect 39228 25394 39284 25396
rect 39228 25342 39230 25394
rect 39230 25342 39282 25394
rect 39282 25342 39284 25394
rect 39228 25340 39284 25342
rect 41244 34972 41300 35028
rect 40460 34076 40516 34132
rect 40460 32674 40516 32676
rect 40460 32622 40462 32674
rect 40462 32622 40514 32674
rect 40514 32622 40516 32674
rect 40460 32620 40516 32622
rect 40348 29986 40404 29988
rect 40348 29934 40350 29986
rect 40350 29934 40402 29986
rect 40402 29934 40404 29986
rect 40348 29932 40404 29934
rect 39788 29820 39844 29876
rect 40236 29314 40292 29316
rect 40236 29262 40238 29314
rect 40238 29262 40290 29314
rect 40290 29262 40292 29314
rect 40236 29260 40292 29262
rect 40124 29202 40180 29204
rect 40124 29150 40126 29202
rect 40126 29150 40178 29202
rect 40178 29150 40180 29202
rect 40124 29148 40180 29150
rect 40012 27186 40068 27188
rect 40012 27134 40014 27186
rect 40014 27134 40066 27186
rect 40066 27134 40068 27186
rect 40012 27132 40068 27134
rect 41468 34354 41524 34356
rect 41468 34302 41470 34354
rect 41470 34302 41522 34354
rect 41522 34302 41524 34354
rect 41468 34300 41524 34302
rect 41244 34076 41300 34132
rect 41804 33180 41860 33236
rect 40908 32562 40964 32564
rect 40908 32510 40910 32562
rect 40910 32510 40962 32562
rect 40962 32510 40964 32562
rect 40908 32508 40964 32510
rect 41468 31836 41524 31892
rect 41804 32674 41860 32676
rect 41804 32622 41806 32674
rect 41806 32622 41858 32674
rect 41858 32622 41860 32674
rect 41804 32620 41860 32622
rect 42140 44268 42196 44324
rect 42252 43372 42308 43428
rect 42476 43426 42532 43428
rect 42476 43374 42478 43426
rect 42478 43374 42530 43426
rect 42530 43374 42532 43426
rect 42476 43372 42532 43374
rect 42252 42924 42308 42980
rect 42028 42642 42084 42644
rect 42028 42590 42030 42642
rect 42030 42590 42082 42642
rect 42082 42590 42084 42642
rect 42028 42588 42084 42590
rect 42252 41074 42308 41076
rect 42252 41022 42254 41074
rect 42254 41022 42306 41074
rect 42306 41022 42308 41074
rect 42252 41020 42308 41022
rect 42588 41020 42644 41076
rect 42140 40348 42196 40404
rect 42252 39228 42308 39284
rect 42476 35698 42532 35700
rect 42476 35646 42478 35698
rect 42478 35646 42530 35698
rect 42530 35646 42532 35698
rect 42476 35644 42532 35646
rect 42364 34860 42420 34916
rect 42364 34354 42420 34356
rect 42364 34302 42366 34354
rect 42366 34302 42418 34354
rect 42418 34302 42420 34354
rect 42364 34300 42420 34302
rect 42028 34130 42084 34132
rect 42028 34078 42030 34130
rect 42030 34078 42082 34130
rect 42082 34078 42084 34130
rect 42028 34076 42084 34078
rect 42364 33180 42420 33236
rect 41916 32508 41972 32564
rect 42028 32284 42084 32340
rect 42252 32508 42308 32564
rect 42252 32284 42308 32340
rect 43708 51548 43764 51604
rect 45276 51212 45332 51268
rect 44156 50540 44212 50596
rect 44828 50594 44884 50596
rect 44828 50542 44830 50594
rect 44830 50542 44882 50594
rect 44882 50542 44884 50594
rect 44828 50540 44884 50542
rect 43372 49644 43428 49700
rect 43036 48188 43092 48244
rect 43372 48354 43428 48356
rect 43372 48302 43374 48354
rect 43374 48302 43426 48354
rect 43426 48302 43428 48354
rect 43372 48300 43428 48302
rect 42924 47516 42980 47572
rect 43484 48242 43540 48244
rect 43484 48190 43486 48242
rect 43486 48190 43538 48242
rect 43538 48190 43540 48242
rect 43484 48188 43540 48190
rect 43484 47180 43540 47236
rect 43596 47516 43652 47572
rect 43260 46732 43316 46788
rect 44268 47570 44324 47572
rect 44268 47518 44270 47570
rect 44270 47518 44322 47570
rect 44322 47518 44324 47570
rect 44268 47516 44324 47518
rect 44828 47516 44884 47572
rect 43932 46956 43988 47012
rect 44828 47180 44884 47236
rect 44492 46674 44548 46676
rect 44492 46622 44494 46674
rect 44494 46622 44546 46674
rect 44546 46622 44548 46674
rect 44492 46620 44548 46622
rect 45836 50594 45892 50596
rect 45836 50542 45838 50594
rect 45838 50542 45890 50594
rect 45890 50542 45892 50594
rect 45836 50540 45892 50542
rect 46396 54514 46452 54516
rect 46396 54462 46398 54514
rect 46398 54462 46450 54514
rect 46450 54462 46452 54514
rect 46396 54460 46452 54462
rect 46956 54460 47012 54516
rect 46844 54402 46900 54404
rect 46844 54350 46846 54402
rect 46846 54350 46898 54402
rect 46898 54350 46900 54402
rect 46844 54348 46900 54350
rect 47852 54348 47908 54404
rect 47852 53788 47908 53844
rect 47516 53228 47572 53284
rect 46844 53170 46900 53172
rect 46844 53118 46846 53170
rect 46846 53118 46898 53170
rect 46898 53118 46900 53170
rect 46844 53116 46900 53118
rect 46396 52946 46452 52948
rect 46396 52894 46398 52946
rect 46398 52894 46450 52946
rect 46450 52894 46452 52946
rect 46396 52892 46452 52894
rect 46732 52892 46788 52948
rect 46508 52834 46564 52836
rect 46508 52782 46510 52834
rect 46510 52782 46562 52834
rect 46562 52782 46564 52834
rect 46508 52780 46564 52782
rect 46732 52274 46788 52276
rect 46732 52222 46734 52274
rect 46734 52222 46786 52274
rect 46786 52222 46788 52274
rect 46732 52220 46788 52222
rect 47180 52668 47236 52724
rect 47516 52892 47572 52948
rect 47292 51378 47348 51380
rect 47292 51326 47294 51378
rect 47294 51326 47346 51378
rect 47346 51326 47348 51378
rect 47292 51324 47348 51326
rect 46060 50540 46116 50596
rect 46732 50594 46788 50596
rect 46732 50542 46734 50594
rect 46734 50542 46786 50594
rect 46786 50542 46788 50594
rect 46732 50540 46788 50542
rect 50988 60620 51044 60676
rect 51324 63922 51380 63924
rect 51324 63870 51326 63922
rect 51326 63870 51378 63922
rect 51378 63870 51380 63922
rect 51324 63868 51380 63870
rect 52108 64428 52164 64484
rect 51660 62242 51716 62244
rect 51660 62190 51662 62242
rect 51662 62190 51714 62242
rect 51714 62190 51716 62242
rect 51660 62188 51716 62190
rect 51436 60956 51492 61012
rect 51212 60172 51268 60228
rect 51660 60732 51716 60788
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50428 59442 50484 59444
rect 50428 59390 50430 59442
rect 50430 59390 50482 59442
rect 50482 59390 50484 59442
rect 50428 59388 50484 59390
rect 49420 57372 49476 57428
rect 49868 58828 49924 58884
rect 49308 55132 49364 55188
rect 49532 55074 49588 55076
rect 49532 55022 49534 55074
rect 49534 55022 49586 55074
rect 49586 55022 49588 55074
rect 49532 55020 49588 55022
rect 49196 54572 49252 54628
rect 47964 53228 48020 53284
rect 47628 50540 47684 50596
rect 45276 48188 45332 48244
rect 45276 46956 45332 47012
rect 45052 46508 45108 46564
rect 45388 46674 45444 46676
rect 45388 46622 45390 46674
rect 45390 46622 45442 46674
rect 45442 46622 45444 46674
rect 45388 46620 45444 46622
rect 45948 46956 46004 47012
rect 45724 46674 45780 46676
rect 45724 46622 45726 46674
rect 45726 46622 45778 46674
rect 45778 46622 45780 46674
rect 45724 46620 45780 46622
rect 45836 46562 45892 46564
rect 45836 46510 45838 46562
rect 45838 46510 45890 46562
rect 45890 46510 45892 46562
rect 45836 46508 45892 46510
rect 44940 44828 44996 44884
rect 43372 44044 43428 44100
rect 43036 43372 43092 43428
rect 44940 43426 44996 43428
rect 44940 43374 44942 43426
rect 44942 43374 44994 43426
rect 44994 43374 44996 43426
rect 44940 43372 44996 43374
rect 43484 42924 43540 42980
rect 44156 42924 44212 42980
rect 45276 42476 45332 42532
rect 43932 42364 43988 42420
rect 44492 41916 44548 41972
rect 43484 40684 43540 40740
rect 43820 40124 43876 40180
rect 43372 39618 43428 39620
rect 43372 39566 43374 39618
rect 43374 39566 43426 39618
rect 43426 39566 43428 39618
rect 43372 39564 43428 39566
rect 45612 42978 45668 42980
rect 45612 42926 45614 42978
rect 45614 42926 45666 42978
rect 45666 42926 45668 42978
rect 45612 42924 45668 42926
rect 45612 42700 45668 42756
rect 45500 42364 45556 42420
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 49980 56306 50036 56308
rect 49980 56254 49982 56306
rect 49982 56254 50034 56306
rect 50034 56254 50036 56306
rect 49980 56252 50036 56254
rect 50316 56252 50372 56308
rect 51100 57538 51156 57540
rect 51100 57486 51102 57538
rect 51102 57486 51154 57538
rect 51154 57486 51156 57538
rect 51100 57484 51156 57486
rect 50316 56082 50372 56084
rect 50316 56030 50318 56082
rect 50318 56030 50370 56082
rect 50370 56030 50372 56082
rect 50316 56028 50372 56030
rect 49980 55186 50036 55188
rect 49980 55134 49982 55186
rect 49982 55134 50034 55186
rect 50034 55134 50036 55186
rect 49980 55132 50036 55134
rect 50316 54460 50372 54516
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 50876 56252 50932 56308
rect 50428 55020 50484 55076
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50876 54514 50932 54516
rect 50876 54462 50878 54514
rect 50878 54462 50930 54514
rect 50930 54462 50932 54514
rect 50876 54460 50932 54462
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50988 53004 51044 53060
rect 51436 59388 51492 59444
rect 54124 65378 54180 65380
rect 54124 65326 54126 65378
rect 54126 65326 54178 65378
rect 54178 65326 54180 65378
rect 54124 65324 54180 65326
rect 52780 64482 52836 64484
rect 52780 64430 52782 64482
rect 52782 64430 52834 64482
rect 52834 64430 52836 64482
rect 52780 64428 52836 64430
rect 54012 64482 54068 64484
rect 54012 64430 54014 64482
rect 54014 64430 54066 64482
rect 54066 64430 54068 64482
rect 54012 64428 54068 64430
rect 53004 63250 53060 63252
rect 53004 63198 53006 63250
rect 53006 63198 53058 63250
rect 53058 63198 53060 63250
rect 53004 63196 53060 63198
rect 52108 62578 52164 62580
rect 52108 62526 52110 62578
rect 52110 62526 52162 62578
rect 52162 62526 52164 62578
rect 52108 62524 52164 62526
rect 52444 62466 52500 62468
rect 52444 62414 52446 62466
rect 52446 62414 52498 62466
rect 52498 62414 52500 62466
rect 52444 62412 52500 62414
rect 52892 62242 52948 62244
rect 52892 62190 52894 62242
rect 52894 62190 52946 62242
rect 52946 62190 52948 62242
rect 52892 62188 52948 62190
rect 53900 63250 53956 63252
rect 53900 63198 53902 63250
rect 53902 63198 53954 63250
rect 53954 63198 53956 63250
rect 53900 63196 53956 63198
rect 53228 62412 53284 62468
rect 53004 60786 53060 60788
rect 53004 60734 53006 60786
rect 53006 60734 53058 60786
rect 53058 60734 53060 60786
rect 53004 60732 53060 60734
rect 54124 62188 54180 62244
rect 54908 65324 54964 65380
rect 55020 65436 55076 65492
rect 54572 64146 54628 64148
rect 54572 64094 54574 64146
rect 54574 64094 54626 64146
rect 54626 64094 54628 64146
rect 54572 64092 54628 64094
rect 54908 64428 54964 64484
rect 54684 63810 54740 63812
rect 54684 63758 54686 63810
rect 54686 63758 54738 63810
rect 54738 63758 54740 63810
rect 54684 63756 54740 63758
rect 54460 63532 54516 63588
rect 55020 63980 55076 64036
rect 56028 66498 56084 66500
rect 56028 66446 56030 66498
rect 56030 66446 56082 66498
rect 56082 66446 56084 66498
rect 56028 66444 56084 66446
rect 58156 66108 58212 66164
rect 57148 65436 57204 65492
rect 57596 65490 57652 65492
rect 57596 65438 57598 65490
rect 57598 65438 57650 65490
rect 57650 65438 57652 65490
rect 57596 65436 57652 65438
rect 55356 65324 55412 65380
rect 55244 64876 55300 64932
rect 55468 65212 55524 65268
rect 55356 64428 55412 64484
rect 55244 63980 55300 64036
rect 55132 63756 55188 63812
rect 54460 61068 54516 61124
rect 53340 60786 53396 60788
rect 53340 60734 53342 60786
rect 53342 60734 53394 60786
rect 53394 60734 53396 60786
rect 53340 60732 53396 60734
rect 54684 60786 54740 60788
rect 54684 60734 54686 60786
rect 54686 60734 54738 60786
rect 54738 60734 54740 60786
rect 54684 60732 54740 60734
rect 52780 60620 52836 60676
rect 51884 60172 51940 60228
rect 55020 63644 55076 63700
rect 55244 63250 55300 63252
rect 55244 63198 55246 63250
rect 55246 63198 55298 63250
rect 55298 63198 55300 63250
rect 55244 63196 55300 63198
rect 55804 63532 55860 63588
rect 55468 61570 55524 61572
rect 55468 61518 55470 61570
rect 55470 61518 55522 61570
rect 55522 61518 55524 61570
rect 55468 61516 55524 61518
rect 51436 57650 51492 57652
rect 51436 57598 51438 57650
rect 51438 57598 51490 57650
rect 51490 57598 51492 57650
rect 51436 57596 51492 57598
rect 51436 56028 51492 56084
rect 51324 54684 51380 54740
rect 52108 60002 52164 60004
rect 52108 59950 52110 60002
rect 52110 59950 52162 60002
rect 52162 59950 52164 60002
rect 52108 59948 52164 59950
rect 53340 59948 53396 60004
rect 52556 58268 52612 58324
rect 53004 58268 53060 58324
rect 51996 56476 52052 56532
rect 52780 56476 52836 56532
rect 51884 56028 51940 56084
rect 55244 61068 55300 61124
rect 54236 59948 54292 60004
rect 54908 59948 54964 60004
rect 54684 59442 54740 59444
rect 54684 59390 54686 59442
rect 54686 59390 54738 59442
rect 54738 59390 54740 59442
rect 54684 59388 54740 59390
rect 56364 63756 56420 63812
rect 56588 63698 56644 63700
rect 56588 63646 56590 63698
rect 56590 63646 56642 63698
rect 56642 63646 56644 63698
rect 56588 63644 56644 63646
rect 56700 63532 56756 63588
rect 56924 60844 56980 60900
rect 57372 61068 57428 61124
rect 57372 60898 57428 60900
rect 57372 60846 57374 60898
rect 57374 60846 57426 60898
rect 57426 60846 57428 60898
rect 57372 60844 57428 60846
rect 56028 59442 56084 59444
rect 56028 59390 56030 59442
rect 56030 59390 56082 59442
rect 56082 59390 56084 59442
rect 56028 59388 56084 59390
rect 57708 60786 57764 60788
rect 57708 60734 57710 60786
rect 57710 60734 57762 60786
rect 57762 60734 57764 60786
rect 57708 60732 57764 60734
rect 58156 65490 58212 65492
rect 58156 65438 58158 65490
rect 58158 65438 58210 65490
rect 58210 65438 58212 65490
rect 58156 65436 58212 65438
rect 58044 64428 58100 64484
rect 57932 61068 57988 61124
rect 56924 60562 56980 60564
rect 56924 60510 56926 60562
rect 56926 60510 56978 60562
rect 56978 60510 56980 60562
rect 56924 60508 56980 60510
rect 56924 59388 56980 59444
rect 51884 54738 51940 54740
rect 51884 54686 51886 54738
rect 51886 54686 51938 54738
rect 51938 54686 51940 54738
rect 51884 54684 51940 54686
rect 51660 54514 51716 54516
rect 51660 54462 51662 54514
rect 51662 54462 51714 54514
rect 51714 54462 51716 54514
rect 51660 54460 51716 54462
rect 51660 53900 51716 53956
rect 52668 53954 52724 53956
rect 52668 53902 52670 53954
rect 52670 53902 52722 53954
rect 52722 53902 52724 53954
rect 52668 53900 52724 53902
rect 52892 55074 52948 55076
rect 52892 55022 52894 55074
rect 52894 55022 52946 55074
rect 52946 55022 52948 55074
rect 52892 55020 52948 55022
rect 53116 54684 53172 54740
rect 53788 55020 53844 55076
rect 52780 53788 52836 53844
rect 53004 53842 53060 53844
rect 53004 53790 53006 53842
rect 53006 53790 53058 53842
rect 53058 53790 53060 53842
rect 53004 53788 53060 53790
rect 51660 53506 51716 53508
rect 51660 53454 51662 53506
rect 51662 53454 51714 53506
rect 51714 53454 51716 53506
rect 51660 53452 51716 53454
rect 51548 53116 51604 53172
rect 51660 53004 51716 53060
rect 51324 52668 51380 52724
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 47404 49586 47460 49588
rect 47404 49534 47406 49586
rect 47406 49534 47458 49586
rect 47458 49534 47460 49586
rect 47404 49532 47460 49534
rect 48860 49532 48916 49588
rect 47964 48076 48020 48132
rect 47740 47180 47796 47236
rect 47628 46844 47684 46900
rect 47628 46508 47684 46564
rect 47852 46396 47908 46452
rect 46620 43372 46676 43428
rect 46844 43372 46900 43428
rect 46620 42754 46676 42756
rect 46620 42702 46622 42754
rect 46622 42702 46674 42754
rect 46674 42702 46676 42754
rect 46620 42700 46676 42702
rect 45948 42476 46004 42532
rect 46396 42530 46452 42532
rect 46396 42478 46398 42530
rect 46398 42478 46450 42530
rect 46450 42478 46452 42530
rect 46396 42476 46452 42478
rect 45724 41804 45780 41860
rect 46844 41804 46900 41860
rect 45164 41020 45220 41076
rect 45164 40684 45220 40740
rect 44716 39788 44772 39844
rect 44268 39506 44324 39508
rect 44268 39454 44270 39506
rect 44270 39454 44322 39506
rect 44322 39454 44324 39506
rect 44268 39452 44324 39454
rect 43036 37154 43092 37156
rect 43036 37102 43038 37154
rect 43038 37102 43090 37154
rect 43090 37102 43092 37154
rect 43036 37100 43092 37102
rect 42700 36876 42756 36932
rect 42588 35196 42644 35252
rect 47740 40236 47796 40292
rect 47404 40124 47460 40180
rect 45836 39842 45892 39844
rect 45836 39790 45838 39842
rect 45838 39790 45890 39842
rect 45890 39790 45892 39842
rect 45836 39788 45892 39790
rect 45052 39506 45108 39508
rect 45052 39454 45054 39506
rect 45054 39454 45106 39506
rect 45106 39454 45108 39506
rect 45052 39452 45108 39454
rect 45724 39506 45780 39508
rect 45724 39454 45726 39506
rect 45726 39454 45778 39506
rect 45778 39454 45780 39506
rect 45724 39452 45780 39454
rect 46172 38722 46228 38724
rect 46172 38670 46174 38722
rect 46174 38670 46226 38722
rect 46226 38670 46228 38722
rect 46172 38668 46228 38670
rect 45724 38108 45780 38164
rect 46396 38162 46452 38164
rect 46396 38110 46398 38162
rect 46398 38110 46450 38162
rect 46450 38110 46452 38162
rect 46396 38108 46452 38110
rect 46060 37996 46116 38052
rect 46508 37884 46564 37940
rect 43708 35196 43764 35252
rect 44716 35196 44772 35252
rect 43932 34914 43988 34916
rect 43932 34862 43934 34914
rect 43934 34862 43986 34914
rect 43986 34862 43988 34914
rect 43932 34860 43988 34862
rect 44268 34860 44324 34916
rect 42700 34412 42756 34468
rect 43596 34412 43652 34468
rect 44492 34412 44548 34468
rect 44604 34130 44660 34132
rect 44604 34078 44606 34130
rect 44606 34078 44658 34130
rect 44658 34078 44660 34130
rect 44604 34076 44660 34078
rect 45052 34076 45108 34132
rect 43372 33180 43428 33236
rect 43596 32450 43652 32452
rect 43596 32398 43598 32450
rect 43598 32398 43650 32450
rect 43650 32398 43652 32450
rect 43596 32396 43652 32398
rect 42588 32284 42644 32340
rect 41692 30828 41748 30884
rect 41468 29260 41524 29316
rect 40908 28476 40964 28532
rect 41132 27858 41188 27860
rect 41132 27806 41134 27858
rect 41134 27806 41186 27858
rect 41186 27806 41188 27858
rect 41132 27804 41188 27806
rect 40908 27132 40964 27188
rect 42364 30156 42420 30212
rect 44044 32450 44100 32452
rect 44044 32398 44046 32450
rect 44046 32398 44098 32450
rect 44098 32398 44100 32450
rect 44044 32396 44100 32398
rect 46172 37212 46228 37268
rect 45836 36988 45892 37044
rect 45500 35698 45556 35700
rect 45500 35646 45502 35698
rect 45502 35646 45554 35698
rect 45554 35646 45556 35698
rect 45500 35644 45556 35646
rect 45500 35196 45556 35252
rect 45724 34130 45780 34132
rect 45724 34078 45726 34130
rect 45726 34078 45778 34130
rect 45778 34078 45780 34130
rect 45724 34076 45780 34078
rect 44268 31778 44324 31780
rect 44268 31726 44270 31778
rect 44270 31726 44322 31778
rect 44322 31726 44324 31778
rect 44268 31724 44324 31726
rect 41916 29932 41972 29988
rect 41804 29148 41860 29204
rect 41916 27804 41972 27860
rect 41916 27186 41972 27188
rect 41916 27134 41918 27186
rect 41918 27134 41970 27186
rect 41970 27134 41972 27186
rect 41916 27132 41972 27134
rect 40124 26514 40180 26516
rect 40124 26462 40126 26514
rect 40126 26462 40178 26514
rect 40178 26462 40180 26514
rect 40124 26460 40180 26462
rect 39676 26124 39732 26180
rect 39788 26012 39844 26068
rect 40348 25676 40404 25732
rect 40124 25506 40180 25508
rect 40124 25454 40126 25506
rect 40126 25454 40178 25506
rect 40178 25454 40180 25506
rect 40124 25452 40180 25454
rect 39564 25116 39620 25172
rect 38108 23212 38164 23268
rect 37884 23100 37940 23156
rect 37324 22258 37380 22260
rect 37324 22206 37326 22258
rect 37326 22206 37378 22258
rect 37378 22206 37380 22258
rect 37324 22204 37380 22206
rect 36988 19404 37044 19460
rect 37100 19180 37156 19236
rect 37212 20188 37268 20244
rect 37772 20242 37828 20244
rect 37772 20190 37774 20242
rect 37774 20190 37826 20242
rect 37826 20190 37828 20242
rect 37772 20188 37828 20190
rect 37100 18508 37156 18564
rect 36876 18396 36932 18452
rect 37884 18732 37940 18788
rect 37212 17724 37268 17780
rect 37884 18284 37940 18340
rect 35980 16940 36036 16996
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34972 16268 35028 16324
rect 35532 16044 35588 16100
rect 38108 16604 38164 16660
rect 38444 23100 38500 23156
rect 38556 22540 38612 22596
rect 38444 22204 38500 22260
rect 38780 22428 38836 22484
rect 40236 23996 40292 24052
rect 40012 23660 40068 23716
rect 39228 23266 39284 23268
rect 39228 23214 39230 23266
rect 39230 23214 39282 23266
rect 39282 23214 39284 23266
rect 39228 23212 39284 23214
rect 38556 20188 38612 20244
rect 38332 19010 38388 19012
rect 38332 18958 38334 19010
rect 38334 18958 38386 19010
rect 38386 18958 38388 19010
rect 38332 18956 38388 18958
rect 38556 18956 38612 19012
rect 38780 19516 38836 19572
rect 38556 18338 38612 18340
rect 38556 18286 38558 18338
rect 38558 18286 38610 18338
rect 38610 18286 38612 18338
rect 38556 18284 38612 18286
rect 37884 16268 37940 16324
rect 36092 16044 36148 16100
rect 37772 15932 37828 15988
rect 37548 15708 37604 15764
rect 34860 14140 34916 14196
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 37100 14588 37156 14644
rect 33964 13020 34020 13076
rect 33292 11228 33348 11284
rect 32620 10780 32676 10836
rect 33516 11170 33572 11172
rect 33516 11118 33518 11170
rect 33518 11118 33570 11170
rect 33570 11118 33572 11170
rect 33516 11116 33572 11118
rect 33516 10892 33572 10948
rect 32732 9714 32788 9716
rect 32732 9662 32734 9714
rect 32734 9662 32786 9714
rect 32786 9662 32788 9714
rect 32732 9660 32788 9662
rect 32844 9212 32900 9268
rect 31164 8146 31220 8148
rect 31164 8094 31166 8146
rect 31166 8094 31218 8146
rect 31218 8094 31220 8146
rect 31164 8092 31220 8094
rect 32508 8370 32564 8372
rect 32508 8318 32510 8370
rect 32510 8318 32562 8370
rect 32562 8318 32564 8370
rect 32508 8316 32564 8318
rect 31612 8146 31668 8148
rect 31612 8094 31614 8146
rect 31614 8094 31666 8146
rect 31666 8094 31668 8146
rect 31612 8092 31668 8094
rect 30940 7644 30996 7700
rect 31500 7698 31556 7700
rect 31500 7646 31502 7698
rect 31502 7646 31554 7698
rect 31554 7646 31556 7698
rect 31500 7644 31556 7646
rect 31724 7308 31780 7364
rect 31836 6636 31892 6692
rect 30716 6076 30772 6132
rect 31276 6188 31332 6244
rect 30828 5964 30884 6020
rect 30828 5516 30884 5572
rect 30940 5180 30996 5236
rect 30828 5122 30884 5124
rect 30828 5070 30830 5122
rect 30830 5070 30882 5122
rect 30882 5070 30884 5122
rect 30828 5068 30884 5070
rect 30492 4508 30548 4564
rect 31500 5404 31556 5460
rect 32396 6636 32452 6692
rect 31948 6524 32004 6580
rect 32284 6524 32340 6580
rect 32060 6188 32116 6244
rect 32172 5628 32228 5684
rect 33292 9884 33348 9940
rect 33404 9996 33460 10052
rect 33180 9826 33236 9828
rect 33180 9774 33182 9826
rect 33182 9774 33234 9826
rect 33234 9774 33236 9826
rect 33180 9772 33236 9774
rect 33740 9884 33796 9940
rect 33292 9660 33348 9716
rect 33292 9324 33348 9380
rect 33964 11564 34020 11620
rect 34076 9772 34132 9828
rect 33852 9266 33908 9268
rect 33852 9214 33854 9266
rect 33854 9214 33906 9266
rect 33906 9214 33908 9266
rect 33852 9212 33908 9214
rect 34636 13074 34692 13076
rect 34636 13022 34638 13074
rect 34638 13022 34690 13074
rect 34690 13022 34692 13074
rect 34636 13020 34692 13022
rect 34524 12402 34580 12404
rect 34524 12350 34526 12402
rect 34526 12350 34578 12402
rect 34578 12350 34580 12402
rect 34524 12348 34580 12350
rect 34300 12012 34356 12068
rect 34972 13132 35028 13188
rect 35308 13468 35364 13524
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35084 13020 35140 13076
rect 34860 12962 34916 12964
rect 34860 12910 34862 12962
rect 34862 12910 34914 12962
rect 34914 12910 34916 12962
rect 34860 12908 34916 12910
rect 35868 13916 35924 13972
rect 35756 13468 35812 13524
rect 35196 12348 35252 12404
rect 35644 13132 35700 13188
rect 35532 12460 35588 12516
rect 34636 11900 34692 11956
rect 35084 12012 35140 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35532 11452 35588 11508
rect 35532 11228 35588 11284
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34524 9772 34580 9828
rect 34412 9100 34468 9156
rect 34188 8428 34244 8484
rect 33964 7980 34020 8036
rect 33852 7586 33908 7588
rect 33852 7534 33854 7586
rect 33854 7534 33906 7586
rect 33906 7534 33908 7586
rect 33852 7532 33908 7534
rect 34188 7474 34244 7476
rect 34188 7422 34190 7474
rect 34190 7422 34242 7474
rect 34242 7422 34244 7474
rect 34188 7420 34244 7422
rect 32620 6524 32676 6580
rect 33628 6300 33684 6356
rect 35644 9826 35700 9828
rect 35644 9774 35646 9826
rect 35646 9774 35698 9826
rect 35698 9774 35700 9826
rect 35644 9772 35700 9774
rect 35868 13020 35924 13076
rect 37884 15874 37940 15876
rect 37884 15822 37886 15874
rect 37886 15822 37938 15874
rect 37938 15822 37940 15874
rect 37884 15820 37940 15822
rect 38332 16268 38388 16324
rect 38556 15820 38612 15876
rect 38444 15314 38500 15316
rect 38444 15262 38446 15314
rect 38446 15262 38498 15314
rect 38498 15262 38500 15314
rect 38444 15260 38500 15262
rect 37212 13468 37268 13524
rect 37548 13468 37604 13524
rect 37100 13074 37156 13076
rect 37100 13022 37102 13074
rect 37102 13022 37154 13074
rect 37154 13022 37156 13074
rect 37100 13020 37156 13022
rect 36316 12962 36372 12964
rect 36316 12910 36318 12962
rect 36318 12910 36370 12962
rect 36370 12910 36372 12962
rect 36316 12908 36372 12910
rect 35868 12572 35924 12628
rect 35980 12460 36036 12516
rect 37660 11900 37716 11956
rect 35084 9042 35140 9044
rect 35084 8990 35086 9042
rect 35086 8990 35138 9042
rect 35138 8990 35140 9042
rect 35084 8988 35140 8990
rect 32060 5068 32116 5124
rect 34972 8034 35028 8036
rect 34972 7982 34974 8034
rect 34974 7982 35026 8034
rect 35026 7982 35028 8034
rect 34972 7980 35028 7982
rect 34972 7196 35028 7252
rect 35532 9154 35588 9156
rect 35532 9102 35534 9154
rect 35534 9102 35586 9154
rect 35586 9102 35588 9154
rect 35532 9100 35588 9102
rect 36092 9826 36148 9828
rect 36092 9774 36094 9826
rect 36094 9774 36146 9826
rect 36146 9774 36148 9826
rect 36092 9772 36148 9774
rect 37100 9772 37156 9828
rect 36540 9714 36596 9716
rect 36540 9662 36542 9714
rect 36542 9662 36594 9714
rect 36594 9662 36596 9714
rect 36540 9660 36596 9662
rect 38332 14700 38388 14756
rect 37884 13468 37940 13524
rect 38444 13468 38500 13524
rect 38108 11900 38164 11956
rect 38332 11506 38388 11508
rect 38332 11454 38334 11506
rect 38334 11454 38386 11506
rect 38386 11454 38388 11506
rect 38332 11452 38388 11454
rect 37884 11282 37940 11284
rect 37884 11230 37886 11282
rect 37886 11230 37938 11282
rect 37938 11230 37940 11282
rect 37884 11228 37940 11230
rect 38892 19010 38948 19012
rect 38892 18958 38894 19010
rect 38894 18958 38946 19010
rect 38946 18958 38948 19010
rect 38892 18956 38948 18958
rect 39340 19292 39396 19348
rect 39788 19346 39844 19348
rect 39788 19294 39790 19346
rect 39790 19294 39842 19346
rect 39842 19294 39844 19346
rect 39788 19292 39844 19294
rect 39564 18732 39620 18788
rect 39788 17724 39844 17780
rect 39116 16604 39172 16660
rect 39564 15820 39620 15876
rect 39564 15314 39620 15316
rect 39564 15262 39566 15314
rect 39566 15262 39618 15314
rect 39618 15262 39620 15314
rect 39564 15260 39620 15262
rect 39004 13692 39060 13748
rect 38780 12738 38836 12740
rect 38780 12686 38782 12738
rect 38782 12686 38834 12738
rect 38834 12686 38836 12738
rect 38780 12684 38836 12686
rect 39564 14418 39620 14420
rect 39564 14366 39566 14418
rect 39566 14366 39618 14418
rect 39618 14366 39620 14418
rect 39564 14364 39620 14366
rect 39116 13356 39172 13412
rect 39228 13244 39284 13300
rect 39004 12402 39060 12404
rect 39004 12350 39006 12402
rect 39006 12350 39058 12402
rect 39058 12350 39060 12402
rect 39004 12348 39060 12350
rect 39676 12684 39732 12740
rect 39676 12460 39732 12516
rect 39340 12348 39396 12404
rect 38780 11788 38836 11844
rect 39452 11452 39508 11508
rect 38668 11282 38724 11284
rect 38668 11230 38670 11282
rect 38670 11230 38722 11282
rect 38722 11230 38724 11282
rect 38668 11228 38724 11230
rect 39004 10108 39060 10164
rect 37324 9436 37380 9492
rect 35868 8988 35924 9044
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 36316 8204 36372 8260
rect 36764 8092 36820 8148
rect 35532 7644 35588 7700
rect 35644 7586 35700 7588
rect 35644 7534 35646 7586
rect 35646 7534 35698 7586
rect 35698 7534 35700 7586
rect 35644 7532 35700 7534
rect 34524 5180 34580 5236
rect 35420 7474 35476 7476
rect 35420 7422 35422 7474
rect 35422 7422 35474 7474
rect 35474 7422 35476 7474
rect 35420 7420 35476 7422
rect 36092 7644 36148 7700
rect 36428 7586 36484 7588
rect 36428 7534 36430 7586
rect 36430 7534 36482 7586
rect 36482 7534 36484 7586
rect 36428 7532 36484 7534
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35980 7250 36036 7252
rect 35980 7198 35982 7250
rect 35982 7198 36034 7250
rect 36034 7198 36036 7250
rect 35980 7196 36036 7198
rect 37660 9154 37716 9156
rect 37660 9102 37662 9154
rect 37662 9102 37714 9154
rect 37714 9102 37716 9154
rect 37660 9100 37716 9102
rect 39228 9154 39284 9156
rect 39228 9102 39230 9154
rect 39230 9102 39282 9154
rect 39282 9102 39284 9154
rect 39228 9100 39284 9102
rect 37436 7644 37492 7700
rect 39004 8034 39060 8036
rect 39004 7982 39006 8034
rect 39006 7982 39058 8034
rect 39058 7982 39060 8034
rect 39004 7980 39060 7982
rect 38892 7644 38948 7700
rect 38108 7474 38164 7476
rect 38108 7422 38110 7474
rect 38110 7422 38162 7474
rect 38162 7422 38164 7474
rect 38108 7420 38164 7422
rect 38668 7474 38724 7476
rect 38668 7422 38670 7474
rect 38670 7422 38722 7474
rect 38722 7422 38724 7474
rect 38668 7420 38724 7422
rect 38220 7308 38276 7364
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 5234 35700 5236
rect 35644 5182 35646 5234
rect 35646 5182 35698 5234
rect 35698 5182 35700 5234
rect 35644 5180 35700 5182
rect 37996 6972 38052 7028
rect 38780 6972 38836 7028
rect 39116 7474 39172 7476
rect 39116 7422 39118 7474
rect 39118 7422 39170 7474
rect 39170 7422 39172 7474
rect 39116 7420 39172 7422
rect 39004 6860 39060 6916
rect 39340 7308 39396 7364
rect 39340 6636 39396 6692
rect 38556 6578 38612 6580
rect 38556 6526 38558 6578
rect 38558 6526 38610 6578
rect 38610 6526 38612 6578
rect 38556 6524 38612 6526
rect 37660 5292 37716 5348
rect 40348 21810 40404 21812
rect 40348 21758 40350 21810
rect 40350 21758 40402 21810
rect 40402 21758 40404 21810
rect 40348 21756 40404 21758
rect 40348 20130 40404 20132
rect 40348 20078 40350 20130
rect 40350 20078 40402 20130
rect 40402 20078 40404 20130
rect 40348 20076 40404 20078
rect 40348 19180 40404 19236
rect 40236 18844 40292 18900
rect 40236 18284 40292 18340
rect 41916 26514 41972 26516
rect 41916 26462 41918 26514
rect 41918 26462 41970 26514
rect 41970 26462 41972 26514
rect 41916 26460 41972 26462
rect 41468 26402 41524 26404
rect 41468 26350 41470 26402
rect 41470 26350 41522 26402
rect 41522 26350 41524 26402
rect 41468 26348 41524 26350
rect 40684 26236 40740 26292
rect 41132 26290 41188 26292
rect 41132 26238 41134 26290
rect 41134 26238 41186 26290
rect 41186 26238 41188 26290
rect 41132 26236 41188 26238
rect 41020 26066 41076 26068
rect 41020 26014 41022 26066
rect 41022 26014 41074 26066
rect 41074 26014 41076 26066
rect 41020 26012 41076 26014
rect 40684 25452 40740 25508
rect 40572 25394 40628 25396
rect 40572 25342 40574 25394
rect 40574 25342 40626 25394
rect 40626 25342 40628 25394
rect 40572 25340 40628 25342
rect 41356 25340 41412 25396
rect 41468 25282 41524 25284
rect 41468 25230 41470 25282
rect 41470 25230 41522 25282
rect 41522 25230 41524 25282
rect 41468 25228 41524 25230
rect 41132 24834 41188 24836
rect 41132 24782 41134 24834
rect 41134 24782 41186 24834
rect 41186 24782 41188 24834
rect 41132 24780 41188 24782
rect 40460 14588 40516 14644
rect 41244 23436 41300 23492
rect 41020 23154 41076 23156
rect 41020 23102 41022 23154
rect 41022 23102 41074 23154
rect 41074 23102 41076 23154
rect 41020 23100 41076 23102
rect 40684 22482 40740 22484
rect 40684 22430 40686 22482
rect 40686 22430 40738 22482
rect 40738 22430 40740 22482
rect 40684 22428 40740 22430
rect 41468 22204 41524 22260
rect 41580 21756 41636 21812
rect 41244 20130 41300 20132
rect 41244 20078 41246 20130
rect 41246 20078 41298 20130
rect 41298 20078 41300 20130
rect 41244 20076 41300 20078
rect 41468 20018 41524 20020
rect 41468 19966 41470 20018
rect 41470 19966 41522 20018
rect 41522 19966 41524 20018
rect 41468 19964 41524 19966
rect 41916 25228 41972 25284
rect 42140 25004 42196 25060
rect 41804 24722 41860 24724
rect 41804 24670 41806 24722
rect 41806 24670 41858 24722
rect 41858 24670 41860 24722
rect 41804 24668 41860 24670
rect 42812 29202 42868 29204
rect 42812 29150 42814 29202
rect 42814 29150 42866 29202
rect 42866 29150 42868 29202
rect 42812 29148 42868 29150
rect 42588 27132 42644 27188
rect 42476 25394 42532 25396
rect 42476 25342 42478 25394
rect 42478 25342 42530 25394
rect 42530 25342 42532 25394
rect 42476 25340 42532 25342
rect 42700 24722 42756 24724
rect 42700 24670 42702 24722
rect 42702 24670 42754 24722
rect 42754 24670 42756 24722
rect 42700 24668 42756 24670
rect 43372 28418 43428 28420
rect 43372 28366 43374 28418
rect 43374 28366 43426 28418
rect 43426 28366 43428 28418
rect 43372 28364 43428 28366
rect 44044 28364 44100 28420
rect 44380 28700 44436 28756
rect 43932 26850 43988 26852
rect 43932 26798 43934 26850
rect 43934 26798 43986 26850
rect 43986 26798 43988 26850
rect 43932 26796 43988 26798
rect 43708 26460 43764 26516
rect 43036 25004 43092 25060
rect 43708 25340 43764 25396
rect 43372 24668 43428 24724
rect 42924 23548 42980 23604
rect 43260 23772 43316 23828
rect 42252 23154 42308 23156
rect 42252 23102 42254 23154
rect 42254 23102 42306 23154
rect 42306 23102 42308 23154
rect 42252 23100 42308 23102
rect 42028 22258 42084 22260
rect 42028 22206 42030 22258
rect 42030 22206 42082 22258
rect 42082 22206 42084 22258
rect 42028 22204 42084 22206
rect 41020 19906 41076 19908
rect 41020 19854 41022 19906
rect 41022 19854 41074 19906
rect 41074 19854 41076 19906
rect 41020 19852 41076 19854
rect 40908 19516 40964 19572
rect 41244 18732 41300 18788
rect 40908 18508 40964 18564
rect 41356 18450 41412 18452
rect 41356 18398 41358 18450
rect 41358 18398 41410 18450
rect 41410 18398 41412 18450
rect 41356 18396 41412 18398
rect 41468 17836 41524 17892
rect 40684 17778 40740 17780
rect 40684 17726 40686 17778
rect 40686 17726 40738 17778
rect 40738 17726 40740 17778
rect 40684 17724 40740 17726
rect 41804 18284 41860 18340
rect 41692 17612 41748 17668
rect 41020 16268 41076 16324
rect 41020 15260 41076 15316
rect 40572 13468 40628 13524
rect 40908 14418 40964 14420
rect 40908 14366 40910 14418
rect 40910 14366 40962 14418
rect 40962 14366 40964 14418
rect 40908 14364 40964 14366
rect 40012 13356 40068 13412
rect 39900 13244 39956 13300
rect 41132 15820 41188 15876
rect 42140 19964 42196 20020
rect 42588 19906 42644 19908
rect 42588 19854 42590 19906
rect 42590 19854 42642 19906
rect 42642 19854 42644 19906
rect 42588 19852 42644 19854
rect 42252 19404 42308 19460
rect 42028 19010 42084 19012
rect 42028 18958 42030 19010
rect 42030 18958 42082 19010
rect 42082 18958 42084 19010
rect 42028 18956 42084 18958
rect 42364 18620 42420 18676
rect 42140 18562 42196 18564
rect 42140 18510 42142 18562
rect 42142 18510 42194 18562
rect 42194 18510 42196 18562
rect 42140 18508 42196 18510
rect 43148 18620 43204 18676
rect 42588 18450 42644 18452
rect 42588 18398 42590 18450
rect 42590 18398 42642 18450
rect 42642 18398 42644 18450
rect 42588 18396 42644 18398
rect 43036 18172 43092 18228
rect 41916 15708 41972 15764
rect 41916 15314 41972 15316
rect 41916 15262 41918 15314
rect 41918 15262 41970 15314
rect 41970 15262 41972 15314
rect 41916 15260 41972 15262
rect 41468 14642 41524 14644
rect 41468 14590 41470 14642
rect 41470 14590 41522 14642
rect 41522 14590 41524 14642
rect 41468 14588 41524 14590
rect 41692 15036 41748 15092
rect 41916 14530 41972 14532
rect 41916 14478 41918 14530
rect 41918 14478 41970 14530
rect 41970 14478 41972 14530
rect 41916 14476 41972 14478
rect 41468 14252 41524 14308
rect 40236 12012 40292 12068
rect 41132 13804 41188 13860
rect 41916 13916 41972 13972
rect 41132 12796 41188 12852
rect 42812 15036 42868 15092
rect 42588 14588 42644 14644
rect 42700 14306 42756 14308
rect 42700 14254 42702 14306
rect 42702 14254 42754 14306
rect 42754 14254 42756 14306
rect 42700 14252 42756 14254
rect 42140 13634 42196 13636
rect 42140 13582 42142 13634
rect 42142 13582 42194 13634
rect 42194 13582 42196 13634
rect 42140 13580 42196 13582
rect 42028 12850 42084 12852
rect 42028 12798 42030 12850
rect 42030 12798 42082 12850
rect 42082 12798 42084 12850
rect 42028 12796 42084 12798
rect 42476 13468 42532 13524
rect 42140 12460 42196 12516
rect 42364 13244 42420 13300
rect 41692 11788 41748 11844
rect 42140 12066 42196 12068
rect 42140 12014 42142 12066
rect 42142 12014 42194 12066
rect 42194 12014 42196 12066
rect 42140 12012 42196 12014
rect 41020 11452 41076 11508
rect 39676 10892 39732 10948
rect 40236 10108 40292 10164
rect 42364 12348 42420 12404
rect 42252 11004 42308 11060
rect 42252 10498 42308 10500
rect 42252 10446 42254 10498
rect 42254 10446 42306 10498
rect 42306 10446 42308 10498
rect 42252 10444 42308 10446
rect 42140 10332 42196 10388
rect 41804 10108 41860 10164
rect 42252 9884 42308 9940
rect 40348 9714 40404 9716
rect 40348 9662 40350 9714
rect 40350 9662 40402 9714
rect 40402 9662 40404 9714
rect 40348 9660 40404 9662
rect 39788 9100 39844 9156
rect 39564 7756 39620 7812
rect 39676 8034 39732 8036
rect 39676 7982 39678 8034
rect 39678 7982 39730 8034
rect 39730 7982 39732 8034
rect 39676 7980 39732 7982
rect 42588 12796 42644 12852
rect 42812 12348 42868 12404
rect 43036 14476 43092 14532
rect 43260 13970 43316 13972
rect 43260 13918 43262 13970
rect 43262 13918 43314 13970
rect 43314 13918 43316 13970
rect 43260 13916 43316 13918
rect 43372 12908 43428 12964
rect 43484 24556 43540 24612
rect 43596 24444 43652 24500
rect 43708 23772 43764 23828
rect 43596 23660 43652 23716
rect 43708 22204 43764 22260
rect 43596 18172 43652 18228
rect 44268 26962 44324 26964
rect 44268 26910 44270 26962
rect 44270 26910 44322 26962
rect 44322 26910 44324 26962
rect 44268 26908 44324 26910
rect 43932 25730 43988 25732
rect 43932 25678 43934 25730
rect 43934 25678 43986 25730
rect 43986 25678 43988 25730
rect 43932 25676 43988 25678
rect 44044 23772 44100 23828
rect 44156 23378 44212 23380
rect 44156 23326 44158 23378
rect 44158 23326 44210 23378
rect 44210 23326 44212 23378
rect 44156 23324 44212 23326
rect 44156 23100 44212 23156
rect 44156 21868 44212 21924
rect 45388 31890 45444 31892
rect 45388 31838 45390 31890
rect 45390 31838 45442 31890
rect 45442 31838 45444 31890
rect 45388 31836 45444 31838
rect 45164 31724 45220 31780
rect 45276 30156 45332 30212
rect 45612 30156 45668 30212
rect 45276 28754 45332 28756
rect 45276 28702 45278 28754
rect 45278 28702 45330 28754
rect 45330 28702 45332 28754
rect 45276 28700 45332 28702
rect 44828 26796 44884 26852
rect 44940 25676 44996 25732
rect 45164 26908 45220 26964
rect 45052 25506 45108 25508
rect 45052 25454 45054 25506
rect 45054 25454 45106 25506
rect 45106 25454 45108 25506
rect 45052 25452 45108 25454
rect 44828 25228 44884 25284
rect 44828 24610 44884 24612
rect 44828 24558 44830 24610
rect 44830 24558 44882 24610
rect 44882 24558 44884 24610
rect 44828 24556 44884 24558
rect 45948 33516 46004 33572
rect 45948 25506 46004 25508
rect 45948 25454 45950 25506
rect 45950 25454 46002 25506
rect 46002 25454 46004 25506
rect 45948 25452 46004 25454
rect 45836 25228 45892 25284
rect 47740 35196 47796 35252
rect 47292 34300 47348 34356
rect 46732 32562 46788 32564
rect 46732 32510 46734 32562
rect 46734 32510 46786 32562
rect 46786 32510 46788 32562
rect 46732 32508 46788 32510
rect 47404 32562 47460 32564
rect 47404 32510 47406 32562
rect 47406 32510 47458 32562
rect 47458 32510 47460 32562
rect 47404 32508 47460 32510
rect 47516 31666 47572 31668
rect 47516 31614 47518 31666
rect 47518 31614 47570 31666
rect 47570 31614 47572 31666
rect 47516 31612 47572 31614
rect 46956 30322 47012 30324
rect 46956 30270 46958 30322
rect 46958 30270 47010 30322
rect 47010 30270 47012 30322
rect 46956 30268 47012 30270
rect 46508 29260 46564 29316
rect 46396 26348 46452 26404
rect 48860 48130 48916 48132
rect 48860 48078 48862 48130
rect 48862 48078 48914 48130
rect 48914 48078 48916 48130
rect 48860 48076 48916 48078
rect 48412 45890 48468 45892
rect 48412 45838 48414 45890
rect 48414 45838 48466 45890
rect 48466 45838 48468 45890
rect 48412 45836 48468 45838
rect 48076 45666 48132 45668
rect 48076 45614 48078 45666
rect 48078 45614 48130 45666
rect 48130 45614 48132 45666
rect 48076 45612 48132 45614
rect 48748 46786 48804 46788
rect 48748 46734 48750 46786
rect 48750 46734 48802 46786
rect 48802 46734 48804 46786
rect 48748 46732 48804 46734
rect 49196 48300 49252 48356
rect 49084 48188 49140 48244
rect 49196 48076 49252 48132
rect 49644 48188 49700 48244
rect 49756 47852 49812 47908
rect 49084 45218 49140 45220
rect 49084 45166 49086 45218
rect 49086 45166 49138 45218
rect 49138 45166 49140 45218
rect 49084 45164 49140 45166
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 49868 47404 49924 47460
rect 49308 46674 49364 46676
rect 49308 46622 49310 46674
rect 49310 46622 49362 46674
rect 49362 46622 49364 46674
rect 49308 46620 49364 46622
rect 49308 45724 49364 45780
rect 49756 46674 49812 46676
rect 49756 46622 49758 46674
rect 49758 46622 49810 46674
rect 49810 46622 49812 46674
rect 49756 46620 49812 46622
rect 49532 45836 49588 45892
rect 49980 48972 50036 49028
rect 50764 49922 50820 49924
rect 50764 49870 50766 49922
rect 50766 49870 50818 49922
rect 50818 49870 50820 49922
rect 50764 49868 50820 49870
rect 50876 49308 50932 49364
rect 50652 49026 50708 49028
rect 50652 48974 50654 49026
rect 50654 48974 50706 49026
rect 50706 48974 50708 49026
rect 50652 48972 50708 48974
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 51100 51100 51156 51156
rect 52780 53506 52836 53508
rect 52780 53454 52782 53506
rect 52782 53454 52834 53506
rect 52834 53454 52836 53506
rect 52780 53452 52836 53454
rect 53676 53452 53732 53508
rect 53900 55468 53956 55524
rect 53340 52220 53396 52276
rect 53228 52108 53284 52164
rect 51772 51154 51828 51156
rect 51772 51102 51774 51154
rect 51774 51102 51826 51154
rect 51826 51102 51828 51154
rect 51772 51100 51828 51102
rect 52444 51378 52500 51380
rect 52444 51326 52446 51378
rect 52446 51326 52498 51378
rect 52498 51326 52500 51378
rect 52444 51324 52500 51326
rect 51212 50652 51268 50708
rect 53228 50764 53284 50820
rect 52668 49868 52724 49924
rect 51660 49308 51716 49364
rect 51548 49026 51604 49028
rect 51548 48974 51550 49026
rect 51550 48974 51602 49026
rect 51602 48974 51604 49026
rect 51548 48972 51604 48974
rect 50092 47852 50148 47908
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50540 46674 50596 46676
rect 50540 46622 50542 46674
rect 50542 46622 50594 46674
rect 50594 46622 50596 46674
rect 50540 46620 50596 46622
rect 50092 46396 50148 46452
rect 49980 45778 50036 45780
rect 49980 45726 49982 45778
rect 49982 45726 50034 45778
rect 50034 45726 50036 45778
rect 49980 45724 50036 45726
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50988 45164 51044 45220
rect 49980 45106 50036 45108
rect 49980 45054 49982 45106
rect 49982 45054 50034 45106
rect 50034 45054 50036 45106
rect 49980 45052 50036 45054
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 48188 43426 48244 43428
rect 48188 43374 48190 43426
rect 48190 43374 48242 43426
rect 48242 43374 48244 43426
rect 48188 43372 48244 43374
rect 48188 40572 48244 40628
rect 48076 40290 48132 40292
rect 48076 40238 48078 40290
rect 48078 40238 48130 40290
rect 48130 40238 48132 40290
rect 48076 40236 48132 40238
rect 49084 41916 49140 41972
rect 49196 40348 49252 40404
rect 50204 42642 50260 42644
rect 50204 42590 50206 42642
rect 50206 42590 50258 42642
rect 50258 42590 50260 42642
rect 50204 42588 50260 42590
rect 49644 41916 49700 41972
rect 49868 41356 49924 41412
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50540 41356 50596 41412
rect 50876 40908 50932 40964
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 53676 52108 53732 52164
rect 54124 52162 54180 52164
rect 54124 52110 54126 52162
rect 54126 52110 54178 52162
rect 54178 52110 54180 52162
rect 54124 52108 54180 52110
rect 54012 50764 54068 50820
rect 54908 55468 54964 55524
rect 55132 55468 55188 55524
rect 55020 55244 55076 55300
rect 54796 54124 54852 54180
rect 54908 54290 54964 54292
rect 54908 54238 54910 54290
rect 54910 54238 54962 54290
rect 54962 54238 54964 54290
rect 54908 54236 54964 54238
rect 55132 54572 55188 54628
rect 55132 54124 55188 54180
rect 56476 55356 56532 55412
rect 55804 53788 55860 53844
rect 56140 54348 56196 54404
rect 56812 54572 56868 54628
rect 56700 54402 56756 54404
rect 56700 54350 56702 54402
rect 56702 54350 56754 54402
rect 56754 54350 56756 54402
rect 56700 54348 56756 54350
rect 56140 52386 56196 52388
rect 56140 52334 56142 52386
rect 56142 52334 56194 52386
rect 56194 52334 56196 52386
rect 56140 52332 56196 52334
rect 56588 52332 56644 52388
rect 55132 52108 55188 52164
rect 54684 51436 54740 51492
rect 54460 49868 54516 49924
rect 55468 51548 55524 51604
rect 55356 51212 55412 51268
rect 54908 49026 54964 49028
rect 54908 48974 54910 49026
rect 54910 48974 54962 49026
rect 54962 48974 54964 49026
rect 54908 48972 54964 48974
rect 54684 48636 54740 48692
rect 53900 48300 53956 48356
rect 54796 48300 54852 48356
rect 52108 46396 52164 46452
rect 54236 48130 54292 48132
rect 54236 48078 54238 48130
rect 54238 48078 54290 48130
rect 54290 48078 54292 48130
rect 54236 48076 54292 48078
rect 51884 44940 51940 44996
rect 51772 43708 51828 43764
rect 51436 42476 51492 42532
rect 50316 40348 50372 40404
rect 48860 39228 48916 39284
rect 47964 28924 48020 28980
rect 48524 37938 48580 37940
rect 48524 37886 48526 37938
rect 48526 37886 48578 37938
rect 48578 37886 48580 37938
rect 48524 37884 48580 37886
rect 48860 34972 48916 35028
rect 48188 34300 48244 34356
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 49420 38722 49476 38724
rect 49420 38670 49422 38722
rect 49422 38670 49474 38722
rect 49474 38670 49476 38722
rect 49420 38668 49476 38670
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50316 35474 50372 35476
rect 50316 35422 50318 35474
rect 50318 35422 50370 35474
rect 50370 35422 50372 35474
rect 50316 35420 50372 35422
rect 49756 34972 49812 35028
rect 49420 34802 49476 34804
rect 49420 34750 49422 34802
rect 49422 34750 49474 34802
rect 49474 34750 49476 34802
rect 49420 34748 49476 34750
rect 51660 42588 51716 42644
rect 51660 40962 51716 40964
rect 51660 40910 51662 40962
rect 51662 40910 51714 40962
rect 51714 40910 51716 40962
rect 51660 40908 51716 40910
rect 51660 40460 51716 40516
rect 51884 41356 51940 41412
rect 51996 41244 52052 41300
rect 52668 47458 52724 47460
rect 52668 47406 52670 47458
rect 52670 47406 52722 47458
rect 52722 47406 52724 47458
rect 52668 47404 52724 47406
rect 56812 51436 56868 51492
rect 56476 51378 56532 51380
rect 56476 51326 56478 51378
rect 56478 51326 56530 51378
rect 56530 51326 56532 51378
rect 56476 51324 56532 51326
rect 55356 48972 55412 49028
rect 56140 49084 56196 49140
rect 55692 48636 55748 48692
rect 55468 48354 55524 48356
rect 55468 48302 55470 48354
rect 55470 48302 55522 48354
rect 55522 48302 55524 48354
rect 55468 48300 55524 48302
rect 57708 54572 57764 54628
rect 57148 54236 57204 54292
rect 57372 52834 57428 52836
rect 57372 52782 57374 52834
rect 57374 52782 57426 52834
rect 57426 52782 57428 52834
rect 57372 52780 57428 52782
rect 57596 52220 57652 52276
rect 57036 51548 57092 51604
rect 54908 48130 54964 48132
rect 54908 48078 54910 48130
rect 54910 48078 54962 48130
rect 54962 48078 54964 48130
rect 54908 48076 54964 48078
rect 53676 47404 53732 47460
rect 56252 47458 56308 47460
rect 56252 47406 56254 47458
rect 56254 47406 56306 47458
rect 56306 47406 56308 47458
rect 56252 47404 56308 47406
rect 53004 46562 53060 46564
rect 53004 46510 53006 46562
rect 53006 46510 53058 46562
rect 53058 46510 53060 46562
rect 53004 46508 53060 46510
rect 54908 46562 54964 46564
rect 54908 46510 54910 46562
rect 54910 46510 54962 46562
rect 54962 46510 54964 46562
rect 54908 46508 54964 46510
rect 54908 45836 54964 45892
rect 55692 46508 55748 46564
rect 55020 45276 55076 45332
rect 53340 45106 53396 45108
rect 53340 45054 53342 45106
rect 53342 45054 53394 45106
rect 53394 45054 53396 45106
rect 53340 45052 53396 45054
rect 54908 45052 54964 45108
rect 55692 45276 55748 45332
rect 52892 44994 52948 44996
rect 52892 44942 52894 44994
rect 52894 44942 52946 44994
rect 52946 44942 52948 44994
rect 52892 44940 52948 44942
rect 54572 44546 54628 44548
rect 54572 44494 54574 44546
rect 54574 44494 54626 44546
rect 54626 44494 54628 44546
rect 54572 44492 54628 44494
rect 53564 43596 53620 43652
rect 52780 43538 52836 43540
rect 52780 43486 52782 43538
rect 52782 43486 52834 43538
rect 52834 43486 52836 43538
rect 52780 43484 52836 43486
rect 53228 43538 53284 43540
rect 53228 43486 53230 43538
rect 53230 43486 53282 43538
rect 53282 43486 53284 43538
rect 53228 43484 53284 43486
rect 54348 44098 54404 44100
rect 54348 44046 54350 44098
rect 54350 44046 54402 44098
rect 54402 44046 54404 44098
rect 54348 44044 54404 44046
rect 55132 44994 55188 44996
rect 55132 44942 55134 44994
rect 55134 44942 55186 44994
rect 55186 44942 55188 44994
rect 55132 44940 55188 44942
rect 54908 43708 54964 43764
rect 53116 42530 53172 42532
rect 53116 42478 53118 42530
rect 53118 42478 53170 42530
rect 53170 42478 53172 42530
rect 53116 42476 53172 42478
rect 53900 42476 53956 42532
rect 52444 41970 52500 41972
rect 52444 41918 52446 41970
rect 52446 41918 52498 41970
rect 52498 41918 52500 41970
rect 52444 41916 52500 41918
rect 53116 41970 53172 41972
rect 53116 41918 53118 41970
rect 53118 41918 53170 41970
rect 53170 41918 53172 41970
rect 53116 41916 53172 41918
rect 55244 44546 55300 44548
rect 55244 44494 55246 44546
rect 55246 44494 55298 44546
rect 55298 44494 55300 44546
rect 55244 44492 55300 44494
rect 55356 44268 55412 44324
rect 56924 45276 56980 45332
rect 57036 45106 57092 45108
rect 57036 45054 57038 45106
rect 57038 45054 57090 45106
rect 57090 45054 57092 45106
rect 57036 45052 57092 45054
rect 56140 44546 56196 44548
rect 56140 44494 56142 44546
rect 56142 44494 56194 44546
rect 56194 44494 56196 44546
rect 56140 44492 56196 44494
rect 56028 44156 56084 44212
rect 56252 44380 56308 44436
rect 55468 44044 55524 44100
rect 55132 42476 55188 42532
rect 53564 41916 53620 41972
rect 52892 41410 52948 41412
rect 52892 41358 52894 41410
rect 52894 41358 52946 41410
rect 52946 41358 52948 41410
rect 52892 41356 52948 41358
rect 52668 41298 52724 41300
rect 52668 41246 52670 41298
rect 52670 41246 52722 41298
rect 52722 41246 52724 41298
rect 52668 41244 52724 41246
rect 53564 40962 53620 40964
rect 53564 40910 53566 40962
rect 53566 40910 53618 40962
rect 53618 40910 53620 40962
rect 53564 40908 53620 40910
rect 53116 40460 53172 40516
rect 54796 41916 54852 41972
rect 55356 41804 55412 41860
rect 55916 40908 55972 40964
rect 56028 40572 56084 40628
rect 55916 40514 55972 40516
rect 55916 40462 55918 40514
rect 55918 40462 55970 40514
rect 55970 40462 55972 40514
rect 55916 40460 55972 40462
rect 53676 40348 53732 40404
rect 54012 40348 54068 40404
rect 52332 36652 52388 36708
rect 53676 38668 53732 38724
rect 51772 35474 51828 35476
rect 51772 35422 51774 35474
rect 51774 35422 51826 35474
rect 51826 35422 51828 35474
rect 51772 35420 51828 35422
rect 50876 35196 50932 35252
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 53116 35474 53172 35476
rect 53116 35422 53118 35474
rect 53118 35422 53170 35474
rect 53170 35422 53172 35474
rect 53116 35420 53172 35422
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 48972 32562 49028 32564
rect 48972 32510 48974 32562
rect 48974 32510 49026 32562
rect 49026 32510 49028 32562
rect 48972 32508 49028 32510
rect 49644 32562 49700 32564
rect 49644 32510 49646 32562
rect 49646 32510 49698 32562
rect 49698 32510 49700 32562
rect 49644 32508 49700 32510
rect 49308 31778 49364 31780
rect 49308 31726 49310 31778
rect 49310 31726 49362 31778
rect 49362 31726 49364 31778
rect 49308 31724 49364 31726
rect 49420 31666 49476 31668
rect 49420 31614 49422 31666
rect 49422 31614 49474 31666
rect 49474 31614 49476 31666
rect 49420 31612 49476 31614
rect 48972 31500 49028 31556
rect 49532 31500 49588 31556
rect 48748 30156 48804 30212
rect 49084 29596 49140 29652
rect 50428 32562 50484 32564
rect 50428 32510 50430 32562
rect 50430 32510 50482 32562
rect 50482 32510 50484 32562
rect 50428 32508 50484 32510
rect 50092 31836 50148 31892
rect 51436 32060 51492 32116
rect 50876 31836 50932 31892
rect 51884 33346 51940 33348
rect 51884 33294 51886 33346
rect 51886 33294 51938 33346
rect 51938 33294 51940 33346
rect 51884 33292 51940 33294
rect 51996 33234 52052 33236
rect 51996 33182 51998 33234
rect 51998 33182 52050 33234
rect 52050 33182 52052 33234
rect 51996 33180 52052 33182
rect 52220 32620 52276 32676
rect 52668 32620 52724 32676
rect 51772 31836 51828 31892
rect 50428 31724 50484 31780
rect 50204 30770 50260 30772
rect 50204 30718 50206 30770
rect 50206 30718 50258 30770
rect 50258 30718 50260 30770
rect 50204 30716 50260 30718
rect 50764 31554 50820 31556
rect 50764 31502 50766 31554
rect 50766 31502 50818 31554
rect 50818 31502 50820 31554
rect 50764 31500 50820 31502
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50876 30716 50932 30772
rect 49980 30268 50036 30324
rect 49868 30210 49924 30212
rect 49868 30158 49870 30210
rect 49870 30158 49922 30210
rect 49922 30158 49924 30210
rect 49868 30156 49924 30158
rect 51548 30380 51604 30436
rect 50876 30210 50932 30212
rect 50876 30158 50878 30210
rect 50878 30158 50930 30210
rect 50930 30158 50932 30210
rect 50876 30156 50932 30158
rect 52780 32060 52836 32116
rect 53452 34690 53508 34692
rect 53452 34638 53454 34690
rect 53454 34638 53506 34690
rect 53506 34638 53508 34690
rect 53452 34636 53508 34638
rect 53452 33234 53508 33236
rect 53452 33182 53454 33234
rect 53454 33182 53506 33234
rect 53506 33182 53508 33234
rect 53452 33180 53508 33182
rect 53116 31500 53172 31556
rect 51772 30268 51828 30324
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 51100 29650 51156 29652
rect 51100 29598 51102 29650
rect 51102 29598 51154 29650
rect 51154 29598 51156 29650
rect 51100 29596 51156 29598
rect 50988 29426 51044 29428
rect 50988 29374 50990 29426
rect 50990 29374 51042 29426
rect 51042 29374 51044 29426
rect 50988 29372 51044 29374
rect 49644 28812 49700 28868
rect 48524 28754 48580 28756
rect 48524 28702 48526 28754
rect 48526 28702 48578 28754
rect 48578 28702 48580 28754
rect 48524 28700 48580 28702
rect 50652 28812 50708 28868
rect 49756 28754 49812 28756
rect 49756 28702 49758 28754
rect 49758 28702 49810 28754
rect 49810 28702 49812 28754
rect 49756 28700 49812 28702
rect 51548 29538 51604 29540
rect 51548 29486 51550 29538
rect 51550 29486 51602 29538
rect 51602 29486 51604 29538
rect 51548 29484 51604 29486
rect 51436 28700 51492 28756
rect 50092 28418 50148 28420
rect 50092 28366 50094 28418
rect 50094 28366 50146 28418
rect 50146 28366 50148 28418
rect 50092 28364 50148 28366
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50316 27804 50372 27860
rect 47852 26460 47908 26516
rect 46620 25506 46676 25508
rect 46620 25454 46622 25506
rect 46622 25454 46674 25506
rect 46674 25454 46676 25506
rect 46620 25452 46676 25454
rect 47628 26066 47684 26068
rect 47628 26014 47630 26066
rect 47630 26014 47682 26066
rect 47682 26014 47684 26066
rect 47628 26012 47684 26014
rect 47292 25452 47348 25508
rect 46956 25340 47012 25396
rect 45276 24444 45332 24500
rect 44604 23996 44660 24052
rect 45500 23996 45556 24052
rect 49084 26012 49140 26068
rect 52668 30268 52724 30324
rect 51660 28364 51716 28420
rect 53228 29932 53284 29988
rect 53004 29484 53060 29540
rect 53228 29372 53284 29428
rect 52780 27916 52836 27972
rect 53004 28476 53060 28532
rect 51436 27858 51492 27860
rect 51436 27806 51438 27858
rect 51438 27806 51490 27858
rect 51490 27806 51492 27858
rect 51436 27804 51492 27806
rect 52108 26908 52164 26964
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 53564 28530 53620 28532
rect 53564 28478 53566 28530
rect 53566 28478 53618 28530
rect 53618 28478 53620 28530
rect 53564 28476 53620 28478
rect 53340 27804 53396 27860
rect 56028 40236 56084 40292
rect 54124 39058 54180 39060
rect 54124 39006 54126 39058
rect 54126 39006 54178 39058
rect 54178 39006 54180 39058
rect 54124 39004 54180 39006
rect 56588 44322 56644 44324
rect 56588 44270 56590 44322
rect 56590 44270 56642 44322
rect 56642 44270 56644 44322
rect 56588 44268 56644 44270
rect 57596 44380 57652 44436
rect 56700 44210 56756 44212
rect 56700 44158 56702 44210
rect 56702 44158 56754 44210
rect 56754 44158 56756 44210
rect 56700 44156 56756 44158
rect 58044 60562 58100 60564
rect 58044 60510 58046 60562
rect 58046 60510 58098 60562
rect 58098 60510 58100 60562
rect 58044 60508 58100 60510
rect 58044 60002 58100 60004
rect 58044 59950 58046 60002
rect 58046 59950 58098 60002
rect 58098 59950 58100 60002
rect 58044 59948 58100 59950
rect 58156 59218 58212 59220
rect 58156 59166 58158 59218
rect 58158 59166 58210 59218
rect 58210 59166 58212 59218
rect 58156 59164 58212 59166
rect 58156 55298 58212 55300
rect 58156 55246 58158 55298
rect 58158 55246 58210 55298
rect 58210 55246 58212 55298
rect 58156 55244 58212 55246
rect 58156 54236 58212 54292
rect 58156 52780 58212 52836
rect 58156 52220 58212 52276
rect 58156 51548 58212 51604
rect 58156 49138 58212 49140
rect 58156 49086 58158 49138
rect 58158 49086 58210 49138
rect 58210 49086 58212 49138
rect 58156 49084 58212 49086
rect 58044 45890 58100 45892
rect 58044 45838 58046 45890
rect 58046 45838 58098 45890
rect 58098 45838 58100 45890
rect 58044 45836 58100 45838
rect 58156 45330 58212 45332
rect 58156 45278 58158 45330
rect 58158 45278 58210 45330
rect 58210 45278 58212 45330
rect 58156 45276 58212 45278
rect 56700 41858 56756 41860
rect 56700 41806 56702 41858
rect 56702 41806 56754 41858
rect 56754 41806 56756 41858
rect 56700 41804 56756 41806
rect 56700 40514 56756 40516
rect 56700 40462 56702 40514
rect 56702 40462 56754 40514
rect 56754 40462 56756 40514
rect 56700 40460 56756 40462
rect 57036 41804 57092 41860
rect 57260 41132 57316 41188
rect 56588 39564 56644 39620
rect 56924 40348 56980 40404
rect 56364 39452 56420 39508
rect 57036 40236 57092 40292
rect 57036 39618 57092 39620
rect 57036 39566 57038 39618
rect 57038 39566 57090 39618
rect 57090 39566 57092 39618
rect 57036 39564 57092 39566
rect 56812 39506 56868 39508
rect 56812 39454 56814 39506
rect 56814 39454 56866 39506
rect 56866 39454 56868 39506
rect 56812 39452 56868 39454
rect 57708 41132 57764 41188
rect 54908 38050 54964 38052
rect 54908 37998 54910 38050
rect 54910 37998 54962 38050
rect 54962 37998 54964 38050
rect 54908 37996 54964 37998
rect 55356 38050 55412 38052
rect 55356 37998 55358 38050
rect 55358 37998 55410 38050
rect 55410 37998 55412 38050
rect 55356 37996 55412 37998
rect 54012 36988 54068 37044
rect 54012 34636 54068 34692
rect 53788 33292 53844 33348
rect 53900 32786 53956 32788
rect 53900 32734 53902 32786
rect 53902 32734 53954 32786
rect 53954 32734 53956 32786
rect 53900 32732 53956 32734
rect 55580 35532 55636 35588
rect 57596 38722 57652 38724
rect 57596 38670 57598 38722
rect 57598 38670 57650 38722
rect 57650 38670 57652 38722
rect 57596 38668 57652 38670
rect 58156 38668 58212 38724
rect 58156 38556 58212 38612
rect 56700 37996 56756 38052
rect 54908 32732 54964 32788
rect 55020 34188 55076 34244
rect 56924 35868 56980 35924
rect 55804 34636 55860 34692
rect 56252 34802 56308 34804
rect 56252 34750 56254 34802
rect 56254 34750 56306 34802
rect 56306 34750 56308 34802
rect 56252 34748 56308 34750
rect 57708 35922 57764 35924
rect 57708 35870 57710 35922
rect 57710 35870 57762 35922
rect 57762 35870 57764 35922
rect 57708 35868 57764 35870
rect 57036 35698 57092 35700
rect 57036 35646 57038 35698
rect 57038 35646 57090 35698
rect 57090 35646 57092 35698
rect 57036 35644 57092 35646
rect 57148 35532 57204 35588
rect 57036 34802 57092 34804
rect 57036 34750 57038 34802
rect 57038 34750 57090 34802
rect 57090 34750 57092 34802
rect 57036 34748 57092 34750
rect 56252 34188 56308 34244
rect 55020 33292 55076 33348
rect 54796 32674 54852 32676
rect 54796 32622 54798 32674
rect 54798 32622 54850 32674
rect 54850 32622 54852 32674
rect 54796 32620 54852 32622
rect 55244 32060 55300 32116
rect 55132 30380 55188 30436
rect 54572 29986 54628 29988
rect 54572 29934 54574 29986
rect 54574 29934 54626 29986
rect 54626 29934 54628 29986
rect 54572 29932 54628 29934
rect 54908 29986 54964 29988
rect 54908 29934 54910 29986
rect 54910 29934 54962 29986
rect 54962 29934 54964 29986
rect 54908 29932 54964 29934
rect 53900 28588 53956 28644
rect 54236 28642 54292 28644
rect 54236 28590 54238 28642
rect 54238 28590 54290 28642
rect 54290 28590 54292 28642
rect 54236 28588 54292 28590
rect 55356 30940 55412 30996
rect 55132 28476 55188 28532
rect 55356 28700 55412 28756
rect 53452 27692 53508 27748
rect 52780 26962 52836 26964
rect 52780 26910 52782 26962
rect 52782 26910 52834 26962
rect 52834 26910 52836 26962
rect 52780 26908 52836 26910
rect 50204 25228 50260 25284
rect 48300 24556 48356 24612
rect 48748 24556 48804 24612
rect 44940 23548 44996 23604
rect 45388 23548 45444 23604
rect 45052 23324 45108 23380
rect 44940 23266 44996 23268
rect 44940 23214 44942 23266
rect 44942 23214 44994 23266
rect 44994 23214 44996 23266
rect 44940 23212 44996 23214
rect 45836 23436 45892 23492
rect 45612 23212 45668 23268
rect 45612 22370 45668 22372
rect 45612 22318 45614 22370
rect 45614 22318 45666 22370
rect 45666 22318 45668 22370
rect 45612 22316 45668 22318
rect 45388 22204 45444 22260
rect 44492 18450 44548 18452
rect 44492 18398 44494 18450
rect 44494 18398 44546 18450
rect 44546 18398 44548 18450
rect 44492 18396 44548 18398
rect 44604 19964 44660 20020
rect 45276 19964 45332 20020
rect 44604 19292 44660 19348
rect 43932 18172 43988 18228
rect 44268 17836 44324 17892
rect 44268 17388 44324 17444
rect 43708 13634 43764 13636
rect 43708 13582 43710 13634
rect 43710 13582 43762 13634
rect 43762 13582 43764 13634
rect 43708 13580 43764 13582
rect 44044 14476 44100 14532
rect 43708 12962 43764 12964
rect 43708 12910 43710 12962
rect 43710 12910 43762 12962
rect 43762 12910 43764 12962
rect 43708 12908 43764 12910
rect 43484 12348 43540 12404
rect 44156 13356 44212 13412
rect 43036 11506 43092 11508
rect 43036 11454 43038 11506
rect 43038 11454 43090 11506
rect 43090 11454 43092 11506
rect 43036 11452 43092 11454
rect 43148 10610 43204 10612
rect 43148 10558 43150 10610
rect 43150 10558 43202 10610
rect 43202 10558 43204 10610
rect 43148 10556 43204 10558
rect 42588 9938 42644 9940
rect 42588 9886 42590 9938
rect 42590 9886 42642 9938
rect 42642 9886 42644 9938
rect 42588 9884 42644 9886
rect 43036 10108 43092 10164
rect 42476 9660 42532 9716
rect 44044 12572 44100 12628
rect 45724 22428 45780 22484
rect 44716 18956 44772 19012
rect 45276 18620 45332 18676
rect 44716 18508 44772 18564
rect 46508 22988 46564 23044
rect 46844 23436 46900 23492
rect 46732 22370 46788 22372
rect 46732 22318 46734 22370
rect 46734 22318 46786 22370
rect 46786 22318 46788 22370
rect 46732 22316 46788 22318
rect 45948 22204 46004 22260
rect 46396 22092 46452 22148
rect 46284 19964 46340 20020
rect 46172 19404 46228 19460
rect 45948 18620 46004 18676
rect 45724 18060 45780 18116
rect 44940 17666 44996 17668
rect 44940 17614 44942 17666
rect 44942 17614 44994 17666
rect 44994 17614 44996 17666
rect 44940 17612 44996 17614
rect 45276 17836 45332 17892
rect 45052 15820 45108 15876
rect 45388 15874 45444 15876
rect 45388 15822 45390 15874
rect 45390 15822 45442 15874
rect 45442 15822 45444 15874
rect 45388 15820 45444 15822
rect 45724 15874 45780 15876
rect 45724 15822 45726 15874
rect 45726 15822 45778 15874
rect 45778 15822 45780 15874
rect 45724 15820 45780 15822
rect 45724 15260 45780 15316
rect 44716 15202 44772 15204
rect 44716 15150 44718 15202
rect 44718 15150 44770 15202
rect 44770 15150 44772 15202
rect 44716 15148 44772 15150
rect 44716 14530 44772 14532
rect 44716 14478 44718 14530
rect 44718 14478 44770 14530
rect 44770 14478 44772 14530
rect 44716 14476 44772 14478
rect 44940 13858 44996 13860
rect 44940 13806 44942 13858
rect 44942 13806 44994 13858
rect 44994 13806 44996 13858
rect 44940 13804 44996 13806
rect 44604 13468 44660 13524
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 52220 24668 52276 24724
rect 52332 25340 52388 25396
rect 52780 25282 52836 25284
rect 52780 25230 52782 25282
rect 52782 25230 52834 25282
rect 52834 25230 52836 25282
rect 52780 25228 52836 25230
rect 55580 32732 55636 32788
rect 56028 32060 56084 32116
rect 57260 34636 57316 34692
rect 57932 35698 57988 35700
rect 57932 35646 57934 35698
rect 57934 35646 57986 35698
rect 57986 35646 57988 35698
rect 57932 35644 57988 35646
rect 57596 34636 57652 34692
rect 57036 33122 57092 33124
rect 57036 33070 57038 33122
rect 57038 33070 57090 33122
rect 57090 33070 57092 33122
rect 57036 33068 57092 33070
rect 56588 30994 56644 30996
rect 56588 30942 56590 30994
rect 56590 30942 56642 30994
rect 56642 30942 56644 30994
rect 56588 30940 56644 30942
rect 56924 30940 56980 30996
rect 57484 33346 57540 33348
rect 57484 33294 57486 33346
rect 57486 33294 57538 33346
rect 57538 33294 57540 33346
rect 57484 33292 57540 33294
rect 57596 33122 57652 33124
rect 57596 33070 57598 33122
rect 57598 33070 57650 33122
rect 57650 33070 57652 33122
rect 57596 33068 57652 33070
rect 58156 32060 58212 32116
rect 58156 31388 58212 31444
rect 57820 31106 57876 31108
rect 57820 31054 57822 31106
rect 57822 31054 57874 31106
rect 57874 31054 57876 31106
rect 57820 31052 57876 31054
rect 57036 29932 57092 29988
rect 56924 29650 56980 29652
rect 56924 29598 56926 29650
rect 56926 29598 56978 29650
rect 56978 29598 56980 29650
rect 56924 29596 56980 29598
rect 57484 29932 57540 29988
rect 57372 29596 57428 29652
rect 56588 28754 56644 28756
rect 56588 28702 56590 28754
rect 56590 28702 56642 28754
rect 56642 28702 56644 28754
rect 56588 28700 56644 28702
rect 55468 28140 55524 28196
rect 56588 28476 56644 28532
rect 53676 27804 53732 27860
rect 55132 27858 55188 27860
rect 55132 27806 55134 27858
rect 55134 27806 55186 27858
rect 55186 27806 55188 27858
rect 55132 27804 55188 27806
rect 54236 27746 54292 27748
rect 54236 27694 54238 27746
rect 54238 27694 54290 27746
rect 54290 27694 54292 27746
rect 54236 27692 54292 27694
rect 53676 26850 53732 26852
rect 53676 26798 53678 26850
rect 53678 26798 53730 26850
rect 53730 26798 53732 26850
rect 53676 26796 53732 26798
rect 54236 26908 54292 26964
rect 55020 27244 55076 27300
rect 53676 25394 53732 25396
rect 53676 25342 53678 25394
rect 53678 25342 53730 25394
rect 53730 25342 53732 25394
rect 53676 25340 53732 25342
rect 52892 24722 52948 24724
rect 52892 24670 52894 24722
rect 52894 24670 52946 24722
rect 52946 24670 52948 24722
rect 52892 24668 52948 24670
rect 52780 23996 52836 24052
rect 52892 23826 52948 23828
rect 52892 23774 52894 23826
rect 52894 23774 52946 23826
rect 52946 23774 52948 23826
rect 52892 23772 52948 23774
rect 51436 23660 51492 23716
rect 48748 23324 48804 23380
rect 47964 23100 48020 23156
rect 46956 21756 47012 21812
rect 47180 22092 47236 22148
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 53004 23714 53060 23716
rect 53004 23662 53006 23714
rect 53006 23662 53058 23714
rect 53058 23662 53060 23714
rect 53004 23660 53060 23662
rect 53228 23938 53284 23940
rect 53228 23886 53230 23938
rect 53230 23886 53282 23938
rect 53282 23886 53284 23938
rect 53228 23884 53284 23886
rect 52220 23212 52276 23268
rect 50428 23100 50484 23156
rect 48188 23042 48244 23044
rect 48188 22990 48190 23042
rect 48190 22990 48242 23042
rect 48242 22990 48244 23042
rect 48188 22988 48244 22990
rect 50764 22988 50820 23044
rect 51212 22988 51268 23044
rect 48188 22428 48244 22484
rect 50204 22428 50260 22484
rect 49084 21868 49140 21924
rect 46844 20018 46900 20020
rect 46844 19966 46846 20018
rect 46846 19966 46898 20018
rect 46898 19966 46900 20018
rect 46844 19964 46900 19966
rect 46732 19906 46788 19908
rect 46732 19854 46734 19906
rect 46734 19854 46786 19906
rect 46786 19854 46788 19906
rect 46732 19852 46788 19854
rect 46956 19740 47012 19796
rect 46732 18508 46788 18564
rect 46620 17442 46676 17444
rect 46620 17390 46622 17442
rect 46622 17390 46674 17442
rect 46674 17390 46676 17442
rect 46620 17388 46676 17390
rect 45500 12850 45556 12852
rect 45500 12798 45502 12850
rect 45502 12798 45554 12850
rect 45554 12798 45556 12850
rect 45500 12796 45556 12798
rect 45276 12572 45332 12628
rect 44716 12290 44772 12292
rect 44716 12238 44718 12290
rect 44718 12238 44770 12290
rect 44770 12238 44772 12290
rect 44716 12236 44772 12238
rect 45612 12236 45668 12292
rect 43820 9826 43876 9828
rect 43820 9774 43822 9826
rect 43822 9774 43874 9826
rect 43874 9774 43876 9826
rect 43820 9772 43876 9774
rect 42812 9154 42868 9156
rect 42812 9102 42814 9154
rect 42814 9102 42866 9154
rect 42866 9102 42868 9154
rect 42812 9100 42868 9102
rect 42140 8204 42196 8260
rect 41468 7868 41524 7924
rect 43596 9212 43652 9268
rect 42924 8092 42980 8148
rect 40012 7698 40068 7700
rect 40012 7646 40014 7698
rect 40014 7646 40066 7698
rect 40066 7646 40068 7698
rect 40012 7644 40068 7646
rect 40124 7586 40180 7588
rect 40124 7534 40126 7586
rect 40126 7534 40178 7586
rect 40178 7534 40180 7586
rect 40124 7532 40180 7534
rect 39900 7420 39956 7476
rect 39676 7196 39732 7252
rect 40236 6690 40292 6692
rect 40236 6638 40238 6690
rect 40238 6638 40290 6690
rect 40290 6638 40292 6690
rect 40236 6636 40292 6638
rect 40012 6300 40068 6356
rect 40796 7474 40852 7476
rect 40796 7422 40798 7474
rect 40798 7422 40850 7474
rect 40850 7422 40852 7474
rect 40796 7420 40852 7422
rect 40796 6914 40852 6916
rect 40796 6862 40798 6914
rect 40798 6862 40850 6914
rect 40850 6862 40852 6914
rect 40796 6860 40852 6862
rect 41468 7698 41524 7700
rect 41468 7646 41470 7698
rect 41470 7646 41522 7698
rect 41522 7646 41524 7698
rect 41468 7644 41524 7646
rect 41244 7474 41300 7476
rect 41244 7422 41246 7474
rect 41246 7422 41298 7474
rect 41298 7422 41300 7474
rect 41244 7420 41300 7422
rect 41692 7532 41748 7588
rect 41244 6802 41300 6804
rect 41244 6750 41246 6802
rect 41246 6750 41298 6802
rect 41298 6750 41300 6802
rect 41244 6748 41300 6750
rect 40572 6636 40628 6692
rect 40348 6300 40404 6356
rect 39452 5292 39508 5348
rect 39900 5292 39956 5348
rect 38220 5068 38276 5124
rect 39116 5122 39172 5124
rect 39116 5070 39118 5122
rect 39118 5070 39170 5122
rect 39170 5070 39172 5122
rect 39116 5068 39172 5070
rect 40908 5292 40964 5348
rect 40796 4396 40852 4452
rect 41804 7420 41860 7476
rect 43484 9154 43540 9156
rect 43484 9102 43486 9154
rect 43486 9102 43538 9154
rect 43538 9102 43540 9154
rect 43484 9100 43540 9102
rect 43708 7980 43764 8036
rect 43820 7586 43876 7588
rect 43820 7534 43822 7586
rect 43822 7534 43874 7586
rect 43874 7534 43876 7586
rect 43820 7532 43876 7534
rect 43260 7084 43316 7140
rect 43260 6748 43316 6804
rect 43036 6636 43092 6692
rect 44268 10556 44324 10612
rect 41804 6524 41860 6580
rect 43820 6412 43876 6468
rect 41244 5292 41300 5348
rect 41692 4450 41748 4452
rect 41692 4398 41694 4450
rect 41694 4398 41746 4450
rect 41746 4398 41748 4450
rect 41692 4396 41748 4398
rect 43932 6188 43988 6244
rect 44940 8370 44996 8372
rect 44940 8318 44942 8370
rect 44942 8318 44994 8370
rect 44994 8318 44996 8370
rect 44940 8316 44996 8318
rect 45612 8316 45668 8372
rect 45724 8204 45780 8260
rect 46396 8258 46452 8260
rect 46396 8206 46398 8258
rect 46398 8206 46450 8258
rect 46450 8206 46452 8258
rect 46396 8204 46452 8206
rect 46172 8034 46228 8036
rect 46172 7982 46174 8034
rect 46174 7982 46226 8034
rect 46226 7982 46228 8034
rect 46172 7980 46228 7982
rect 45164 6636 45220 6692
rect 45052 6076 45108 6132
rect 46620 15202 46676 15204
rect 46620 15150 46622 15202
rect 46622 15150 46674 15202
rect 46674 15150 46676 15202
rect 46620 15148 46676 15150
rect 47292 19964 47348 20020
rect 47180 19234 47236 19236
rect 47180 19182 47182 19234
rect 47182 19182 47234 19234
rect 47234 19182 47236 19234
rect 47180 19180 47236 19182
rect 47180 17666 47236 17668
rect 47180 17614 47182 17666
rect 47182 17614 47234 17666
rect 47234 17614 47236 17666
rect 47180 17612 47236 17614
rect 47516 19740 47572 19796
rect 47628 19404 47684 19460
rect 47964 19964 48020 20020
rect 47852 19852 47908 19908
rect 47740 19068 47796 19124
rect 47852 18060 47908 18116
rect 47404 17442 47460 17444
rect 47404 17390 47406 17442
rect 47406 17390 47458 17442
rect 47458 17390 47460 17442
rect 47404 17388 47460 17390
rect 47740 15932 47796 15988
rect 47180 15820 47236 15876
rect 46844 15314 46900 15316
rect 46844 15262 46846 15314
rect 46846 15262 46898 15314
rect 46898 15262 46900 15314
rect 46844 15260 46900 15262
rect 47292 15484 47348 15540
rect 48972 15820 49028 15876
rect 48972 15484 49028 15540
rect 49644 21810 49700 21812
rect 49644 21758 49646 21810
rect 49646 21758 49698 21810
rect 49698 21758 49700 21810
rect 49644 21756 49700 21758
rect 49756 21698 49812 21700
rect 49756 21646 49758 21698
rect 49758 21646 49810 21698
rect 49810 21646 49812 21698
rect 49756 21644 49812 21646
rect 50092 19180 50148 19236
rect 49868 17612 49924 17668
rect 49308 17500 49364 17556
rect 49420 15820 49476 15876
rect 47628 14252 47684 14308
rect 48076 14530 48132 14532
rect 48076 14478 48078 14530
rect 48078 14478 48130 14530
rect 48130 14478 48132 14530
rect 48076 14476 48132 14478
rect 48300 14364 48356 14420
rect 47516 13804 47572 13860
rect 47292 13746 47348 13748
rect 47292 13694 47294 13746
rect 47294 13694 47346 13746
rect 47346 13694 47348 13746
rect 47292 13692 47348 13694
rect 47516 12850 47572 12852
rect 47516 12798 47518 12850
rect 47518 12798 47570 12850
rect 47570 12798 47572 12850
rect 47516 12796 47572 12798
rect 47852 12572 47908 12628
rect 47852 11452 47908 11508
rect 46620 10668 46676 10724
rect 46620 8146 46676 8148
rect 46620 8094 46622 8146
rect 46622 8094 46674 8146
rect 46674 8094 46676 8146
rect 46620 8092 46676 8094
rect 49308 14700 49364 14756
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50988 21644 51044 21700
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50092 15820 50148 15876
rect 50876 19122 50932 19124
rect 50876 19070 50878 19122
rect 50878 19070 50930 19122
rect 50930 19070 50932 19122
rect 50876 19068 50932 19070
rect 50764 19010 50820 19012
rect 50764 18958 50766 19010
rect 50766 18958 50818 19010
rect 50818 18958 50820 19010
rect 50764 18956 50820 18958
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 51212 18956 51268 19012
rect 51100 18508 51156 18564
rect 50652 17948 50708 18004
rect 50988 17724 51044 17780
rect 50652 17666 50708 17668
rect 50652 17614 50654 17666
rect 50654 17614 50706 17666
rect 50706 17614 50708 17666
rect 50652 17612 50708 17614
rect 50428 17500 50484 17556
rect 51324 18172 51380 18228
rect 51548 18396 51604 18452
rect 51436 17948 51492 18004
rect 51100 17388 51156 17444
rect 51884 19010 51940 19012
rect 51884 18958 51886 19010
rect 51886 18958 51938 19010
rect 51938 18958 51940 19010
rect 51884 18956 51940 18958
rect 52220 18450 52276 18452
rect 52220 18398 52222 18450
rect 52222 18398 52274 18450
rect 52274 18398 52276 18450
rect 52220 18396 52276 18398
rect 52556 18284 52612 18340
rect 51772 18172 51828 18228
rect 51324 17388 51380 17444
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 51436 16882 51492 16884
rect 51436 16830 51438 16882
rect 51438 16830 51490 16882
rect 51490 16830 51492 16882
rect 51436 16828 51492 16830
rect 51660 16828 51716 16884
rect 50540 15986 50596 15988
rect 50540 15934 50542 15986
rect 50542 15934 50594 15986
rect 50594 15934 50596 15986
rect 50540 15932 50596 15934
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50204 15202 50260 15204
rect 50204 15150 50206 15202
rect 50206 15150 50258 15202
rect 50258 15150 50260 15202
rect 50204 15148 50260 15150
rect 49532 13244 49588 13300
rect 49868 12348 49924 12404
rect 50652 15036 50708 15092
rect 52332 18226 52388 18228
rect 52332 18174 52334 18226
rect 52334 18174 52386 18226
rect 52386 18174 52388 18226
rect 52332 18172 52388 18174
rect 52108 17836 52164 17892
rect 51996 17052 52052 17108
rect 51772 16716 51828 16772
rect 52332 17388 52388 17444
rect 52780 17890 52836 17892
rect 52780 17838 52782 17890
rect 52782 17838 52834 17890
rect 52834 17838 52836 17890
rect 52780 17836 52836 17838
rect 52332 16716 52388 16772
rect 51772 15372 51828 15428
rect 51548 15202 51604 15204
rect 51548 15150 51550 15202
rect 51550 15150 51602 15202
rect 51602 15150 51604 15202
rect 51548 15148 51604 15150
rect 51100 14924 51156 14980
rect 51996 14924 52052 14980
rect 52108 15484 52164 15540
rect 50540 14754 50596 14756
rect 50540 14702 50542 14754
rect 50542 14702 50594 14754
rect 50594 14702 50596 14754
rect 50540 14700 50596 14702
rect 50428 14588 50484 14644
rect 50204 14530 50260 14532
rect 50204 14478 50206 14530
rect 50206 14478 50258 14530
rect 50258 14478 50260 14530
rect 50204 14476 50260 14478
rect 51212 14700 51268 14756
rect 50764 14642 50820 14644
rect 50764 14590 50766 14642
rect 50766 14590 50818 14642
rect 50818 14590 50820 14642
rect 50764 14588 50820 14590
rect 50540 14252 50596 14308
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 51212 14530 51268 14532
rect 51212 14478 51214 14530
rect 51214 14478 51266 14530
rect 51266 14478 51268 14530
rect 51212 14476 51268 14478
rect 51772 14418 51828 14420
rect 51772 14366 51774 14418
rect 51774 14366 51826 14418
rect 51826 14366 51828 14418
rect 51772 14364 51828 14366
rect 50988 14252 51044 14308
rect 50204 13746 50260 13748
rect 50204 13694 50206 13746
rect 50206 13694 50258 13746
rect 50258 13694 50260 13746
rect 50204 13692 50260 13694
rect 51548 14306 51604 14308
rect 51548 14254 51550 14306
rect 51550 14254 51602 14306
rect 51602 14254 51604 14306
rect 51548 14252 51604 14254
rect 50316 13580 50372 13636
rect 50092 11676 50148 11732
rect 48860 11506 48916 11508
rect 48860 11454 48862 11506
rect 48862 11454 48914 11506
rect 48914 11454 48916 11506
rect 48860 11452 48916 11454
rect 50204 12796 50260 12852
rect 48300 10668 48356 10724
rect 50876 13468 50932 13524
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50316 12236 50372 12292
rect 50652 12402 50708 12404
rect 50652 12350 50654 12402
rect 50654 12350 50706 12402
rect 50706 12350 50708 12402
rect 50652 12348 50708 12350
rect 50764 11788 50820 11844
rect 51436 12348 51492 12404
rect 51884 13692 51940 13748
rect 52220 13580 52276 13636
rect 52556 17388 52612 17444
rect 52892 17500 52948 17556
rect 53452 23996 53508 24052
rect 53452 23826 53508 23828
rect 53452 23774 53454 23826
rect 53454 23774 53506 23826
rect 53506 23774 53508 23826
rect 53452 23772 53508 23774
rect 53340 22988 53396 23044
rect 54124 24668 54180 24724
rect 54460 23938 54516 23940
rect 54460 23886 54462 23938
rect 54462 23886 54514 23938
rect 54514 23886 54516 23938
rect 54460 23884 54516 23886
rect 54124 23266 54180 23268
rect 54124 23214 54126 23266
rect 54126 23214 54178 23266
rect 54178 23214 54180 23266
rect 54124 23212 54180 23214
rect 54684 23042 54740 23044
rect 54684 22990 54686 23042
rect 54686 22990 54738 23042
rect 54738 22990 54740 23042
rect 54684 22988 54740 22990
rect 54572 22258 54628 22260
rect 54572 22206 54574 22258
rect 54574 22206 54626 22258
rect 54626 22206 54628 22258
rect 54572 22204 54628 22206
rect 54796 21532 54852 21588
rect 53452 18396 53508 18452
rect 53228 18338 53284 18340
rect 53228 18286 53230 18338
rect 53230 18286 53282 18338
rect 53282 18286 53284 18338
rect 53228 18284 53284 18286
rect 53116 17948 53172 18004
rect 54460 18338 54516 18340
rect 54460 18286 54462 18338
rect 54462 18286 54514 18338
rect 54514 18286 54516 18338
rect 54460 18284 54516 18286
rect 53564 18172 53620 18228
rect 53788 18060 53844 18116
rect 54572 18226 54628 18228
rect 54572 18174 54574 18226
rect 54574 18174 54626 18226
rect 54626 18174 54628 18226
rect 54572 18172 54628 18174
rect 54124 17836 54180 17892
rect 53228 17500 53284 17556
rect 53116 17442 53172 17444
rect 53116 17390 53118 17442
rect 53118 17390 53170 17442
rect 53170 17390 53172 17442
rect 53116 17388 53172 17390
rect 52668 17052 52724 17108
rect 52892 16882 52948 16884
rect 52892 16830 52894 16882
rect 52894 16830 52946 16882
rect 52946 16830 52948 16882
rect 52892 16828 52948 16830
rect 52444 15372 52500 15428
rect 52668 15148 52724 15204
rect 52780 14754 52836 14756
rect 52780 14702 52782 14754
rect 52782 14702 52834 14754
rect 52834 14702 52836 14754
rect 52780 14700 52836 14702
rect 52780 13858 52836 13860
rect 52780 13806 52782 13858
rect 52782 13806 52834 13858
rect 52834 13806 52836 13858
rect 52780 13804 52836 13806
rect 52668 13746 52724 13748
rect 52668 13694 52670 13746
rect 52670 13694 52722 13746
rect 52722 13694 52724 13746
rect 52668 13692 52724 13694
rect 52220 12290 52276 12292
rect 52220 12238 52222 12290
rect 52222 12238 52274 12290
rect 52274 12238 52276 12290
rect 52220 12236 52276 12238
rect 50988 11788 51044 11844
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 46844 10108 46900 10164
rect 49868 10610 49924 10612
rect 49868 10558 49870 10610
rect 49870 10558 49922 10610
rect 49922 10558 49924 10610
rect 49868 10556 49924 10558
rect 47180 9100 47236 9156
rect 47404 8370 47460 8372
rect 47404 8318 47406 8370
rect 47406 8318 47458 8370
rect 47458 8318 47460 8370
rect 47404 8316 47460 8318
rect 47516 8258 47572 8260
rect 47516 8206 47518 8258
rect 47518 8206 47570 8258
rect 47570 8206 47572 8258
rect 47516 8204 47572 8206
rect 47852 8146 47908 8148
rect 47852 8094 47854 8146
rect 47854 8094 47906 8146
rect 47906 8094 47908 8146
rect 47852 8092 47908 8094
rect 47180 7980 47236 8036
rect 47180 7756 47236 7812
rect 46508 6636 46564 6692
rect 47292 6636 47348 6692
rect 46620 6300 46676 6356
rect 46732 6130 46788 6132
rect 46732 6078 46734 6130
rect 46734 6078 46786 6130
rect 46786 6078 46788 6130
rect 46732 6076 46788 6078
rect 44604 5180 44660 5236
rect 44940 5628 44996 5684
rect 45276 5628 45332 5684
rect 45500 5234 45556 5236
rect 45500 5182 45502 5234
rect 45502 5182 45554 5234
rect 45554 5182 45556 5234
rect 45500 5180 45556 5182
rect 46508 6018 46564 6020
rect 46508 5966 46510 6018
rect 46510 5966 46562 6018
rect 46562 5966 46564 6018
rect 46508 5964 46564 5966
rect 46508 5180 46564 5236
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 47068 6018 47124 6020
rect 47068 5966 47070 6018
rect 47070 5966 47122 6018
rect 47122 5966 47124 6018
rect 47068 5964 47124 5966
rect 48188 6412 48244 6468
rect 48860 8258 48916 8260
rect 48860 8206 48862 8258
rect 48862 8206 48914 8258
rect 48914 8206 48916 8258
rect 48860 8204 48916 8206
rect 48636 8092 48692 8148
rect 48524 7980 48580 8036
rect 49308 7868 49364 7924
rect 48636 7308 48692 7364
rect 50876 10668 50932 10724
rect 51660 11506 51716 11508
rect 51660 11454 51662 11506
rect 51662 11454 51714 11506
rect 51714 11454 51716 11506
rect 51660 11452 51716 11454
rect 52668 12290 52724 12292
rect 52668 12238 52670 12290
rect 52670 12238 52722 12290
rect 52722 12238 52724 12290
rect 52668 12236 52724 12238
rect 52108 11394 52164 11396
rect 52108 11342 52110 11394
rect 52110 11342 52162 11394
rect 52162 11342 52164 11394
rect 52108 11340 52164 11342
rect 53452 17164 53508 17220
rect 53564 17276 53620 17332
rect 54348 17612 54404 17668
rect 55468 27970 55524 27972
rect 55468 27918 55470 27970
rect 55470 27918 55522 27970
rect 55522 27918 55524 27970
rect 55468 27916 55524 27918
rect 57260 27970 57316 27972
rect 57260 27918 57262 27970
rect 57262 27918 57314 27970
rect 57314 27918 57316 27970
rect 57260 27916 57316 27918
rect 58156 29596 58212 29652
rect 58044 28700 58100 28756
rect 57932 27970 57988 27972
rect 57932 27918 57934 27970
rect 57934 27918 57986 27970
rect 57986 27918 57988 27970
rect 57932 27916 57988 27918
rect 56812 27692 56868 27748
rect 56028 26460 56084 26516
rect 56700 27132 56756 27188
rect 56924 27580 56980 27636
rect 57036 26514 57092 26516
rect 57036 26462 57038 26514
rect 57038 26462 57090 26514
rect 57090 26462 57092 26514
rect 57036 26460 57092 26462
rect 57932 27634 57988 27636
rect 57932 27582 57934 27634
rect 57934 27582 57986 27634
rect 57986 27582 57988 27634
rect 57932 27580 57988 27582
rect 56588 24668 56644 24724
rect 57596 25282 57652 25284
rect 57596 25230 57598 25282
rect 57598 25230 57650 25282
rect 57650 25230 57652 25282
rect 57596 25228 57652 25230
rect 55132 23324 55188 23380
rect 56700 23378 56756 23380
rect 56700 23326 56702 23378
rect 56702 23326 56754 23378
rect 56754 23326 56756 23378
rect 56700 23324 56756 23326
rect 56588 23266 56644 23268
rect 56588 23214 56590 23266
rect 56590 23214 56642 23266
rect 56642 23214 56644 23266
rect 56588 23212 56644 23214
rect 57148 24722 57204 24724
rect 57148 24670 57150 24722
rect 57150 24670 57202 24722
rect 57202 24670 57204 24722
rect 57148 24668 57204 24670
rect 56812 22370 56868 22372
rect 56812 22318 56814 22370
rect 56814 22318 56866 22370
rect 56866 22318 56868 22370
rect 56812 22316 56868 22318
rect 57036 22258 57092 22260
rect 57036 22206 57038 22258
rect 57038 22206 57090 22258
rect 57090 22206 57092 22258
rect 57036 22204 57092 22206
rect 55132 21980 55188 22036
rect 55132 21586 55188 21588
rect 55132 21534 55134 21586
rect 55134 21534 55186 21586
rect 55186 21534 55188 21586
rect 55132 21532 55188 21534
rect 56924 22092 56980 22148
rect 57484 24610 57540 24612
rect 57484 24558 57486 24610
rect 57486 24558 57538 24610
rect 57538 24558 57540 24610
rect 57484 24556 57540 24558
rect 57932 23212 57988 23268
rect 57372 22370 57428 22372
rect 57372 22318 57374 22370
rect 57374 22318 57426 22370
rect 57426 22318 57428 22370
rect 57372 22316 57428 22318
rect 58156 27916 58212 27972
rect 58156 27186 58212 27188
rect 58156 27134 58158 27186
rect 58158 27134 58210 27186
rect 58210 27134 58212 27186
rect 58156 27132 58212 27134
rect 58268 25564 58324 25620
rect 58156 25228 58212 25284
rect 58156 24444 58212 24500
rect 57148 21980 57204 22036
rect 57596 22146 57652 22148
rect 57596 22094 57598 22146
rect 57598 22094 57650 22146
rect 57650 22094 57652 22146
rect 57596 22092 57652 22094
rect 55020 17500 55076 17556
rect 55132 17164 55188 17220
rect 53788 16828 53844 16884
rect 53340 16770 53396 16772
rect 53340 16718 53342 16770
rect 53342 16718 53394 16770
rect 53394 16718 53396 16770
rect 53340 16716 53396 16718
rect 55132 16828 55188 16884
rect 53564 15036 53620 15092
rect 56476 18172 56532 18228
rect 57820 17554 57876 17556
rect 57820 17502 57822 17554
rect 57822 17502 57874 17554
rect 57874 17502 57876 17554
rect 57820 17500 57876 17502
rect 58156 17554 58212 17556
rect 58156 17502 58158 17554
rect 58158 17502 58210 17554
rect 58210 17502 58212 17554
rect 58156 17500 58212 17502
rect 55244 16716 55300 16772
rect 57036 16940 57092 16996
rect 54012 15036 54068 15092
rect 54460 15036 54516 15092
rect 53340 14418 53396 14420
rect 53340 14366 53342 14418
rect 53342 14366 53394 14418
rect 53394 14366 53396 14418
rect 53340 14364 53396 14366
rect 54124 14418 54180 14420
rect 54124 14366 54126 14418
rect 54126 14366 54178 14418
rect 54178 14366 54180 14418
rect 54124 14364 54180 14366
rect 56588 14418 56644 14420
rect 56588 14366 56590 14418
rect 56590 14366 56642 14418
rect 56642 14366 56644 14418
rect 56588 14364 56644 14366
rect 53116 14306 53172 14308
rect 53116 14254 53118 14306
rect 53118 14254 53170 14306
rect 53170 14254 53172 14306
rect 53116 14252 53172 14254
rect 55244 13858 55300 13860
rect 55244 13806 55246 13858
rect 55246 13806 55298 13858
rect 55298 13806 55300 13858
rect 55244 13804 55300 13806
rect 53116 13634 53172 13636
rect 53116 13582 53118 13634
rect 53118 13582 53170 13634
rect 53170 13582 53172 13634
rect 53116 13580 53172 13582
rect 54460 13580 54516 13636
rect 53004 12738 53060 12740
rect 53004 12686 53006 12738
rect 53006 12686 53058 12738
rect 53058 12686 53060 12738
rect 53004 12684 53060 12686
rect 55916 13580 55972 13636
rect 56700 13634 56756 13636
rect 56700 13582 56702 13634
rect 56702 13582 56754 13634
rect 56754 13582 56756 13634
rect 56700 13580 56756 13582
rect 54460 11676 54516 11732
rect 55580 11676 55636 11732
rect 57372 16716 57428 16772
rect 57260 14364 57316 14420
rect 57820 14418 57876 14420
rect 57820 14366 57822 14418
rect 57822 14366 57874 14418
rect 57874 14366 57876 14418
rect 57820 14364 57876 14366
rect 57260 13580 57316 13636
rect 54796 11506 54852 11508
rect 54796 11454 54798 11506
rect 54798 11454 54850 11506
rect 54850 11454 54852 11506
rect 54796 11452 54852 11454
rect 52892 11340 52948 11396
rect 51324 10722 51380 10724
rect 51324 10670 51326 10722
rect 51326 10670 51378 10722
rect 51378 10670 51380 10722
rect 51324 10668 51380 10670
rect 51212 10556 51268 10612
rect 50652 10498 50708 10500
rect 50652 10446 50654 10498
rect 50654 10446 50706 10498
rect 50706 10446 50708 10498
rect 50652 10444 50708 10446
rect 50204 9996 50260 10052
rect 50988 9996 51044 10052
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 49980 9154 50036 9156
rect 49980 9102 49982 9154
rect 49982 9102 50034 9154
rect 50034 9102 50036 9154
rect 49980 9100 50036 9102
rect 49868 8146 49924 8148
rect 49868 8094 49870 8146
rect 49870 8094 49922 8146
rect 49922 8094 49924 8146
rect 49868 8092 49924 8094
rect 49532 7980 49588 8036
rect 49420 7196 49476 7252
rect 48412 6076 48468 6132
rect 47068 5122 47124 5124
rect 47068 5070 47070 5122
rect 47070 5070 47122 5122
rect 47122 5070 47124 5122
rect 47068 5068 47124 5070
rect 46956 4508 47012 4564
rect 46060 4172 46116 4228
rect 47068 4226 47124 4228
rect 47068 4174 47070 4226
rect 47070 4174 47122 4226
rect 47122 4174 47124 4226
rect 47068 4172 47124 4174
rect 48748 6802 48804 6804
rect 48748 6750 48750 6802
rect 48750 6750 48802 6802
rect 48802 6750 48804 6802
rect 48748 6748 48804 6750
rect 49868 7474 49924 7476
rect 49868 7422 49870 7474
rect 49870 7422 49922 7474
rect 49922 7422 49924 7474
rect 49868 7420 49924 7422
rect 50428 8428 50484 8484
rect 50428 8258 50484 8260
rect 50428 8206 50430 8258
rect 50430 8206 50482 8258
rect 50482 8206 50484 8258
rect 50428 8204 50484 8206
rect 51548 9884 51604 9940
rect 51324 9266 51380 9268
rect 51324 9214 51326 9266
rect 51326 9214 51378 9266
rect 51378 9214 51380 9266
rect 51324 9212 51380 9214
rect 52444 10722 52500 10724
rect 52444 10670 52446 10722
rect 52446 10670 52498 10722
rect 52498 10670 52500 10722
rect 52444 10668 52500 10670
rect 51996 10332 52052 10388
rect 52668 9938 52724 9940
rect 52668 9886 52670 9938
rect 52670 9886 52722 9938
rect 52722 9886 52724 9938
rect 52668 9884 52724 9886
rect 51660 9714 51716 9716
rect 51660 9662 51662 9714
rect 51662 9662 51714 9714
rect 51714 9662 51716 9714
rect 51660 9660 51716 9662
rect 54796 9714 54852 9716
rect 54796 9662 54798 9714
rect 54798 9662 54850 9714
rect 54850 9662 54852 9714
rect 54796 9660 54852 9662
rect 58156 10610 58212 10612
rect 58156 10558 58158 10610
rect 58158 10558 58210 10610
rect 58210 10558 58212 10610
rect 58156 10556 58212 10558
rect 51996 9212 52052 9268
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50652 7532 50708 7588
rect 50652 7196 50708 7252
rect 50876 7308 50932 7364
rect 49980 6802 50036 6804
rect 49980 6750 49982 6802
rect 49982 6750 50034 6802
rect 50034 6750 50036 6802
rect 49980 6748 50036 6750
rect 49756 6690 49812 6692
rect 49756 6638 49758 6690
rect 49758 6638 49810 6690
rect 49810 6638 49812 6690
rect 49756 6636 49812 6638
rect 49420 6578 49476 6580
rect 49420 6526 49422 6578
rect 49422 6526 49474 6578
rect 49474 6526 49476 6578
rect 49420 6524 49476 6526
rect 50428 6524 50484 6580
rect 51212 8370 51268 8372
rect 51212 8318 51214 8370
rect 51214 8318 51266 8370
rect 51266 8318 51268 8370
rect 51212 8316 51268 8318
rect 51324 8204 51380 8260
rect 51548 7532 51604 7588
rect 51436 7474 51492 7476
rect 51436 7422 51438 7474
rect 51438 7422 51490 7474
rect 51490 7422 51492 7474
rect 51436 7420 51492 7422
rect 51548 7362 51604 7364
rect 51548 7310 51550 7362
rect 51550 7310 51602 7362
rect 51602 7310 51604 7362
rect 51548 7308 51604 7310
rect 52444 7362 52500 7364
rect 52444 7310 52446 7362
rect 52446 7310 52498 7362
rect 52498 7310 52500 7362
rect 52444 7308 52500 7310
rect 51548 6748 51604 6804
rect 52668 6802 52724 6804
rect 52668 6750 52670 6802
rect 52670 6750 52722 6802
rect 52722 6750 52724 6802
rect 52668 6748 52724 6750
rect 52556 6636 52612 6692
rect 54796 6690 54852 6692
rect 54796 6638 54798 6690
rect 54798 6638 54850 6690
rect 54850 6638 54852 6690
rect 54796 6636 54852 6638
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50428 6076 50484 6132
rect 49868 5852 49924 5908
rect 48860 5180 48916 5236
rect 48748 4562 48804 4564
rect 48748 4510 48750 4562
rect 48750 4510 48802 4562
rect 48802 4510 48804 4562
rect 48748 4508 48804 4510
rect 49868 5234 49924 5236
rect 49868 5182 49870 5234
rect 49870 5182 49922 5234
rect 49922 5182 49924 5234
rect 49868 5180 49924 5182
rect 50316 5122 50372 5124
rect 50316 5070 50318 5122
rect 50318 5070 50370 5122
rect 50370 5070 50372 5122
rect 50316 5068 50372 5070
rect 48524 4172 48580 4228
rect 51212 6076 51268 6132
rect 54012 6412 54068 6468
rect 53340 4956 53396 5012
rect 51324 4898 51380 4900
rect 51324 4846 51326 4898
rect 51326 4846 51378 4898
rect 51378 4846 51380 4898
rect 51324 4844 51380 4846
rect 52668 4844 52724 4900
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 55468 4956 55524 5012
rect 54012 4284 54068 4340
rect 57596 4338 57652 4340
rect 57596 4286 57598 4338
rect 57598 4286 57650 4338
rect 57650 4286 57652 4338
rect 57596 4284 57652 4286
rect 57372 4226 57428 4228
rect 57372 4174 57374 4226
rect 57374 4174 57426 4226
rect 57426 4174 57428 4226
rect 57372 4172 57428 4174
rect 58156 4172 58212 4228
rect 58156 3612 58212 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 4722 66780 4732 66836
rect 4788 66780 5516 66836
rect 5572 66780 5582 66836
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 24882 66444 24892 66500
rect 24948 66444 26124 66500
rect 26180 66444 26190 66500
rect 38994 66444 39004 66500
rect 39060 66444 40796 66500
rect 40852 66444 40862 66500
rect 45042 66444 45052 66500
rect 45108 66444 48412 66500
rect 48468 66444 48478 66500
rect 49074 66444 49084 66500
rect 49140 66444 52220 66500
rect 52276 66444 52286 66500
rect 53106 66444 53116 66500
rect 53172 66444 56028 66500
rect 56084 66444 56094 66500
rect 59200 66164 60000 66192
rect 43026 66108 43036 66164
rect 43092 66108 46172 66164
rect 46228 66108 46238 66164
rect 58146 66108 58156 66164
rect 58212 66108 60000 66164
rect 59200 66080 60000 66108
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 51090 65548 51100 65604
rect 51156 65548 51166 65604
rect 51100 65492 51156 65548
rect 20178 65436 20188 65492
rect 20244 65436 20860 65492
rect 20916 65436 20926 65492
rect 33842 65436 33852 65492
rect 33908 65436 34860 65492
rect 34916 65436 35532 65492
rect 35588 65436 35598 65492
rect 41010 65436 41020 65492
rect 41076 65436 42700 65492
rect 42756 65436 42766 65492
rect 51100 65436 52332 65492
rect 52388 65436 52398 65492
rect 55010 65436 55020 65492
rect 55076 65436 57148 65492
rect 57204 65436 57214 65492
rect 57586 65436 57596 65492
rect 57652 65436 58156 65492
rect 58212 65436 58222 65492
rect 17602 65324 17612 65380
rect 17668 65324 19516 65380
rect 19572 65324 19582 65380
rect 34962 65324 34972 65380
rect 35028 65324 35644 65380
rect 35700 65324 35710 65380
rect 38546 65324 38556 65380
rect 38612 65324 41132 65380
rect 41188 65324 42028 65380
rect 42084 65324 44380 65380
rect 44436 65324 44446 65380
rect 46498 65324 46508 65380
rect 46564 65324 47740 65380
rect 47796 65324 47806 65380
rect 51762 65324 51772 65380
rect 51828 65324 54124 65380
rect 54180 65324 54190 65380
rect 54898 65324 54908 65380
rect 54964 65324 55356 65380
rect 37426 65212 37436 65268
rect 37492 65212 40124 65268
rect 40180 65212 40190 65268
rect 55412 65212 55468 65380
rect 55524 65212 55534 65268
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 22530 64876 22540 64932
rect 22596 64876 23548 64932
rect 23604 64876 23614 64932
rect 30258 64876 30268 64932
rect 30324 64876 55244 64932
rect 55300 64876 55310 64932
rect 5730 64652 5740 64708
rect 5796 64652 8876 64708
rect 8932 64652 9324 64708
rect 9380 64652 12572 64708
rect 12628 64652 12638 64708
rect 17938 64652 17948 64708
rect 18004 64652 20188 64708
rect 20244 64652 20254 64708
rect 27794 64652 27804 64708
rect 27860 64652 29148 64708
rect 29204 64652 29484 64708
rect 29540 64652 30380 64708
rect 30436 64652 30446 64708
rect 36642 64652 36652 64708
rect 36708 64652 37100 64708
rect 37156 64652 38556 64708
rect 38612 64652 38622 64708
rect 11778 64540 11788 64596
rect 11844 64540 12684 64596
rect 12740 64540 13804 64596
rect 13860 64540 13870 64596
rect 30930 64540 30940 64596
rect 30996 64540 32956 64596
rect 33012 64540 33022 64596
rect 12226 64428 12236 64484
rect 12292 64428 12796 64484
rect 12852 64428 13468 64484
rect 13524 64428 13534 64484
rect 20850 64428 20860 64484
rect 20916 64428 21420 64484
rect 21476 64428 21868 64484
rect 21924 64428 23212 64484
rect 23268 64428 23996 64484
rect 24052 64428 25452 64484
rect 25508 64428 25518 64484
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 26674 64204 26684 64260
rect 26740 64204 27468 64260
rect 27524 64204 28140 64260
rect 28196 64204 28206 64260
rect 11442 63980 11452 64036
rect 11508 63980 12124 64036
rect 12180 63980 12190 64036
rect 16706 63980 16716 64036
rect 16772 63980 17724 64036
rect 17780 63980 17790 64036
rect 32284 63924 32340 64540
rect 33282 64428 33292 64484
rect 33348 64428 34636 64484
rect 34692 64428 34702 64484
rect 52098 64428 52108 64484
rect 52164 64428 52780 64484
rect 52836 64428 54012 64484
rect 54068 64428 54908 64484
rect 54964 64428 55356 64484
rect 55412 64428 58044 64484
rect 58100 64428 58110 64484
rect 43652 64316 47516 64372
rect 47572 64316 47582 64372
rect 43652 64148 43708 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 44930 64204 44940 64260
rect 44996 64204 49532 64260
rect 49588 64204 49598 64260
rect 39218 64092 39228 64148
rect 39284 64092 41580 64148
rect 41636 64092 43708 64148
rect 45602 64092 45612 64148
rect 45668 64092 46508 64148
rect 46564 64092 46574 64148
rect 46722 64092 46732 64148
rect 46788 64092 54572 64148
rect 54628 64092 54638 64148
rect 44818 63980 44828 64036
rect 44884 63980 46844 64036
rect 46900 63980 46910 64036
rect 55010 63980 55020 64036
rect 55076 63980 55244 64036
rect 55300 63980 55310 64036
rect 12562 63868 12572 63924
rect 12628 63868 13580 63924
rect 13636 63868 16828 63924
rect 16884 63868 16894 63924
rect 23650 63868 23660 63924
rect 23716 63868 26852 63924
rect 32274 63868 32284 63924
rect 32340 63868 32350 63924
rect 32498 63868 32508 63924
rect 32564 63868 33180 63924
rect 33236 63868 33246 63924
rect 43362 63868 43372 63924
rect 43428 63868 43820 63924
rect 43876 63868 43886 63924
rect 45154 63868 45164 63924
rect 45220 63868 46396 63924
rect 46452 63868 46462 63924
rect 49522 63868 49532 63924
rect 49588 63868 51324 63924
rect 51380 63868 51390 63924
rect 26796 63812 26852 63868
rect 26796 63756 31724 63812
rect 31780 63756 31790 63812
rect 54674 63756 54684 63812
rect 54740 63756 54750 63812
rect 55122 63756 55132 63812
rect 55188 63756 56364 63812
rect 56420 63756 56430 63812
rect 26338 63644 26348 63700
rect 26404 63644 27244 63700
rect 27300 63644 28252 63700
rect 28308 63644 28318 63700
rect 54684 63588 54740 63756
rect 55010 63644 55020 63700
rect 55076 63644 56588 63700
rect 56644 63644 56654 63700
rect 31938 63532 31948 63588
rect 32004 63532 32844 63588
rect 32900 63532 32910 63588
rect 47730 63532 47740 63588
rect 47796 63532 50652 63588
rect 50708 63532 54460 63588
rect 54516 63532 54526 63588
rect 54684 63532 55804 63588
rect 55860 63532 56700 63588
rect 56756 63532 56766 63588
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 9986 63308 9996 63364
rect 10052 63308 12348 63364
rect 12404 63308 12414 63364
rect 21074 63308 21084 63364
rect 21140 63308 22316 63364
rect 22372 63308 22382 63364
rect 31266 63308 31276 63364
rect 31332 63308 31948 63364
rect 32004 63308 33068 63364
rect 33124 63308 33134 63364
rect 24770 63196 24780 63252
rect 24836 63196 26236 63252
rect 26292 63196 26302 63252
rect 49970 63196 49980 63252
rect 50036 63196 51100 63252
rect 51156 63196 51166 63252
rect 52994 63196 53004 63252
rect 53060 63196 53900 63252
rect 53956 63196 55244 63252
rect 55300 63196 55310 63252
rect 13906 63084 13916 63140
rect 13972 63084 15484 63140
rect 15540 63084 17276 63140
rect 17332 63084 17342 63140
rect 26674 63084 26684 63140
rect 26740 63084 27132 63140
rect 27188 63084 27198 63140
rect 30146 63084 30156 63140
rect 30212 63084 30940 63140
rect 30996 63084 31276 63140
rect 31332 63084 31342 63140
rect 43474 63084 43484 63140
rect 43540 63084 44044 63140
rect 44100 63084 44940 63140
rect 44996 63084 45006 63140
rect 46050 63084 46060 63140
rect 46116 63084 47292 63140
rect 47348 63084 47740 63140
rect 47796 63084 47806 63140
rect 49074 63084 49084 63140
rect 49140 63084 49644 63140
rect 49700 63084 50764 63140
rect 50820 63084 50830 63140
rect 6514 62972 6524 63028
rect 6580 62972 7308 63028
rect 7364 62972 7644 63028
rect 7700 62972 7710 63028
rect 16370 62972 16380 63028
rect 16436 62972 17612 63028
rect 17668 62972 17678 63028
rect 26450 62972 26460 63028
rect 26516 62972 27244 63028
rect 27300 62972 27310 63028
rect 41010 62972 41020 63028
rect 41076 62972 41804 63028
rect 41860 62972 44156 63028
rect 44212 62972 45052 63028
rect 45108 62972 45118 63028
rect 12450 62860 12460 62916
rect 12516 62860 13692 62916
rect 13748 62860 13758 62916
rect 16258 62860 16268 62916
rect 16324 62860 17388 62916
rect 17444 62860 17454 62916
rect 17826 62860 17836 62916
rect 17892 62860 18508 62916
rect 18564 62860 22092 62916
rect 22148 62860 22158 62916
rect 26114 62860 26124 62916
rect 26180 62860 27020 62916
rect 27076 62860 27086 62916
rect 27570 62860 27580 62916
rect 27636 62860 28476 62916
rect 28532 62860 28542 62916
rect 28914 62860 28924 62916
rect 28980 62860 29484 62916
rect 29540 62860 29550 62916
rect 41906 62860 41916 62916
rect 41972 62860 42924 62916
rect 42980 62860 42990 62916
rect 43652 62860 45276 62916
rect 45332 62860 47180 62916
rect 47236 62860 47246 62916
rect 43652 62804 43708 62860
rect 37874 62748 37884 62804
rect 37940 62748 43708 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 45602 62524 45612 62580
rect 45668 62524 46508 62580
rect 46564 62524 46574 62580
rect 48850 62524 48860 62580
rect 48916 62524 52108 62580
rect 52164 62524 52174 62580
rect 7084 62412 8540 62468
rect 8596 62412 8606 62468
rect 10882 62412 10892 62468
rect 10948 62412 18956 62468
rect 19012 62412 19022 62468
rect 37426 62412 37436 62468
rect 37492 62412 38220 62468
rect 38276 62412 38286 62468
rect 39442 62412 39452 62468
rect 39508 62412 52444 62468
rect 52500 62412 53228 62468
rect 53284 62412 53294 62468
rect 7084 62356 7140 62412
rect 6738 62300 6748 62356
rect 6804 62300 7084 62356
rect 7140 62300 7150 62356
rect 8082 62300 8092 62356
rect 8148 62300 10220 62356
rect 10276 62300 10286 62356
rect 13682 62300 13692 62356
rect 13748 62300 15148 62356
rect 15204 62300 15214 62356
rect 18162 62300 18172 62356
rect 18228 62300 19516 62356
rect 19572 62300 19582 62356
rect 27234 62300 27244 62356
rect 27300 62300 28364 62356
rect 28420 62300 29484 62356
rect 29540 62300 29550 62356
rect 35858 62300 35868 62356
rect 35924 62300 41244 62356
rect 41300 62300 41310 62356
rect 42690 62300 42700 62356
rect 42756 62300 43484 62356
rect 43540 62300 43550 62356
rect 43652 62300 43932 62356
rect 43988 62300 43998 62356
rect 44930 62300 44940 62356
rect 44996 62300 45724 62356
rect 45780 62300 45790 62356
rect 7858 62188 7868 62244
rect 7924 62188 10556 62244
rect 10612 62188 10622 62244
rect 20402 62188 20412 62244
rect 20468 62188 20860 62244
rect 20916 62188 32956 62244
rect 33012 62188 33022 62244
rect 36754 62188 36764 62244
rect 36820 62188 41020 62244
rect 41076 62188 42252 62244
rect 42308 62188 42318 62244
rect 43586 62188 43596 62244
rect 43652 62188 43708 62300
rect 50082 62188 50092 62244
rect 50148 62188 51660 62244
rect 51716 62188 51726 62244
rect 52882 62188 52892 62244
rect 52948 62188 54124 62244
rect 54180 62188 54190 62244
rect 25890 62076 25900 62132
rect 25956 62076 27692 62132
rect 27748 62076 27758 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 48850 61852 48860 61908
rect 48916 61852 50988 61908
rect 51044 61852 51054 61908
rect 54124 61572 54180 62188
rect 54124 61516 55468 61572
rect 55524 61516 55534 61572
rect 42018 61404 42028 61460
rect 42084 61404 43708 61460
rect 43764 61404 44156 61460
rect 44212 61404 44222 61460
rect 6178 61292 6188 61348
rect 6244 61292 6860 61348
rect 6916 61292 6926 61348
rect 22642 61292 22652 61348
rect 22708 61292 25564 61348
rect 25620 61292 31052 61348
rect 31108 61292 31118 61348
rect 32386 61292 32396 61348
rect 32452 61292 37772 61348
rect 37828 61292 37838 61348
rect 38322 61292 38332 61348
rect 38388 61292 39900 61348
rect 39956 61292 39966 61348
rect 28130 61180 28140 61236
rect 28196 61180 34524 61236
rect 34580 61180 35196 61236
rect 35252 61180 36092 61236
rect 36148 61180 36158 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 25106 61068 25116 61124
rect 25172 61068 26908 61124
rect 29586 61068 29596 61124
rect 29652 61068 34412 61124
rect 34468 61068 34972 61124
rect 35028 61068 35868 61124
rect 35924 61068 35934 61124
rect 37884 61068 38668 61124
rect 38724 61068 38734 61124
rect 54450 61068 54460 61124
rect 54516 61068 55244 61124
rect 55300 61068 57372 61124
rect 57428 61068 57932 61124
rect 57988 61068 57998 61124
rect 26852 61012 26908 61068
rect 37884 61012 37940 61068
rect 25442 60956 25452 61012
rect 25508 60956 26012 61012
rect 26068 60956 26078 61012
rect 26852 60956 37324 61012
rect 37380 60956 37884 61012
rect 37940 60956 37950 61012
rect 49046 60956 49084 61012
rect 49140 60956 49150 61012
rect 49746 60956 49756 61012
rect 49812 60956 50428 61012
rect 50484 60956 50988 61012
rect 51044 60956 51436 61012
rect 51492 60956 51502 61012
rect 49084 60900 49140 60956
rect 10994 60844 11004 60900
rect 11060 60844 13244 60900
rect 13300 60844 13310 60900
rect 16258 60844 16268 60900
rect 16324 60844 17500 60900
rect 17556 60844 17566 60900
rect 27794 60844 27804 60900
rect 27860 60844 33852 60900
rect 33908 60844 34748 60900
rect 34804 60844 34814 60900
rect 35410 60844 35420 60900
rect 35476 60844 37548 60900
rect 37604 60844 37614 60900
rect 37762 60844 37772 60900
rect 37828 60844 39116 60900
rect 39172 60844 39182 60900
rect 49084 60844 50204 60900
rect 50260 60844 50270 60900
rect 56914 60844 56924 60900
rect 56980 60844 57372 60900
rect 57428 60844 57438 60900
rect 10210 60732 10220 60788
rect 10276 60732 10780 60788
rect 10836 60732 13356 60788
rect 13412 60732 13422 60788
rect 14578 60732 14588 60788
rect 14644 60732 22652 60788
rect 22708 60732 22718 60788
rect 25442 60732 25452 60788
rect 25508 60732 25900 60788
rect 25956 60732 27132 60788
rect 27188 60732 27198 60788
rect 27906 60732 27916 60788
rect 27972 60732 28924 60788
rect 28980 60732 28990 60788
rect 40002 60732 40012 60788
rect 40068 60732 51660 60788
rect 51716 60732 53004 60788
rect 53060 60732 53070 60788
rect 53330 60732 53340 60788
rect 53396 60732 54684 60788
rect 54740 60732 57708 60788
rect 57764 60732 57774 60788
rect 5618 60620 5628 60676
rect 5684 60620 6300 60676
rect 6356 60620 6366 60676
rect 21746 60620 21756 60676
rect 21812 60620 23212 60676
rect 23268 60620 23548 60676
rect 23604 60620 25676 60676
rect 25732 60620 25742 60676
rect 26852 60620 27692 60676
rect 27748 60620 28700 60676
rect 28756 60620 28766 60676
rect 30034 60620 30044 60676
rect 30100 60620 30492 60676
rect 30548 60620 30828 60676
rect 30884 60620 31276 60676
rect 31332 60620 31342 60676
rect 40450 60620 40460 60676
rect 40516 60620 41916 60676
rect 41972 60620 44940 60676
rect 44996 60620 45006 60676
rect 49522 60620 49532 60676
rect 49588 60620 49756 60676
rect 49812 60620 49822 60676
rect 50978 60620 50988 60676
rect 51044 60620 52780 60676
rect 52836 60620 52846 60676
rect 26852 60564 26908 60620
rect 15698 60508 15708 60564
rect 15764 60508 26908 60564
rect 27234 60508 27244 60564
rect 27300 60508 28028 60564
rect 28084 60508 29932 60564
rect 29988 60508 29998 60564
rect 32050 60508 32060 60564
rect 32116 60508 33292 60564
rect 33348 60508 33358 60564
rect 34738 60508 34748 60564
rect 34804 60508 36988 60564
rect 37044 60508 37054 60564
rect 39890 60508 39900 60564
rect 39956 60508 41468 60564
rect 41524 60508 41804 60564
rect 41860 60508 42476 60564
rect 42532 60508 42542 60564
rect 56914 60508 56924 60564
rect 56980 60508 58044 60564
rect 58100 60508 58110 60564
rect 18834 60396 18844 60452
rect 18900 60396 20188 60452
rect 20244 60396 20254 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 20132 60284 33180 60340
rect 33236 60284 33404 60340
rect 33460 60284 33470 60340
rect 20132 60228 20188 60284
rect 10546 60172 10556 60228
rect 10612 60172 12964 60228
rect 17602 60172 17612 60228
rect 17668 60172 20188 60228
rect 28354 60172 28364 60228
rect 28420 60172 29260 60228
rect 29316 60172 29326 60228
rect 44258 60172 44268 60228
rect 44324 60172 48860 60228
rect 48916 60172 48926 60228
rect 51202 60172 51212 60228
rect 51268 60172 51884 60228
rect 51940 60172 51950 60228
rect 9090 60060 9100 60116
rect 9156 60060 11788 60116
rect 11844 60060 11854 60116
rect 12908 60004 12964 60172
rect 15586 60060 15596 60116
rect 15652 60060 38108 60116
rect 38164 60060 38174 60116
rect 8418 59948 8428 60004
rect 8484 59948 8652 60004
rect 8708 59948 11340 60004
rect 11396 59948 11406 60004
rect 12898 59948 12908 60004
rect 12964 59948 15148 60004
rect 15204 59948 15214 60004
rect 27458 59948 27468 60004
rect 27524 59948 29372 60004
rect 29428 59948 29438 60004
rect 31154 59948 31164 60004
rect 31220 59948 33628 60004
rect 33684 59948 33694 60004
rect 52098 59948 52108 60004
rect 52164 59948 53340 60004
rect 53396 59948 54236 60004
rect 54292 59948 54302 60004
rect 54898 59948 54908 60004
rect 54964 59948 58044 60004
rect 58100 59948 58110 60004
rect 16146 59836 16156 59892
rect 16212 59836 18060 59892
rect 18116 59836 18126 59892
rect 23986 59836 23996 59892
rect 24052 59836 26572 59892
rect 26628 59836 26638 59892
rect 30370 59836 30380 59892
rect 30436 59836 32396 59892
rect 32452 59836 32462 59892
rect 12450 59724 12460 59780
rect 12516 59724 14028 59780
rect 14084 59724 14094 59780
rect 16706 59724 16716 59780
rect 16772 59724 18172 59780
rect 18228 59724 19852 59780
rect 19908 59724 19918 59780
rect 31042 59724 31052 59780
rect 31108 59724 40012 59780
rect 40068 59724 41692 59780
rect 41748 59724 41758 59780
rect 39442 59612 39452 59668
rect 39508 59612 41916 59668
rect 41972 59612 42812 59668
rect 42868 59612 44156 59668
rect 44212 59612 44222 59668
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 24658 59500 24668 59556
rect 24724 59500 30380 59556
rect 30436 59500 30446 59556
rect 40674 59500 40684 59556
rect 40740 59500 40750 59556
rect 3490 59388 3500 59444
rect 3556 59388 7644 59444
rect 7700 59388 7710 59444
rect 15026 59388 15036 59444
rect 15092 59388 17164 59444
rect 17220 59388 17230 59444
rect 7522 59276 7532 59332
rect 7588 59276 8204 59332
rect 8260 59276 8428 59332
rect 11330 59276 11340 59332
rect 11396 59276 12796 59332
rect 12852 59276 12862 59332
rect 17602 59276 17612 59332
rect 17668 59276 18060 59332
rect 18116 59276 18126 59332
rect 8372 58996 8428 59276
rect 40684 59220 40740 59500
rect 47058 59388 47068 59444
rect 47124 59388 48300 59444
rect 48356 59388 50428 59444
rect 50484 59388 51436 59444
rect 51492 59388 54684 59444
rect 54740 59388 54750 59444
rect 55412 59388 56028 59444
rect 56084 59388 56924 59444
rect 56980 59388 56990 59444
rect 55412 59332 55468 59388
rect 42354 59276 42364 59332
rect 42420 59276 43036 59332
rect 43092 59276 43102 59332
rect 48178 59276 48188 59332
rect 48244 59276 49532 59332
rect 49588 59276 49598 59332
rect 50372 59276 55468 59332
rect 34850 59164 34860 59220
rect 34916 59164 37100 59220
rect 37156 59164 37166 59220
rect 40684 59164 41244 59220
rect 41300 59164 43260 59220
rect 43316 59164 43326 59220
rect 43810 59164 43820 59220
rect 43876 59164 45276 59220
rect 45332 59164 45342 59220
rect 18050 59052 18060 59108
rect 18116 59052 25116 59108
rect 25172 59052 25182 59108
rect 31378 59052 31388 59108
rect 31444 59052 32284 59108
rect 32340 59052 32350 59108
rect 39218 59052 39228 59108
rect 39284 59052 41020 59108
rect 41076 59052 41086 59108
rect 8372 58940 20300 58996
rect 20356 58940 21084 58996
rect 21140 58940 21150 58996
rect 40338 58940 40348 58996
rect 40404 58940 40796 58996
rect 40852 58940 40862 58996
rect 50372 58884 50428 59276
rect 59200 59220 60000 59248
rect 58146 59164 58156 59220
rect 58212 59164 60000 59220
rect 59200 59136 60000 59164
rect 12786 58828 12796 58884
rect 12852 58828 16212 58884
rect 45714 58828 45724 58884
rect 45780 58828 49868 58884
rect 49924 58828 50428 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 16156 58772 16212 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 4834 58716 4844 58772
rect 4900 58716 5852 58772
rect 5908 58716 6636 58772
rect 6692 58716 6702 58772
rect 12226 58716 12236 58772
rect 12292 58716 14588 58772
rect 14644 58716 14654 58772
rect 16146 58716 16156 58772
rect 16212 58716 16222 58772
rect 43250 58716 43260 58772
rect 43316 58716 48860 58772
rect 48916 58716 48926 58772
rect 4844 58660 4900 58716
rect 1810 58604 1820 58660
rect 1876 58604 2828 58660
rect 2884 58604 4900 58660
rect 37762 58492 37772 58548
rect 37828 58492 38556 58548
rect 38612 58492 41020 58548
rect 41076 58492 41804 58548
rect 41860 58492 42364 58548
rect 42420 58492 42430 58548
rect 45266 58492 45276 58548
rect 45332 58492 46956 58548
rect 47012 58492 47022 58548
rect 25666 58380 25676 58436
rect 25732 58380 26684 58436
rect 26740 58380 26750 58436
rect 43138 58380 43148 58436
rect 43204 58380 44828 58436
rect 44884 58380 44894 58436
rect 0 58324 800 58352
rect 0 58268 1708 58324
rect 1764 58268 1774 58324
rect 3826 58268 3836 58324
rect 3892 58268 4060 58324
rect 4116 58268 4956 58324
rect 5012 58268 5022 58324
rect 10994 58268 11004 58324
rect 11060 58268 11788 58324
rect 11844 58268 11854 58324
rect 20738 58268 20748 58324
rect 20804 58268 26012 58324
rect 26068 58268 26078 58324
rect 29810 58268 29820 58324
rect 29876 58268 30492 58324
rect 30548 58268 30558 58324
rect 41682 58268 41692 58324
rect 41748 58268 52556 58324
rect 52612 58268 53004 58324
rect 53060 58268 53070 58324
rect 0 58240 800 58268
rect 2482 58156 2492 58212
rect 2548 58156 3948 58212
rect 4004 58156 4014 58212
rect 15362 58156 15372 58212
rect 15428 58156 16156 58212
rect 16212 58156 16492 58212
rect 16548 58156 26236 58212
rect 26292 58156 26302 58212
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 19730 57820 19740 57876
rect 19796 57820 20300 57876
rect 20356 57820 24668 57876
rect 24724 57820 24734 57876
rect 13794 57708 13804 57764
rect 13860 57708 14924 57764
rect 14980 57708 16604 57764
rect 16660 57708 16670 57764
rect 27682 57708 27692 57764
rect 27748 57708 35532 57764
rect 35588 57708 36204 57764
rect 36260 57708 37660 57764
rect 37716 57708 37726 57764
rect 8418 57596 8428 57652
rect 8484 57596 9436 57652
rect 9492 57596 9502 57652
rect 10098 57596 10108 57652
rect 10164 57596 10668 57652
rect 10724 57596 10734 57652
rect 13346 57596 13356 57652
rect 13412 57596 13916 57652
rect 13972 57596 13982 57652
rect 19394 57596 19404 57652
rect 19460 57596 20300 57652
rect 20356 57596 20366 57652
rect 20738 57596 20748 57652
rect 20804 57596 20814 57652
rect 26852 57596 28252 57652
rect 28308 57596 28318 57652
rect 30146 57596 30156 57652
rect 30212 57596 30940 57652
rect 30996 57596 31006 57652
rect 32386 57596 32396 57652
rect 32452 57596 33180 57652
rect 33236 57596 33740 57652
rect 33796 57596 33806 57652
rect 43586 57596 43596 57652
rect 43652 57596 44492 57652
rect 44548 57596 44558 57652
rect 51426 57596 51436 57652
rect 51492 57596 51502 57652
rect 20748 57540 20804 57596
rect 4610 57484 4620 57540
rect 4676 57484 5628 57540
rect 5684 57484 5694 57540
rect 19058 57484 19068 57540
rect 19124 57484 20804 57540
rect 26852 57428 26908 57596
rect 51436 57540 51492 57596
rect 42578 57484 42588 57540
rect 42644 57484 43148 57540
rect 43204 57484 43214 57540
rect 51090 57484 51100 57540
rect 51156 57484 51492 57540
rect 17948 57372 26460 57428
rect 26516 57372 26908 57428
rect 34962 57372 34972 57428
rect 35028 57372 37772 57428
rect 37828 57372 37838 57428
rect 47058 57372 47068 57428
rect 47124 57372 48188 57428
rect 48244 57372 49420 57428
rect 49476 57372 49486 57428
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 17948 57092 18004 57372
rect 30034 57260 30044 57316
rect 30100 57260 30604 57316
rect 30660 57260 31612 57316
rect 31668 57260 31678 57316
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 5842 57036 5852 57092
rect 5908 57036 6188 57092
rect 6244 57036 6254 57092
rect 9986 57036 9996 57092
rect 10052 57036 10444 57092
rect 10500 57036 10510 57092
rect 10770 57036 10780 57092
rect 10836 57036 12236 57092
rect 12292 57036 12302 57092
rect 16034 57036 16044 57092
rect 16100 57036 18004 57092
rect 25666 57036 25676 57092
rect 25732 57036 26740 57092
rect 32274 57036 32284 57092
rect 32340 57036 36876 57092
rect 36932 57036 36942 57092
rect 4834 56924 4844 56980
rect 4900 56924 5516 56980
rect 5572 56924 5582 56980
rect 26684 56868 26740 57036
rect 32386 56924 32396 56980
rect 32452 56924 33740 56980
rect 33796 56924 33806 56980
rect 5282 56812 5292 56868
rect 5348 56812 6748 56868
rect 6804 56812 8652 56868
rect 8708 56812 9772 56868
rect 9828 56812 9838 56868
rect 19842 56812 19852 56868
rect 19908 56812 20748 56868
rect 20804 56812 20814 56868
rect 26674 56812 26684 56868
rect 26740 56812 27692 56868
rect 27748 56812 27758 56868
rect 36418 56812 36428 56868
rect 36484 56812 37100 56868
rect 37156 56812 37166 56868
rect 37986 56812 37996 56868
rect 38052 56812 42252 56868
rect 42308 56812 42318 56868
rect 6850 56700 6860 56756
rect 6916 56700 8428 56756
rect 8754 56700 8764 56756
rect 8820 56700 9884 56756
rect 9940 56700 9950 56756
rect 13682 56700 13692 56756
rect 13748 56700 14252 56756
rect 14308 56700 15148 56756
rect 15204 56700 15214 56756
rect 35186 56700 35196 56756
rect 35252 56700 36092 56756
rect 36148 56700 37324 56756
rect 37380 56700 38220 56756
rect 38276 56700 38286 56756
rect 42914 56700 42924 56756
rect 42980 56700 43260 56756
rect 43316 56700 43326 56756
rect 8372 56644 8428 56700
rect 8372 56588 11228 56644
rect 11284 56588 12012 56644
rect 12068 56588 12078 56644
rect 12562 56588 12572 56644
rect 12628 56588 13916 56644
rect 13972 56588 14700 56644
rect 14756 56588 14766 56644
rect 51986 56476 51996 56532
rect 52052 56476 52780 56532
rect 52836 56476 52846 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 8194 56252 8204 56308
rect 8260 56252 8764 56308
rect 8820 56252 8830 56308
rect 47618 56252 47628 56308
rect 47684 56252 47964 56308
rect 48020 56252 49980 56308
rect 50036 56252 50046 56308
rect 50306 56252 50316 56308
rect 50372 56252 50876 56308
rect 50932 56252 50942 56308
rect 8306 56140 8316 56196
rect 8372 56140 9212 56196
rect 9268 56140 9278 56196
rect 13346 56140 13356 56196
rect 13412 56140 14028 56196
rect 14084 56140 14094 56196
rect 22978 56140 22988 56196
rect 23044 56140 23660 56196
rect 23716 56140 24164 56196
rect 32498 56140 32508 56196
rect 32564 56140 35644 56196
rect 35700 56140 36204 56196
rect 36260 56140 36270 56196
rect 37090 56140 37100 56196
rect 37156 56140 38668 56196
rect 11778 56028 11788 56084
rect 11844 56028 12908 56084
rect 12964 56028 14588 56084
rect 14644 56028 14654 56084
rect 13132 55972 13188 56028
rect 24108 55972 24164 56140
rect 38612 56084 38668 56140
rect 35970 56028 35980 56084
rect 36036 56028 37212 56084
rect 37268 56028 37278 56084
rect 38612 56028 39004 56084
rect 39060 56028 39070 56084
rect 50306 56028 50316 56084
rect 50372 56028 51436 56084
rect 51492 56028 51884 56084
rect 51940 56028 51950 56084
rect 4610 55916 4620 55972
rect 4676 55916 5180 55972
rect 5236 55916 6636 55972
rect 6692 55916 6702 55972
rect 13122 55916 13132 55972
rect 13188 55916 13198 55972
rect 14242 55916 14252 55972
rect 14308 55916 15260 55972
rect 15316 55916 15326 55972
rect 24098 55916 24108 55972
rect 24164 55916 24174 55972
rect 41682 55916 41692 55972
rect 41748 55916 42924 55972
rect 42980 55916 42990 55972
rect 45490 55916 45500 55972
rect 45556 55916 46396 55972
rect 46452 55916 46462 55972
rect 23650 55804 23660 55860
rect 23716 55804 24444 55860
rect 24500 55804 24510 55860
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 6178 55468 6188 55524
rect 6244 55468 10332 55524
rect 10388 55468 11004 55524
rect 11060 55468 11070 55524
rect 21298 55468 21308 55524
rect 21364 55468 25228 55524
rect 25284 55468 25294 55524
rect 35186 55468 35196 55524
rect 35252 55468 35980 55524
rect 36036 55468 36046 55524
rect 53890 55468 53900 55524
rect 53956 55468 54908 55524
rect 54964 55468 54974 55524
rect 55122 55468 55132 55524
rect 55188 55468 55198 55524
rect 55132 55412 55188 55468
rect 33618 55356 33628 55412
rect 33684 55356 34860 55412
rect 34916 55356 34926 55412
rect 41570 55356 41580 55412
rect 41636 55356 42140 55412
rect 42196 55356 46732 55412
rect 46788 55356 46798 55412
rect 55132 55356 56476 55412
rect 56532 55356 56542 55412
rect 11330 55244 11340 55300
rect 11396 55244 13468 55300
rect 13524 55244 14476 55300
rect 14532 55244 14542 55300
rect 44258 55244 44268 55300
rect 44324 55244 44940 55300
rect 44996 55244 45006 55300
rect 55010 55244 55020 55300
rect 55076 55244 58156 55300
rect 58212 55244 58222 55300
rect 31602 55132 31612 55188
rect 31668 55132 32284 55188
rect 32340 55132 33068 55188
rect 33124 55132 33134 55188
rect 38322 55132 38332 55188
rect 38388 55132 39564 55188
rect 39620 55132 39630 55188
rect 46946 55132 46956 55188
rect 47012 55132 49308 55188
rect 49364 55132 49980 55188
rect 50036 55132 50046 55188
rect 3154 55020 3164 55076
rect 3220 55020 3836 55076
rect 3892 55020 3902 55076
rect 12674 55020 12684 55076
rect 12740 55020 13580 55076
rect 13636 55020 16940 55076
rect 16996 55020 17006 55076
rect 27010 55020 27020 55076
rect 27076 55020 27916 55076
rect 27972 55020 29372 55076
rect 29428 55020 29438 55076
rect 30818 55020 30828 55076
rect 30884 55020 31500 55076
rect 31556 55020 31566 55076
rect 40450 55020 40460 55076
rect 40516 55020 41468 55076
rect 41524 55020 42364 55076
rect 42420 55020 42430 55076
rect 49522 55020 49532 55076
rect 49588 55020 50428 55076
rect 50484 55020 50494 55076
rect 52882 55020 52892 55076
rect 52948 55020 53788 55076
rect 53844 55020 53854 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 30370 54684 30380 54740
rect 30436 54684 31388 54740
rect 31444 54684 31454 54740
rect 41794 54684 41804 54740
rect 41860 54684 42476 54740
rect 42532 54684 42542 54740
rect 51314 54684 51324 54740
rect 51380 54684 51884 54740
rect 51940 54684 53116 54740
rect 53172 54684 53182 54740
rect 3266 54572 3276 54628
rect 3332 54572 4060 54628
rect 4116 54572 5404 54628
rect 5460 54572 5470 54628
rect 26674 54572 26684 54628
rect 26740 54572 26908 54628
rect 30930 54572 30940 54628
rect 30996 54572 31948 54628
rect 32004 54572 32014 54628
rect 39442 54572 39452 54628
rect 39508 54572 39900 54628
rect 39956 54572 40796 54628
rect 40852 54572 40862 54628
rect 46050 54572 46060 54628
rect 46116 54572 46844 54628
rect 46900 54572 49196 54628
rect 49252 54572 49262 54628
rect 55122 54572 55132 54628
rect 55188 54572 56812 54628
rect 56868 54572 57708 54628
rect 57764 54572 57774 54628
rect 26852 54516 26908 54572
rect 4610 54460 4620 54516
rect 4676 54460 5180 54516
rect 5236 54460 5246 54516
rect 12562 54460 12572 54516
rect 12628 54460 14476 54516
rect 14532 54460 15484 54516
rect 15540 54460 15550 54516
rect 16380 54460 18284 54516
rect 18340 54460 19068 54516
rect 19124 54460 19628 54516
rect 19684 54460 19694 54516
rect 26852 54460 27580 54516
rect 27636 54460 27646 54516
rect 46386 54460 46396 54516
rect 46452 54460 46956 54516
rect 47012 54460 47022 54516
rect 50306 54460 50316 54516
rect 50372 54460 50876 54516
rect 50932 54460 51660 54516
rect 51716 54460 51726 54516
rect 16380 54404 16436 54460
rect 6738 54348 6748 54404
rect 6804 54348 16436 54404
rect 16706 54348 16716 54404
rect 16772 54348 20188 54404
rect 28466 54348 28476 54404
rect 28532 54348 29148 54404
rect 29204 54348 29214 54404
rect 46834 54348 46844 54404
rect 46900 54348 47852 54404
rect 47908 54348 47918 54404
rect 56130 54348 56140 54404
rect 56196 54348 56700 54404
rect 56756 54348 56766 54404
rect 20132 54292 20188 54348
rect 20132 54236 32396 54292
rect 32452 54236 32462 54292
rect 54898 54236 54908 54292
rect 54964 54236 57148 54292
rect 57204 54236 58156 54292
rect 58212 54236 58222 54292
rect 13346 54124 13356 54180
rect 13412 54124 14140 54180
rect 14196 54124 14206 54180
rect 54786 54124 54796 54180
rect 54852 54124 55132 54180
rect 55188 54124 55198 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 23314 54012 23324 54068
rect 23380 54012 24780 54068
rect 24836 54012 30380 54068
rect 30436 54012 30446 54068
rect 41010 54012 41020 54068
rect 41076 54012 42476 54068
rect 42532 54012 44268 54068
rect 44324 54012 44334 54068
rect 3378 53900 3388 53956
rect 3444 53900 4284 53956
rect 4340 53900 4350 53956
rect 29362 53900 29372 53956
rect 29428 53900 31276 53956
rect 31332 53900 31342 53956
rect 40114 53900 40124 53956
rect 40180 53900 43148 53956
rect 43204 53900 43214 53956
rect 51650 53900 51660 53956
rect 51716 53900 52668 53956
rect 52724 53900 52734 53956
rect 17826 53788 17836 53844
rect 17892 53788 18732 53844
rect 18788 53788 18798 53844
rect 20514 53788 20524 53844
rect 20580 53788 20590 53844
rect 21186 53788 21196 53844
rect 21252 53788 22316 53844
rect 22372 53788 22382 53844
rect 28130 53788 28140 53844
rect 28196 53788 28924 53844
rect 28980 53788 28990 53844
rect 36194 53788 36204 53844
rect 36260 53788 37100 53844
rect 37156 53788 37166 53844
rect 37986 53788 37996 53844
rect 38052 53788 42028 53844
rect 42084 53788 42094 53844
rect 47842 53788 47852 53844
rect 47908 53788 52780 53844
rect 52836 53788 52846 53844
rect 52994 53788 53004 53844
rect 53060 53788 55804 53844
rect 55860 53788 55870 53844
rect 20524 53732 20580 53788
rect 19842 53676 19852 53732
rect 19908 53676 20580 53732
rect 20636 53676 30716 53732
rect 30772 53676 30782 53732
rect 34514 53676 34524 53732
rect 34580 53676 36428 53732
rect 36484 53676 36494 53732
rect 44258 53676 44268 53732
rect 44324 53676 45836 53732
rect 45892 53676 45902 53732
rect 20636 53620 20692 53676
rect 7410 53564 7420 53620
rect 7476 53564 7868 53620
rect 7924 53564 9100 53620
rect 9156 53564 9166 53620
rect 19394 53564 19404 53620
rect 19460 53564 20636 53620
rect 20692 53564 20702 53620
rect 23090 53564 23100 53620
rect 23156 53564 23548 53620
rect 23604 53564 24332 53620
rect 24388 53564 24398 53620
rect 39554 53564 39564 53620
rect 39620 53564 40908 53620
rect 40964 53564 45500 53620
rect 45556 53564 45566 53620
rect 20076 53508 20132 53564
rect 51660 53508 51716 53788
rect 5954 53452 5964 53508
rect 6020 53452 7196 53508
rect 7252 53452 7262 53508
rect 17938 53452 17948 53508
rect 18004 53452 18844 53508
rect 18900 53452 19628 53508
rect 19684 53452 19694 53508
rect 20066 53452 20076 53508
rect 20132 53452 20142 53508
rect 23202 53452 23212 53508
rect 23268 53452 23884 53508
rect 23940 53452 23950 53508
rect 29026 53452 29036 53508
rect 29092 53452 30044 53508
rect 30100 53452 30604 53508
rect 30660 53452 30670 53508
rect 40114 53452 40124 53508
rect 40180 53452 41356 53508
rect 41412 53452 41422 53508
rect 51650 53452 51660 53508
rect 51716 53452 51726 53508
rect 52770 53452 52780 53508
rect 52836 53452 53676 53508
rect 53732 53452 53742 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 20626 53228 20636 53284
rect 20692 53228 21308 53284
rect 21364 53228 21374 53284
rect 47506 53228 47516 53284
rect 47572 53228 47964 53284
rect 48020 53228 48030 53284
rect 7634 53116 7644 53172
rect 7700 53116 8652 53172
rect 8708 53116 8718 53172
rect 24658 53116 24668 53172
rect 24724 53116 25340 53172
rect 25396 53116 25406 53172
rect 31266 53116 31276 53172
rect 31332 53116 32172 53172
rect 32228 53116 32238 53172
rect 35970 53116 35980 53172
rect 36036 53116 36316 53172
rect 36372 53116 37324 53172
rect 37380 53116 37390 53172
rect 46834 53116 46844 53172
rect 46900 53116 51548 53172
rect 51604 53116 51614 53172
rect 4274 53004 4284 53060
rect 4340 53004 4956 53060
rect 5012 53004 9996 53060
rect 10052 53004 10332 53060
rect 10388 53004 10398 53060
rect 12898 53004 12908 53060
rect 12964 53004 14812 53060
rect 14868 53004 14878 53060
rect 35634 53004 35644 53060
rect 35700 53004 36652 53060
rect 36708 53004 36718 53060
rect 38546 53004 38556 53060
rect 38612 53004 41020 53060
rect 41076 53004 41086 53060
rect 50978 53004 50988 53060
rect 51044 53004 51660 53060
rect 51716 53004 51726 53060
rect 8372 52836 8428 52948
rect 8484 52892 8494 52948
rect 8642 52892 8652 52948
rect 8708 52892 9100 52948
rect 9156 52892 9166 52948
rect 17490 52892 17500 52948
rect 17556 52892 20636 52948
rect 20692 52892 20702 52948
rect 23090 52892 23100 52948
rect 23156 52892 24220 52948
rect 24276 52892 24286 52948
rect 34402 52892 34412 52948
rect 34468 52892 35980 52948
rect 36036 52892 36764 52948
rect 36820 52892 36830 52948
rect 46386 52892 46396 52948
rect 46452 52892 46732 52948
rect 46788 52892 47516 52948
rect 47572 52892 47582 52948
rect 7298 52780 7308 52836
rect 7364 52780 8428 52836
rect 10658 52780 10668 52836
rect 10724 52780 12348 52836
rect 12404 52780 12414 52836
rect 20290 52780 20300 52836
rect 20356 52780 20524 52836
rect 20580 52780 20590 52836
rect 30706 52780 30716 52836
rect 30772 52780 31948 52836
rect 32004 52780 32014 52836
rect 43810 52780 43820 52836
rect 43876 52780 46508 52836
rect 46564 52780 46574 52836
rect 57362 52780 57372 52836
rect 57428 52780 58156 52836
rect 58212 52780 58222 52836
rect 47170 52668 47180 52724
rect 47236 52668 51324 52724
rect 51380 52668 51390 52724
rect 19618 52556 19628 52612
rect 19684 52556 20524 52612
rect 20580 52556 20590 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 16482 52444 16492 52500
rect 16548 52444 32508 52500
rect 32564 52444 33292 52500
rect 33348 52444 33516 52500
rect 33572 52444 33582 52500
rect 20738 52332 20748 52388
rect 20804 52332 23100 52388
rect 23156 52332 23166 52388
rect 33170 52332 33180 52388
rect 33236 52332 35644 52388
rect 35700 52332 35710 52388
rect 56130 52332 56140 52388
rect 56196 52332 56588 52388
rect 56644 52332 56654 52388
rect 59200 52276 60000 52304
rect 8194 52220 8204 52276
rect 8260 52220 8652 52276
rect 8708 52220 10108 52276
rect 10164 52220 11452 52276
rect 11508 52220 11518 52276
rect 14914 52220 14924 52276
rect 14980 52220 15988 52276
rect 30930 52220 30940 52276
rect 30996 52220 31948 52276
rect 32004 52220 32014 52276
rect 32386 52220 32396 52276
rect 32452 52220 33740 52276
rect 33796 52220 33806 52276
rect 45490 52220 45500 52276
rect 45556 52220 46732 52276
rect 46788 52220 46798 52276
rect 53330 52220 53340 52276
rect 53396 52220 57596 52276
rect 57652 52220 57662 52276
rect 58146 52220 58156 52276
rect 58212 52220 60000 52276
rect 15932 52164 15988 52220
rect 59200 52192 60000 52220
rect 3826 52108 3836 52164
rect 3892 52108 4620 52164
rect 4676 52108 6748 52164
rect 6804 52108 6814 52164
rect 9650 52108 9660 52164
rect 9716 52108 10220 52164
rect 10276 52108 12964 52164
rect 14466 52108 14476 52164
rect 14532 52108 15260 52164
rect 15316 52108 15326 52164
rect 15922 52108 15932 52164
rect 15988 52108 15998 52164
rect 19170 52108 19180 52164
rect 19236 52108 20300 52164
rect 20356 52108 20366 52164
rect 31826 52108 31836 52164
rect 31892 52108 32284 52164
rect 32340 52108 33852 52164
rect 33908 52108 33918 52164
rect 53218 52108 53228 52164
rect 53284 52108 53676 52164
rect 53732 52108 54124 52164
rect 54180 52108 55132 52164
rect 55188 52108 55198 52164
rect 7970 51996 7980 52052
rect 8036 51996 8764 52052
rect 8820 51996 8830 52052
rect 12908 51828 12964 52108
rect 43138 51996 43148 52052
rect 43204 51996 44156 52052
rect 44212 51996 44222 52052
rect 12898 51772 12908 51828
rect 12964 51772 13468 51828
rect 13524 51772 13534 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 11778 51548 11788 51604
rect 11844 51548 13356 51604
rect 13412 51548 13916 51604
rect 13972 51548 13982 51604
rect 42466 51548 42476 51604
rect 42532 51548 43260 51604
rect 43316 51548 43708 51604
rect 43764 51548 43774 51604
rect 55458 51548 55468 51604
rect 55524 51548 57036 51604
rect 57092 51548 58156 51604
rect 58212 51548 58222 51604
rect 14354 51436 14364 51492
rect 14420 51436 15036 51492
rect 15092 51436 15102 51492
rect 22418 51436 22428 51492
rect 22484 51436 23772 51492
rect 23828 51436 23838 51492
rect 54674 51436 54684 51492
rect 54740 51436 56812 51492
rect 56868 51436 56878 51492
rect 3378 51324 3388 51380
rect 3444 51324 5068 51380
rect 5124 51324 5134 51380
rect 43250 51324 43260 51380
rect 43316 51324 47292 51380
rect 47348 51324 47358 51380
rect 52434 51324 52444 51380
rect 52500 51324 52510 51380
rect 56466 51324 56476 51380
rect 56532 51324 56542 51380
rect 3266 51212 3276 51268
rect 3332 51212 3948 51268
rect 4004 51212 5516 51268
rect 5572 51212 5582 51268
rect 28018 51212 28028 51268
rect 28084 51212 36148 51268
rect 36754 51212 36764 51268
rect 36820 51212 37772 51268
rect 37828 51212 38556 51268
rect 38612 51212 38622 51268
rect 41794 51212 41804 51268
rect 41860 51212 42252 51268
rect 42308 51212 45276 51268
rect 45332 51212 45342 51268
rect 36092 51156 36148 51212
rect 52444 51156 52500 51324
rect 56476 51268 56532 51324
rect 55346 51212 55356 51268
rect 55412 51212 56532 51268
rect 4274 51100 4284 51156
rect 4340 51100 4396 51156
rect 4452 51100 4462 51156
rect 7634 51100 7644 51156
rect 7700 51100 11116 51156
rect 11172 51100 11182 51156
rect 28578 51100 28588 51156
rect 28644 51100 29260 51156
rect 29316 51100 29326 51156
rect 36082 51100 36092 51156
rect 36148 51100 36158 51156
rect 51090 51100 51100 51156
rect 51156 51100 51772 51156
rect 51828 51100 52500 51156
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 11554 50876 11564 50932
rect 11620 50876 17500 50932
rect 17556 50876 17566 50932
rect 28242 50876 28252 50932
rect 28308 50876 29708 50932
rect 29764 50876 32284 50932
rect 32340 50876 32350 50932
rect 29362 50764 29372 50820
rect 29428 50764 30940 50820
rect 30996 50764 31006 50820
rect 41010 50764 41020 50820
rect 41076 50764 41804 50820
rect 41860 50764 41870 50820
rect 53218 50764 53228 50820
rect 53284 50764 54012 50820
rect 54068 50764 54078 50820
rect 5506 50652 5516 50708
rect 5572 50652 11564 50708
rect 11620 50652 12236 50708
rect 12292 50652 12302 50708
rect 29810 50652 29820 50708
rect 29876 50652 30716 50708
rect 30772 50652 30782 50708
rect 45836 50652 51212 50708
rect 51268 50652 51278 50708
rect 45836 50596 45892 50652
rect 3602 50540 3612 50596
rect 3668 50540 5628 50596
rect 5684 50540 5694 50596
rect 29586 50540 29596 50596
rect 29652 50540 30156 50596
rect 30212 50540 30222 50596
rect 41458 50540 41468 50596
rect 41524 50540 42812 50596
rect 42868 50540 42878 50596
rect 44146 50540 44156 50596
rect 44212 50540 44828 50596
rect 44884 50540 45836 50596
rect 45892 50540 45902 50596
rect 46050 50540 46060 50596
rect 46116 50540 46732 50596
rect 46788 50540 47628 50596
rect 47684 50540 47694 50596
rect 4050 50428 4060 50484
rect 4116 50428 5740 50484
rect 5796 50428 5806 50484
rect 26226 50428 26236 50484
rect 26292 50428 30604 50484
rect 30660 50428 30670 50484
rect 4246 50316 4284 50372
rect 4340 50316 4350 50372
rect 4620 50260 4676 50428
rect 4620 50204 4732 50260
rect 4788 50204 4798 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 2482 49980 2492 50036
rect 2548 49980 4508 50036
rect 4564 49980 4574 50036
rect 21970 49980 21980 50036
rect 22036 49980 28812 50036
rect 28868 49980 30492 50036
rect 30548 49980 30558 50036
rect 39330 49980 39340 50036
rect 39396 49980 41020 50036
rect 41076 49980 42140 50036
rect 42196 49980 42206 50036
rect 8642 49868 8652 49924
rect 8708 49868 9212 49924
rect 9268 49868 10220 49924
rect 10276 49868 10286 49924
rect 19282 49868 19292 49924
rect 19348 49868 20300 49924
rect 20356 49868 20366 49924
rect 31892 49868 32508 49924
rect 32564 49868 32574 49924
rect 37762 49868 37772 49924
rect 37828 49868 38556 49924
rect 38612 49868 38622 49924
rect 50754 49868 50764 49924
rect 50820 49868 52668 49924
rect 52724 49868 54460 49924
rect 54516 49868 54526 49924
rect 8866 49756 8876 49812
rect 8932 49756 9324 49812
rect 9380 49756 10332 49812
rect 10388 49756 12684 49812
rect 12740 49756 12750 49812
rect 13234 49756 13244 49812
rect 13300 49756 14364 49812
rect 14420 49756 14430 49812
rect 19394 49756 19404 49812
rect 19460 49756 21420 49812
rect 21476 49756 21486 49812
rect 28690 49756 28700 49812
rect 28756 49756 29820 49812
rect 29876 49756 29886 49812
rect 31892 49700 31948 49868
rect 32722 49756 32732 49812
rect 32788 49756 33404 49812
rect 33460 49756 33470 49812
rect 34178 49756 34188 49812
rect 34244 49756 35084 49812
rect 35140 49756 35150 49812
rect 41458 49756 41468 49812
rect 41524 49756 42252 49812
rect 42308 49756 42318 49812
rect 10770 49644 10780 49700
rect 10836 49644 12348 49700
rect 12404 49644 13692 49700
rect 13748 49644 13916 49700
rect 13972 49644 13982 49700
rect 19170 49644 19180 49700
rect 19236 49644 19740 49700
rect 19796 49644 20524 49700
rect 20580 49644 31164 49700
rect 31220 49644 31948 49700
rect 42130 49644 42140 49700
rect 42196 49644 43372 49700
rect 43428 49644 43438 49700
rect 47394 49532 47404 49588
rect 47460 49532 48860 49588
rect 48916 49532 48926 49588
rect 27346 49420 27356 49476
rect 27412 49420 34860 49476
rect 34916 49420 34926 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 39666 49308 39676 49364
rect 39732 49308 50876 49364
rect 50932 49308 51660 49364
rect 51716 49308 51726 49364
rect 16258 49196 16268 49252
rect 16324 49196 33012 49252
rect 32956 49140 33012 49196
rect 8530 49084 8540 49140
rect 8596 49084 9100 49140
rect 9156 49084 9166 49140
rect 16706 49084 16716 49140
rect 16772 49084 19068 49140
rect 19124 49084 22540 49140
rect 22596 49084 22988 49140
rect 23044 49084 25116 49140
rect 25172 49084 25182 49140
rect 30482 49084 30492 49140
rect 30548 49084 31948 49140
rect 32946 49084 32956 49140
rect 33012 49084 33740 49140
rect 33796 49084 33806 49140
rect 55412 49084 56140 49140
rect 56196 49084 58156 49140
rect 58212 49084 58222 49140
rect 31892 49028 31948 49084
rect 5394 48972 5404 49028
rect 5460 48972 6076 49028
rect 6132 48972 10108 49028
rect 10164 48972 10174 49028
rect 31892 48972 35084 49028
rect 35140 48972 35150 49028
rect 49970 48972 49980 49028
rect 50036 48972 50652 49028
rect 50708 48972 51548 49028
rect 51604 48972 51614 49028
rect 54898 48972 54908 49028
rect 54964 48972 55356 49028
rect 55412 48972 55468 49084
rect 6738 48860 6748 48916
rect 6804 48860 9324 48916
rect 9380 48860 9390 48916
rect 17378 48860 17388 48916
rect 17444 48860 20188 48916
rect 20244 48860 20254 48916
rect 20626 48860 20636 48916
rect 20692 48860 21420 48916
rect 21476 48860 21486 48916
rect 8418 48748 8428 48804
rect 8484 48748 9660 48804
rect 9716 48748 9726 48804
rect 20066 48748 20076 48804
rect 20132 48748 20524 48804
rect 20580 48748 21308 48804
rect 21364 48748 21374 48804
rect 23650 48748 23660 48804
rect 23716 48748 24444 48804
rect 24500 48748 25788 48804
rect 25844 48748 25854 48804
rect 20402 48636 20412 48692
rect 20468 48636 21532 48692
rect 21588 48636 21598 48692
rect 54674 48636 54684 48692
rect 54740 48636 55692 48692
rect 55748 48636 55758 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 8306 48412 8316 48468
rect 8372 48412 9548 48468
rect 9604 48412 9614 48468
rect 8082 48300 8092 48356
rect 8148 48300 8764 48356
rect 8820 48300 8830 48356
rect 9986 48300 9996 48356
rect 10052 48300 10556 48356
rect 10612 48300 11340 48356
rect 11396 48300 11406 48356
rect 28354 48300 28364 48356
rect 28420 48300 29372 48356
rect 29428 48300 29438 48356
rect 42354 48300 42364 48356
rect 42420 48300 43372 48356
rect 43428 48300 43438 48356
rect 49186 48300 49196 48356
rect 49252 48300 53900 48356
rect 53956 48300 53966 48356
rect 54786 48300 54796 48356
rect 54852 48300 55468 48356
rect 55524 48300 55534 48356
rect 11106 48188 11116 48244
rect 11172 48188 12572 48244
rect 12628 48188 13356 48244
rect 13412 48188 13422 48244
rect 26114 48188 26124 48244
rect 26180 48188 27468 48244
rect 27524 48188 27534 48244
rect 27682 48188 27692 48244
rect 27748 48188 28252 48244
rect 28308 48188 28318 48244
rect 43026 48188 43036 48244
rect 43092 48188 43484 48244
rect 43540 48188 43550 48244
rect 45266 48188 45276 48244
rect 45332 48188 49084 48244
rect 49140 48188 49644 48244
rect 49700 48188 49710 48244
rect 13682 48076 13692 48132
rect 13748 48076 14812 48132
rect 14868 48076 16604 48132
rect 16660 48076 16670 48132
rect 20962 48076 20972 48132
rect 21028 48076 21980 48132
rect 22036 48076 23436 48132
rect 23492 48076 23502 48132
rect 41570 48076 41580 48132
rect 41636 48076 42588 48132
rect 42644 48076 42654 48132
rect 47954 48076 47964 48132
rect 48020 48076 48860 48132
rect 48916 48076 49196 48132
rect 49252 48076 49262 48132
rect 54226 48076 54236 48132
rect 54292 48076 54908 48132
rect 54964 48076 54974 48132
rect 23762 47964 23772 48020
rect 23828 47964 24668 48020
rect 24724 47964 24734 48020
rect 27906 47964 27916 48020
rect 27972 47964 28364 48020
rect 28420 47964 28430 48020
rect 13346 47852 13356 47908
rect 13412 47852 13692 47908
rect 13748 47852 13758 47908
rect 42690 47852 42700 47908
rect 42756 47852 49756 47908
rect 49812 47852 50092 47908
rect 50148 47852 50158 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 9538 47628 9548 47684
rect 9604 47628 11116 47684
rect 11172 47628 11182 47684
rect 21522 47628 21532 47684
rect 21588 47628 22652 47684
rect 22708 47628 22718 47684
rect 35410 47628 35420 47684
rect 35476 47628 36652 47684
rect 36708 47628 37436 47684
rect 37492 47628 37502 47684
rect 1810 47516 1820 47572
rect 1876 47516 5068 47572
rect 5124 47516 5134 47572
rect 15250 47516 15260 47572
rect 15316 47516 16492 47572
rect 16548 47516 16558 47572
rect 23090 47516 23100 47572
rect 23156 47516 24332 47572
rect 24388 47516 24398 47572
rect 28466 47516 28476 47572
rect 28532 47516 34636 47572
rect 34692 47516 34972 47572
rect 35028 47516 35038 47572
rect 38098 47516 38108 47572
rect 38164 47516 41692 47572
rect 41748 47516 41758 47572
rect 42130 47516 42140 47572
rect 42196 47516 42924 47572
rect 42980 47516 43596 47572
rect 43652 47516 44268 47572
rect 44324 47516 44828 47572
rect 44884 47516 44894 47572
rect 9650 47404 9660 47460
rect 9716 47404 11116 47460
rect 11172 47404 11788 47460
rect 11844 47404 11854 47460
rect 12226 47404 12236 47460
rect 12292 47404 13356 47460
rect 13412 47404 13422 47460
rect 14018 47404 14028 47460
rect 14084 47404 16380 47460
rect 16436 47404 17612 47460
rect 17668 47404 17678 47460
rect 18162 47404 18172 47460
rect 18228 47404 19068 47460
rect 19124 47404 19134 47460
rect 23650 47404 23660 47460
rect 23716 47404 24556 47460
rect 24612 47404 24622 47460
rect 36418 47404 36428 47460
rect 36484 47404 38444 47460
rect 38500 47404 38510 47460
rect 49858 47404 49868 47460
rect 49924 47404 52668 47460
rect 52724 47404 53676 47460
rect 53732 47404 56252 47460
rect 56308 47404 56318 47460
rect 4610 47292 4620 47348
rect 4676 47292 5292 47348
rect 5348 47292 5740 47348
rect 5796 47292 5806 47348
rect 11330 47292 11340 47348
rect 11396 47292 13580 47348
rect 13636 47292 13646 47348
rect 36082 47292 36092 47348
rect 36148 47292 39004 47348
rect 39060 47292 39070 47348
rect 18274 47180 18284 47236
rect 18340 47180 23660 47236
rect 23716 47180 23726 47236
rect 24882 47180 24892 47236
rect 24948 47180 27244 47236
rect 27300 47180 27692 47236
rect 27748 47180 27758 47236
rect 37090 47180 37100 47236
rect 37156 47180 37660 47236
rect 37716 47180 38556 47236
rect 38612 47180 38622 47236
rect 43474 47180 43484 47236
rect 43540 47180 44828 47236
rect 44884 47180 47740 47236
rect 47796 47180 47806 47236
rect 14690 47068 14700 47124
rect 14756 47068 15820 47124
rect 15876 47068 15886 47124
rect 17938 47068 17948 47124
rect 18004 47068 18620 47124
rect 18676 47068 18686 47124
rect 24322 47068 24332 47124
rect 24388 47068 25452 47124
rect 25508 47068 46228 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 46172 47012 46228 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 5506 46956 5516 47012
rect 5572 46956 6300 47012
rect 6356 46956 13468 47012
rect 13524 46956 13534 47012
rect 26450 46956 26460 47012
rect 26516 46956 27468 47012
rect 27524 46956 27534 47012
rect 43922 46956 43932 47012
rect 43988 46956 45276 47012
rect 45332 46956 45948 47012
rect 46004 46956 46014 47012
rect 46172 46956 48804 47012
rect 11778 46844 11788 46900
rect 11844 46844 13132 46900
rect 13188 46844 13198 46900
rect 24546 46844 24556 46900
rect 24612 46844 30100 46900
rect 32050 46844 32060 46900
rect 32116 46844 32508 46900
rect 32564 46844 37548 46900
rect 37604 46844 37614 46900
rect 38322 46844 38332 46900
rect 38388 46844 47628 46900
rect 47684 46844 47694 46900
rect 30044 46788 30100 46844
rect 48748 46788 48804 46956
rect 28690 46732 28700 46788
rect 28756 46732 29820 46788
rect 29876 46732 29886 46788
rect 30044 46732 34748 46788
rect 34804 46732 34814 46788
rect 39890 46732 39900 46788
rect 39956 46732 43260 46788
rect 43316 46732 43708 46788
rect 48738 46732 48748 46788
rect 48804 46732 48814 46788
rect 43652 46676 43708 46732
rect 13122 46620 13132 46676
rect 13188 46620 14476 46676
rect 14532 46620 14542 46676
rect 19394 46620 19404 46676
rect 19460 46620 23548 46676
rect 23604 46620 25228 46676
rect 25284 46620 25294 46676
rect 35858 46620 35868 46676
rect 35924 46620 36652 46676
rect 36708 46620 37436 46676
rect 37492 46620 37502 46676
rect 37650 46620 37660 46676
rect 37716 46620 38892 46676
rect 38948 46620 38958 46676
rect 43652 46620 44492 46676
rect 44548 46620 44558 46676
rect 45378 46620 45388 46676
rect 45444 46620 45724 46676
rect 45780 46620 45790 46676
rect 49298 46620 49308 46676
rect 49364 46620 49756 46676
rect 49812 46620 50540 46676
rect 50596 46620 50606 46676
rect 2706 46508 2716 46564
rect 2772 46508 3500 46564
rect 3556 46508 3566 46564
rect 15922 46508 15932 46564
rect 15988 46508 26012 46564
rect 26068 46508 26078 46564
rect 45042 46508 45052 46564
rect 45108 46508 45836 46564
rect 45892 46508 45902 46564
rect 47618 46508 47628 46564
rect 47684 46508 53004 46564
rect 53060 46508 53070 46564
rect 54898 46508 54908 46564
rect 54964 46508 55692 46564
rect 55748 46508 55758 46564
rect 19730 46396 19740 46452
rect 19796 46396 35756 46452
rect 35812 46396 36316 46452
rect 36372 46396 37100 46452
rect 37156 46396 37166 46452
rect 39554 46396 39564 46452
rect 39620 46396 40908 46452
rect 40964 46396 40974 46452
rect 47842 46396 47852 46452
rect 47908 46396 50092 46452
rect 50148 46396 52108 46452
rect 52164 46396 52174 46452
rect 22978 46284 22988 46340
rect 23044 46284 23660 46340
rect 23716 46284 23726 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 15092 46172 20188 46228
rect 20244 46172 21084 46228
rect 21140 46172 21150 46228
rect 30146 46172 30156 46228
rect 30212 46172 31164 46228
rect 31220 46172 31948 46228
rect 32004 46172 32014 46228
rect 15092 46116 15148 46172
rect 11890 46060 11900 46116
rect 11956 46060 12796 46116
rect 12852 46060 14028 46116
rect 14084 46060 15148 46116
rect 18162 46060 18172 46116
rect 18228 46060 26236 46116
rect 26292 46060 26460 46116
rect 26516 46060 26526 46116
rect 13570 45948 13580 46004
rect 13636 45948 19292 46004
rect 19348 45948 19358 46004
rect 29810 45948 29820 46004
rect 29876 45948 31052 46004
rect 31108 45948 31118 46004
rect 15810 45836 15820 45892
rect 15876 45836 17052 45892
rect 17108 45836 17118 45892
rect 48402 45836 48412 45892
rect 48468 45836 49532 45892
rect 49588 45836 49598 45892
rect 54898 45836 54908 45892
rect 54964 45836 58044 45892
rect 58100 45836 58110 45892
rect 14812 45724 15484 45780
rect 15540 45724 15550 45780
rect 32050 45724 32060 45780
rect 32116 45724 33180 45780
rect 33236 45724 33246 45780
rect 49298 45724 49308 45780
rect 49364 45724 49980 45780
rect 50036 45724 50046 45780
rect 14812 45668 14868 45724
rect 8754 45612 8764 45668
rect 8820 45612 8988 45668
rect 9044 45612 9996 45668
rect 10052 45612 14812 45668
rect 14868 45612 14878 45668
rect 15362 45612 15372 45668
rect 15428 45612 15820 45668
rect 15876 45612 15886 45668
rect 20738 45612 20748 45668
rect 20804 45612 21420 45668
rect 21476 45612 37996 45668
rect 38052 45612 48076 45668
rect 48132 45612 48142 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 9426 45388 9436 45444
rect 9492 45388 12796 45444
rect 12852 45388 13580 45444
rect 13636 45388 13646 45444
rect 37538 45388 37548 45444
rect 37604 45388 38332 45444
rect 38388 45388 38398 45444
rect 59200 45332 60000 45360
rect 8306 45276 8316 45332
rect 8372 45276 8382 45332
rect 8866 45276 8876 45332
rect 8932 45276 9772 45332
rect 9828 45276 9838 45332
rect 12450 45276 12460 45332
rect 12516 45276 18788 45332
rect 22306 45276 22316 45332
rect 22372 45276 23324 45332
rect 23380 45276 23390 45332
rect 34402 45276 34412 45332
rect 34468 45276 36204 45332
rect 36260 45276 36652 45332
rect 36708 45276 38892 45332
rect 38948 45276 38958 45332
rect 40674 45276 40684 45332
rect 40740 45276 41916 45332
rect 41972 45276 41982 45332
rect 55010 45276 55020 45332
rect 55076 45276 55692 45332
rect 55748 45276 56924 45332
rect 56980 45276 56990 45332
rect 58146 45276 58156 45332
rect 58212 45276 60000 45332
rect 8316 45220 8372 45276
rect 7522 45164 7532 45220
rect 7588 45164 10108 45220
rect 10164 45164 10174 45220
rect 14018 45164 14028 45220
rect 14084 45164 14252 45220
rect 14308 45164 14476 45220
rect 14532 45164 14812 45220
rect 14868 45164 14878 45220
rect 6066 45052 6076 45108
rect 6132 45052 9436 45108
rect 9492 45052 9502 45108
rect 15026 45052 15036 45108
rect 15092 45052 15820 45108
rect 15876 45052 15886 45108
rect 18732 44996 18788 45276
rect 59200 45248 60000 45276
rect 21634 45164 21644 45220
rect 21700 45164 22204 45220
rect 22260 45164 22270 45220
rect 31826 45164 31836 45220
rect 31892 45164 34076 45220
rect 34132 45164 34142 45220
rect 49074 45164 49084 45220
rect 49140 45164 50988 45220
rect 51044 45164 51054 45220
rect 21746 45052 21756 45108
rect 21812 45052 22428 45108
rect 22484 45052 22494 45108
rect 24770 45052 24780 45108
rect 24836 45052 25340 45108
rect 25396 45052 26236 45108
rect 26292 45052 26302 45108
rect 27906 45052 27916 45108
rect 27972 45052 28476 45108
rect 28532 45052 29148 45108
rect 29204 45052 29214 45108
rect 49970 45052 49980 45108
rect 50036 45052 53340 45108
rect 53396 45052 54908 45108
rect 54964 45052 54974 45108
rect 55412 45052 57036 45108
rect 57092 45052 57102 45108
rect 55412 44996 55468 45052
rect 18722 44940 18732 44996
rect 18788 44940 20972 44996
rect 21028 44940 30156 44996
rect 30212 44940 30222 44996
rect 33954 44940 33964 44996
rect 34020 44940 35420 44996
rect 35476 44940 35486 44996
rect 51874 44940 51884 44996
rect 51940 44940 52892 44996
rect 52948 44940 52958 44996
rect 55122 44940 55132 44996
rect 55188 44940 55468 44996
rect 22194 44828 22204 44884
rect 22260 44828 23100 44884
rect 23156 44828 23166 44884
rect 40226 44828 40236 44884
rect 40292 44828 44940 44884
rect 44996 44828 45006 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 5282 44492 5292 44548
rect 5348 44492 5964 44548
rect 6020 44492 13524 44548
rect 54562 44492 54572 44548
rect 54628 44492 55244 44548
rect 55300 44492 56140 44548
rect 56196 44492 56206 44548
rect 13468 44436 13524 44492
rect 3378 44380 3388 44436
rect 3444 44380 4508 44436
rect 4564 44380 5628 44436
rect 5684 44380 5694 44436
rect 7186 44380 7196 44436
rect 7252 44380 8092 44436
rect 8148 44380 8158 44436
rect 13458 44380 13468 44436
rect 13524 44380 15372 44436
rect 15428 44380 15438 44436
rect 15810 44380 15820 44436
rect 15876 44380 16156 44436
rect 16212 44380 16222 44436
rect 35634 44380 35644 44436
rect 35700 44380 39116 44436
rect 39172 44380 39182 44436
rect 56242 44380 56252 44436
rect 56308 44380 57596 44436
rect 57652 44380 57662 44436
rect 4834 44268 4844 44324
rect 4900 44268 6188 44324
rect 6244 44268 6254 44324
rect 21634 44268 21644 44324
rect 21700 44268 22092 44324
rect 22148 44268 24444 44324
rect 24500 44268 24510 44324
rect 31154 44268 31164 44324
rect 31220 44268 31836 44324
rect 31892 44268 32620 44324
rect 32676 44268 33292 44324
rect 33348 44268 33358 44324
rect 38882 44268 38892 44324
rect 38948 44268 40796 44324
rect 40852 44268 42140 44324
rect 42196 44268 42206 44324
rect 55346 44268 55356 44324
rect 55412 44268 56588 44324
rect 56644 44268 56654 44324
rect 23314 44156 23324 44212
rect 23380 44156 24108 44212
rect 24164 44156 24174 44212
rect 24658 44156 24668 44212
rect 24724 44156 25564 44212
rect 25620 44156 31388 44212
rect 31444 44156 32172 44212
rect 32228 44156 32238 44212
rect 33058 44156 33068 44212
rect 33124 44156 33628 44212
rect 33684 44156 33694 44212
rect 34066 44156 34076 44212
rect 34132 44156 34916 44212
rect 56018 44156 56028 44212
rect 56084 44156 56700 44212
rect 56756 44156 56766 44212
rect 33628 44100 33684 44156
rect 34860 44100 34916 44156
rect 33628 44044 34636 44100
rect 34692 44044 34702 44100
rect 34850 44044 34860 44100
rect 34916 44044 43372 44100
rect 43428 44044 43438 44100
rect 54338 44044 54348 44100
rect 54404 44044 55468 44100
rect 55524 44044 55534 44100
rect 23202 43932 23212 43988
rect 23268 43932 23660 43988
rect 23716 43932 33628 43988
rect 33684 43932 33694 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 16370 43820 16380 43876
rect 16436 43820 17836 43876
rect 17892 43820 17902 43876
rect 2370 43708 2380 43764
rect 2436 43708 2604 43764
rect 2660 43708 2670 43764
rect 18050 43708 18060 43764
rect 18116 43708 20188 43764
rect 20244 43708 20254 43764
rect 25890 43708 25900 43764
rect 25956 43708 35084 43764
rect 35140 43708 35150 43764
rect 51762 43708 51772 43764
rect 51828 43708 54908 43764
rect 54964 43708 54974 43764
rect 53564 43652 53620 43708
rect 3602 43596 3612 43652
rect 3668 43596 5068 43652
rect 5124 43596 5134 43652
rect 5506 43596 5516 43652
rect 5572 43596 8428 43652
rect 8484 43596 8494 43652
rect 18610 43596 18620 43652
rect 18676 43596 21196 43652
rect 21252 43596 21262 43652
rect 29810 43596 29820 43652
rect 29876 43596 31276 43652
rect 31332 43596 31342 43652
rect 53554 43596 53564 43652
rect 53620 43596 53630 43652
rect 13458 43484 13468 43540
rect 13524 43484 15484 43540
rect 15540 43484 15550 43540
rect 19058 43484 19068 43540
rect 19124 43484 20860 43540
rect 20916 43484 22092 43540
rect 22148 43484 22158 43540
rect 28354 43484 28364 43540
rect 28420 43484 29932 43540
rect 29988 43484 29998 43540
rect 30146 43484 30156 43540
rect 30212 43484 33852 43540
rect 33908 43484 41020 43540
rect 41076 43484 41468 43540
rect 41524 43484 52780 43540
rect 52836 43484 53228 43540
rect 53284 43484 53294 43540
rect 16146 43372 16156 43428
rect 16212 43372 17164 43428
rect 17220 43372 17230 43428
rect 19730 43372 19740 43428
rect 19796 43372 22316 43428
rect 22372 43372 22382 43428
rect 40338 43372 40348 43428
rect 40404 43372 42252 43428
rect 42308 43372 42318 43428
rect 42466 43372 42476 43428
rect 42532 43372 43036 43428
rect 43092 43372 44940 43428
rect 44996 43372 45006 43428
rect 46610 43372 46620 43428
rect 46676 43372 46844 43428
rect 46900 43372 48188 43428
rect 48244 43372 48254 43428
rect 13570 43260 13580 43316
rect 13636 43260 36428 43316
rect 36484 43260 38108 43316
rect 38164 43260 38174 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 14130 43036 14140 43092
rect 14196 43036 32620 43092
rect 32676 43036 33516 43092
rect 33572 43036 33582 43092
rect 16146 42924 16156 42980
rect 16212 42924 18396 42980
rect 18452 42924 20300 42980
rect 20356 42924 20366 42980
rect 37762 42924 37772 42980
rect 37828 42924 39004 42980
rect 39060 42924 40796 42980
rect 40852 42924 40862 42980
rect 42242 42924 42252 42980
rect 42308 42924 43484 42980
rect 43540 42924 43550 42980
rect 44146 42924 44156 42980
rect 44212 42924 45612 42980
rect 45668 42924 45678 42980
rect 14690 42812 14700 42868
rect 14756 42812 16380 42868
rect 16436 42812 16446 42868
rect 27794 42812 27804 42868
rect 27860 42812 29708 42868
rect 29764 42812 31276 42868
rect 31332 42812 31342 42868
rect 8866 42700 8876 42756
rect 8932 42700 9660 42756
rect 9716 42700 9726 42756
rect 15026 42700 15036 42756
rect 15092 42700 15484 42756
rect 15540 42700 16492 42756
rect 16548 42700 16558 42756
rect 26002 42700 26012 42756
rect 26068 42700 27132 42756
rect 27188 42700 29148 42756
rect 29204 42700 29214 42756
rect 45602 42700 45612 42756
rect 45668 42700 46620 42756
rect 46676 42700 46686 42756
rect 14914 42588 14924 42644
rect 14980 42588 21308 42644
rect 21364 42588 21374 42644
rect 39778 42588 39788 42644
rect 39844 42588 40572 42644
rect 40628 42588 40638 42644
rect 41682 42588 41692 42644
rect 41748 42588 42028 42644
rect 42084 42588 42094 42644
rect 50194 42588 50204 42644
rect 50260 42588 51660 42644
rect 51716 42588 51726 42644
rect 8754 42476 8764 42532
rect 8820 42476 9772 42532
rect 9828 42476 12348 42532
rect 12404 42476 12414 42532
rect 12898 42476 12908 42532
rect 12964 42476 13804 42532
rect 13860 42476 13870 42532
rect 15810 42476 15820 42532
rect 15876 42476 21084 42532
rect 21140 42476 21532 42532
rect 21588 42476 21598 42532
rect 28578 42476 28588 42532
rect 28644 42476 30940 42532
rect 30996 42476 31006 42532
rect 45266 42476 45276 42532
rect 45332 42476 45948 42532
rect 46004 42476 46396 42532
rect 46452 42476 46462 42532
rect 51426 42476 51436 42532
rect 51492 42476 53116 42532
rect 53172 42476 53900 42532
rect 53956 42476 55132 42532
rect 55188 42476 55198 42532
rect 33618 42364 33628 42420
rect 33684 42364 39452 42420
rect 39508 42364 39518 42420
rect 43922 42364 43932 42420
rect 43988 42364 45500 42420
rect 45556 42364 45566 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 9874 42140 9884 42196
rect 9940 42140 10556 42196
rect 10612 42140 10622 42196
rect 12114 42140 12124 42196
rect 12180 42140 13468 42196
rect 13524 42140 13534 42196
rect 19954 42140 19964 42196
rect 20020 42140 20748 42196
rect 20804 42140 20814 42196
rect 27244 42140 27916 42196
rect 27972 42140 28364 42196
rect 28420 42140 28430 42196
rect 33618 42140 33628 42196
rect 33684 42140 34076 42196
rect 34132 42140 34142 42196
rect 27244 42084 27300 42140
rect 1810 42028 1820 42084
rect 1876 42028 5068 42084
rect 5124 42028 5404 42084
rect 5460 42028 5470 42084
rect 11554 42028 11564 42084
rect 11620 42028 12236 42084
rect 12292 42028 12302 42084
rect 14690 42028 14700 42084
rect 14756 42028 15148 42084
rect 15204 42028 15596 42084
rect 15652 42028 15662 42084
rect 16818 42028 16828 42084
rect 16884 42028 19180 42084
rect 19236 42028 19246 42084
rect 22642 42028 22652 42084
rect 22708 42028 23660 42084
rect 23716 42028 23726 42084
rect 27234 42028 27244 42084
rect 27300 42028 27310 42084
rect 28578 42028 28588 42084
rect 28644 42028 30044 42084
rect 30100 42028 30110 42084
rect 33730 42028 33740 42084
rect 33796 42028 33806 42084
rect 35522 42028 35532 42084
rect 35588 42028 39340 42084
rect 39396 42028 39406 42084
rect 33740 41972 33796 42028
rect 8194 41916 8204 41972
rect 8260 41916 8876 41972
rect 8932 41916 9436 41972
rect 9492 41916 9502 41972
rect 16706 41916 16716 41972
rect 16772 41916 20300 41972
rect 20356 41916 20366 41972
rect 22306 41916 22316 41972
rect 22372 41916 23996 41972
rect 24052 41916 24062 41972
rect 28018 41916 28028 41972
rect 28084 41916 29484 41972
rect 29540 41916 29550 41972
rect 32162 41916 32172 41972
rect 32228 41916 33796 41972
rect 38210 41916 38220 41972
rect 38276 41916 38444 41972
rect 38500 41916 38892 41972
rect 38948 41916 38958 41972
rect 44482 41916 44492 41972
rect 44548 41916 49084 41972
rect 49140 41916 49644 41972
rect 49700 41916 49710 41972
rect 52434 41916 52444 41972
rect 52500 41916 53116 41972
rect 53172 41916 53564 41972
rect 53620 41916 54796 41972
rect 54852 41916 56756 41972
rect 56700 41860 56756 41916
rect 6066 41804 6076 41860
rect 6132 41804 8764 41860
rect 8820 41804 8830 41860
rect 8978 41804 8988 41860
rect 9044 41804 10332 41860
rect 10388 41804 11900 41860
rect 11956 41804 11966 41860
rect 14130 41804 14140 41860
rect 14196 41804 14588 41860
rect 14644 41804 14654 41860
rect 15586 41804 15596 41860
rect 15652 41804 16380 41860
rect 16436 41804 19964 41860
rect 20020 41804 20030 41860
rect 23650 41804 23660 41860
rect 23716 41804 25116 41860
rect 25172 41804 25182 41860
rect 33730 41804 33740 41860
rect 33796 41804 36876 41860
rect 36932 41804 36942 41860
rect 38098 41804 38108 41860
rect 38164 41804 45724 41860
rect 45780 41804 46844 41860
rect 46900 41804 46910 41860
rect 55346 41804 55356 41860
rect 55412 41748 55468 41860
rect 56690 41804 56700 41860
rect 56756 41804 56766 41860
rect 57026 41804 57036 41860
rect 57092 41804 57102 41860
rect 57036 41748 57092 41804
rect 14466 41692 14476 41748
rect 14532 41692 15260 41748
rect 15316 41692 15326 41748
rect 16482 41692 16492 41748
rect 16548 41692 17276 41748
rect 17332 41692 20748 41748
rect 20804 41692 20814 41748
rect 28578 41692 28588 41748
rect 28644 41692 33404 41748
rect 33460 41692 33964 41748
rect 34020 41692 34030 41748
rect 34972 41692 40348 41748
rect 40404 41692 41692 41748
rect 41748 41692 41758 41748
rect 55412 41692 57092 41748
rect 15362 41580 15372 41636
rect 15428 41580 20636 41636
rect 20692 41580 20702 41636
rect 20850 41580 20860 41636
rect 20916 41580 23324 41636
rect 23380 41580 23390 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 34972 41524 35028 41692
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 15092 41468 18060 41524
rect 18116 41468 21308 41524
rect 21364 41468 21374 41524
rect 23426 41468 23436 41524
rect 23492 41468 35028 41524
rect 15092 41412 15148 41468
rect 2818 41356 2828 41412
rect 2884 41356 3276 41412
rect 3332 41356 15148 41412
rect 19506 41356 19516 41412
rect 19572 41356 20748 41412
rect 20804 41356 21196 41412
rect 21252 41356 21262 41412
rect 23762 41356 23772 41412
rect 23828 41356 25116 41412
rect 25172 41356 25182 41412
rect 27794 41356 27804 41412
rect 27860 41356 28140 41412
rect 28196 41356 30604 41412
rect 30660 41356 30670 41412
rect 34066 41356 34076 41412
rect 34132 41356 36652 41412
rect 36708 41356 36718 41412
rect 49858 41356 49868 41412
rect 49924 41356 50540 41412
rect 50596 41356 50606 41412
rect 51874 41356 51884 41412
rect 51940 41356 52892 41412
rect 52948 41356 52958 41412
rect 18386 41244 18396 41300
rect 18452 41244 18732 41300
rect 18788 41244 20524 41300
rect 20580 41244 22540 41300
rect 22596 41244 22606 41300
rect 24770 41244 24780 41300
rect 24836 41244 25564 41300
rect 25620 41244 27580 41300
rect 27636 41244 27646 41300
rect 32498 41244 32508 41300
rect 32564 41244 33628 41300
rect 33684 41244 33694 41300
rect 51986 41244 51996 41300
rect 52052 41244 52668 41300
rect 52724 41244 52734 41300
rect 8530 41132 8540 41188
rect 8596 41132 10108 41188
rect 10164 41132 10174 41188
rect 23426 41132 23436 41188
rect 23492 41132 24332 41188
rect 24388 41132 24398 41188
rect 24882 41132 24892 41188
rect 24948 41132 26012 41188
rect 26068 41132 26908 41188
rect 26964 41132 26974 41188
rect 33170 41132 33180 41188
rect 33236 41132 34524 41188
rect 34580 41132 34590 41188
rect 36082 41132 36092 41188
rect 36148 41132 37436 41188
rect 37492 41132 40348 41188
rect 40404 41132 40414 41188
rect 57250 41132 57260 41188
rect 57316 41132 57708 41188
rect 57764 41132 57774 41188
rect 11666 41020 11676 41076
rect 11732 41020 12684 41076
rect 12740 41020 13916 41076
rect 13972 41020 13982 41076
rect 19170 41020 19180 41076
rect 19236 41020 20188 41076
rect 20244 41020 20254 41076
rect 26450 41020 26460 41076
rect 26516 41020 26908 41076
rect 41122 41020 41132 41076
rect 41188 41020 42252 41076
rect 42308 41020 42318 41076
rect 42578 41020 42588 41076
rect 42644 41020 45164 41076
rect 45220 41020 45230 41076
rect 26852 40964 26908 41020
rect 5842 40908 5852 40964
rect 5908 40908 6524 40964
rect 6580 40908 12348 40964
rect 12404 40908 12414 40964
rect 14578 40908 14588 40964
rect 14644 40908 15708 40964
rect 15764 40908 15774 40964
rect 19394 40908 19404 40964
rect 19460 40908 19964 40964
rect 20020 40908 20030 40964
rect 26852 40908 27356 40964
rect 27412 40908 28140 40964
rect 28196 40908 28206 40964
rect 31892 40908 35084 40964
rect 35140 40908 35644 40964
rect 35700 40908 35710 40964
rect 50866 40908 50876 40964
rect 50932 40908 51660 40964
rect 51716 40908 51726 40964
rect 53554 40908 53564 40964
rect 53620 40908 55916 40964
rect 55972 40908 55982 40964
rect 24434 40796 24444 40852
rect 24500 40796 26572 40852
rect 26628 40796 26638 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 31892 40740 31948 40908
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 12562 40684 12572 40740
rect 12628 40684 13580 40740
rect 13636 40684 14756 40740
rect 23426 40684 23436 40740
rect 23492 40684 27804 40740
rect 27860 40684 27870 40740
rect 28018 40684 28028 40740
rect 28084 40684 31948 40740
rect 43474 40684 43484 40740
rect 43540 40684 45164 40740
rect 45220 40684 45230 40740
rect 14242 40572 14252 40628
rect 14308 40572 14644 40628
rect 12786 40460 12796 40516
rect 12852 40460 13356 40516
rect 13412 40460 14364 40516
rect 14420 40460 14430 40516
rect 7074 40348 7084 40404
rect 7140 40348 7868 40404
rect 7924 40348 8540 40404
rect 8596 40348 8606 40404
rect 13458 40348 13468 40404
rect 13524 40348 13804 40404
rect 13860 40348 14252 40404
rect 14308 40348 14318 40404
rect 4610 40236 4620 40292
rect 4676 40236 5740 40292
rect 5796 40236 5806 40292
rect 13906 40236 13916 40292
rect 13972 40236 14364 40292
rect 14420 40236 14430 40292
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 14588 39956 14644 40572
rect 14700 40516 14756 40684
rect 14914 40572 14924 40628
rect 14980 40572 15148 40628
rect 15204 40572 15214 40628
rect 26684 40572 27468 40628
rect 27524 40572 27534 40628
rect 28914 40572 28924 40628
rect 28980 40572 29708 40628
rect 29764 40572 29774 40628
rect 48178 40572 48188 40628
rect 48244 40572 56028 40628
rect 56084 40572 56094 40628
rect 26684 40516 26740 40572
rect 28924 40516 28980 40572
rect 14700 40460 17388 40516
rect 17444 40460 17454 40516
rect 18274 40460 18284 40516
rect 18340 40460 21308 40516
rect 21364 40460 21374 40516
rect 24098 40460 24108 40516
rect 24164 40460 26740 40516
rect 26796 40460 28980 40516
rect 30258 40460 30268 40516
rect 30324 40460 31164 40516
rect 31220 40460 34972 40516
rect 35028 40460 35644 40516
rect 35700 40460 35710 40516
rect 51650 40460 51660 40516
rect 51716 40460 53116 40516
rect 53172 40460 53182 40516
rect 55906 40460 55916 40516
rect 55972 40460 56700 40516
rect 56756 40460 56766 40516
rect 14924 40404 14980 40460
rect 26796 40404 26852 40460
rect 14802 40348 14812 40404
rect 14868 40348 14980 40404
rect 17266 40348 17276 40404
rect 17332 40348 17948 40404
rect 18004 40348 19404 40404
rect 19460 40348 20132 40404
rect 20290 40348 20300 40404
rect 20356 40348 21868 40404
rect 21924 40348 21934 40404
rect 22978 40348 22988 40404
rect 23044 40348 23772 40404
rect 23828 40348 23838 40404
rect 23986 40348 23996 40404
rect 24052 40348 26852 40404
rect 27570 40348 27580 40404
rect 27636 40348 29372 40404
rect 29428 40348 29438 40404
rect 40226 40348 40236 40404
rect 40292 40348 41244 40404
rect 41300 40348 41468 40404
rect 41524 40348 41534 40404
rect 41682 40348 41692 40404
rect 41748 40348 42140 40404
rect 42196 40348 42206 40404
rect 49186 40348 49196 40404
rect 49252 40348 50316 40404
rect 50372 40348 53676 40404
rect 53732 40348 53742 40404
rect 54002 40348 54012 40404
rect 54068 40348 56924 40404
rect 56980 40348 56990 40404
rect 20076 40292 20132 40348
rect 15362 40236 15372 40292
rect 15428 40236 16940 40292
rect 16996 40236 17006 40292
rect 20076 40236 20412 40292
rect 20468 40236 20478 40292
rect 47730 40236 47740 40292
rect 47796 40236 48076 40292
rect 48132 40236 48142 40292
rect 56018 40236 56028 40292
rect 56084 40236 57036 40292
rect 57092 40236 57102 40292
rect 16594 40124 16604 40180
rect 16660 40124 18844 40180
rect 18900 40124 18910 40180
rect 43810 40124 43820 40180
rect 43876 40124 47404 40180
rect 47460 40124 47470 40180
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 14578 39900 14588 39956
rect 14644 39900 14654 39956
rect 14802 39900 14812 39956
rect 14868 39900 14924 39956
rect 14980 39900 14990 39956
rect 15092 39900 28588 39956
rect 28644 39900 28654 39956
rect 15092 39844 15148 39900
rect 4162 39788 4172 39844
rect 4228 39788 5628 39844
rect 5684 39788 5694 39844
rect 12786 39788 12796 39844
rect 12852 39788 15148 39844
rect 20626 39788 20636 39844
rect 20692 39788 21084 39844
rect 21140 39788 21150 39844
rect 44706 39788 44716 39844
rect 44772 39788 45836 39844
rect 45892 39788 45902 39844
rect 3826 39676 3836 39732
rect 3892 39676 4396 39732
rect 4452 39676 4462 39732
rect 4610 39676 4620 39732
rect 4676 39676 6188 39732
rect 6244 39676 6254 39732
rect 17714 39676 17724 39732
rect 17780 39676 18732 39732
rect 18788 39676 18798 39732
rect 22642 39676 22652 39732
rect 22708 39676 23436 39732
rect 23492 39676 25004 39732
rect 25060 39676 26124 39732
rect 26180 39676 26190 39732
rect 35186 39676 35196 39732
rect 35252 39676 37100 39732
rect 37156 39676 37166 39732
rect 3154 39564 3164 39620
rect 3220 39564 3948 39620
rect 4004 39564 4014 39620
rect 14242 39564 14252 39620
rect 14308 39564 15148 39620
rect 15204 39564 15932 39620
rect 15988 39564 15998 39620
rect 20178 39564 20188 39620
rect 20244 39564 21196 39620
rect 21252 39564 21262 39620
rect 25554 39564 25564 39620
rect 25620 39564 26460 39620
rect 26516 39564 26526 39620
rect 38098 39564 38108 39620
rect 38164 39564 43372 39620
rect 43428 39564 43438 39620
rect 56578 39564 56588 39620
rect 56644 39564 57036 39620
rect 57092 39564 57102 39620
rect 19618 39452 19628 39508
rect 19684 39452 21308 39508
rect 21364 39452 21374 39508
rect 39778 39452 39788 39508
rect 39844 39452 41692 39508
rect 41748 39452 41758 39508
rect 44258 39452 44268 39508
rect 44324 39452 45052 39508
rect 45108 39452 45724 39508
rect 45780 39452 45790 39508
rect 55412 39452 56364 39508
rect 56420 39452 56812 39508
rect 56868 39452 56878 39508
rect 24210 39340 24220 39396
rect 24276 39340 27468 39396
rect 27524 39340 27916 39396
rect 27972 39340 27982 39396
rect 30818 39340 30828 39396
rect 30884 39340 31612 39396
rect 31668 39340 31678 39396
rect 42242 39228 42252 39284
rect 42308 39228 48860 39284
rect 48916 39228 48926 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 8530 39116 8540 39172
rect 8596 39116 15148 39172
rect 24770 39116 24780 39172
rect 24836 39116 26908 39172
rect 26964 39116 26974 39172
rect 15092 39060 15148 39116
rect 55412 39060 55468 39452
rect 6178 39004 6188 39060
rect 6244 39004 6860 39060
rect 6916 39004 6926 39060
rect 12114 39004 12124 39060
rect 12180 39004 12796 39060
rect 12852 39004 12862 39060
rect 15092 39004 15652 39060
rect 15810 39004 15820 39060
rect 15876 39004 16716 39060
rect 16772 39004 19628 39060
rect 19684 39004 19694 39060
rect 26674 39004 26684 39060
rect 26740 39004 27692 39060
rect 27748 39004 27758 39060
rect 30034 39004 30044 39060
rect 30100 39004 30828 39060
rect 30884 39004 32060 39060
rect 32116 39004 32126 39060
rect 54114 39004 54124 39060
rect 54180 39004 55468 39060
rect 15596 38948 15652 39004
rect 11442 38892 11452 38948
rect 11508 38892 12684 38948
rect 12740 38892 12750 38948
rect 14130 38892 14140 38948
rect 14196 38892 15260 38948
rect 15316 38892 15326 38948
rect 15596 38892 20300 38948
rect 20356 38892 20366 38948
rect 23650 38892 23660 38948
rect 23716 38892 24444 38948
rect 24500 38892 26236 38948
rect 26292 38892 26302 38948
rect 26562 38892 26572 38948
rect 26628 38892 37548 38948
rect 37604 38892 37996 38948
rect 38052 38892 38062 38948
rect 5842 38780 5852 38836
rect 5908 38780 6636 38836
rect 6692 38780 7868 38836
rect 7924 38780 12236 38836
rect 12292 38780 12302 38836
rect 12450 38780 12460 38836
rect 12516 38780 12526 38836
rect 21298 38780 21308 38836
rect 21364 38780 21756 38836
rect 21812 38780 21822 38836
rect 24546 38780 24556 38836
rect 24612 38780 25676 38836
rect 25732 38780 25742 38836
rect 26002 38780 26012 38836
rect 26068 38780 28028 38836
rect 28084 38780 28094 38836
rect 12460 38724 12516 38780
rect 4386 38668 4396 38724
rect 4452 38668 7420 38724
rect 7476 38668 7486 38724
rect 9874 38668 9884 38724
rect 9940 38668 11564 38724
rect 11620 38668 12516 38724
rect 12786 38668 12796 38724
rect 12852 38668 13468 38724
rect 13524 38668 19740 38724
rect 19796 38668 19806 38724
rect 23874 38668 23884 38724
rect 23940 38668 26908 38724
rect 26964 38668 26974 38724
rect 29922 38668 29932 38724
rect 29988 38668 34748 38724
rect 34804 38668 34814 38724
rect 37090 38668 37100 38724
rect 37156 38668 46060 38724
rect 46116 38668 46172 38724
rect 46228 38668 46238 38724
rect 49410 38668 49420 38724
rect 49476 38668 53676 38724
rect 53732 38668 53742 38724
rect 57586 38668 57596 38724
rect 57652 38668 58156 38724
rect 58212 38668 58222 38724
rect 6402 38556 6412 38612
rect 6468 38556 7084 38612
rect 7140 38556 7980 38612
rect 8036 38556 8046 38612
rect 12338 38556 12348 38612
rect 12404 38556 15372 38612
rect 15428 38556 15438 38612
rect 22418 38556 22428 38612
rect 22484 38556 23212 38612
rect 23268 38556 23278 38612
rect 23986 38556 23996 38612
rect 24052 38556 24220 38612
rect 24276 38556 24286 38612
rect 26114 38556 26124 38612
rect 26180 38556 27356 38612
rect 27412 38556 29260 38612
rect 29316 38556 29326 38612
rect 30818 38556 30828 38612
rect 30884 38556 35532 38612
rect 35588 38556 35598 38612
rect 39666 38556 39676 38612
rect 39732 38556 40236 38612
rect 40292 38556 40302 38612
rect 58146 38556 58156 38612
rect 58212 38556 58222 38612
rect 31938 38444 31948 38500
rect 32004 38444 34076 38500
rect 34132 38444 34142 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 58156 38388 58212 38556
rect 59200 38388 60000 38416
rect 15362 38332 15372 38388
rect 15428 38332 16492 38388
rect 16548 38332 19404 38388
rect 19460 38332 21532 38388
rect 21588 38332 21598 38388
rect 58156 38332 60000 38388
rect 59200 38304 60000 38332
rect 19618 38220 19628 38276
rect 19684 38220 21420 38276
rect 21476 38220 21486 38276
rect 21858 38220 21868 38276
rect 21924 38220 22652 38276
rect 22708 38220 22718 38276
rect 16482 38108 16492 38164
rect 16548 38108 17948 38164
rect 18004 38108 18014 38164
rect 18834 38108 18844 38164
rect 18900 38108 21308 38164
rect 21364 38108 21374 38164
rect 24882 38108 24892 38164
rect 24948 38108 27020 38164
rect 27076 38108 27086 38164
rect 36306 38108 36316 38164
rect 36372 38108 37324 38164
rect 37380 38108 37390 38164
rect 37874 38108 37884 38164
rect 37940 38108 38780 38164
rect 38836 38108 38846 38164
rect 45714 38108 45724 38164
rect 45780 38108 46396 38164
rect 46452 38108 46462 38164
rect 4050 37996 4060 38052
rect 4116 37996 11004 38052
rect 11060 37996 11070 38052
rect 15698 37996 15708 38052
rect 15764 37996 17612 38052
rect 17668 37996 17678 38052
rect 20178 37996 20188 38052
rect 20244 37996 20254 38052
rect 24098 37996 24108 38052
rect 24164 37996 25340 38052
rect 25396 37996 25406 38052
rect 26562 37996 26572 38052
rect 26628 37996 27468 38052
rect 27524 37996 28588 38052
rect 28644 37996 29148 38052
rect 29204 37996 29214 38052
rect 35298 37996 35308 38052
rect 35364 37996 36988 38052
rect 37044 37996 37054 38052
rect 46022 37996 46060 38052
rect 46116 37996 46126 38052
rect 54898 37996 54908 38052
rect 54964 37996 55356 38052
rect 55412 37996 56700 38052
rect 56756 37996 56766 38052
rect 14690 37884 14700 37940
rect 14756 37884 17052 37940
rect 17108 37884 17118 37940
rect 20188 37828 20244 37996
rect 20962 37884 20972 37940
rect 21028 37884 22092 37940
rect 22148 37884 22158 37940
rect 23090 37884 23100 37940
rect 23156 37884 23996 37940
rect 24052 37884 24062 37940
rect 24210 37884 24220 37940
rect 24276 37884 24556 37940
rect 24612 37884 24622 37940
rect 27570 37884 27580 37940
rect 27636 37884 28140 37940
rect 28196 37884 29260 37940
rect 29316 37884 29326 37940
rect 30594 37884 30604 37940
rect 30660 37884 31500 37940
rect 31556 37884 31566 37940
rect 33954 37884 33964 37940
rect 34020 37884 35980 37940
rect 36036 37884 38668 37940
rect 38724 37884 38734 37940
rect 46498 37884 46508 37940
rect 46564 37884 48524 37940
rect 48580 37884 48590 37940
rect 15026 37772 15036 37828
rect 15092 37772 20244 37828
rect 20626 37772 20636 37828
rect 20692 37772 21644 37828
rect 21700 37772 21710 37828
rect 26002 37772 26012 37828
rect 26068 37772 28364 37828
rect 28420 37772 28430 37828
rect 33058 37772 33068 37828
rect 33124 37772 36204 37828
rect 36260 37772 36270 37828
rect 14018 37660 14028 37716
rect 14084 37660 15148 37716
rect 16818 37660 16828 37716
rect 16884 37660 17500 37716
rect 17556 37660 18396 37716
rect 18452 37660 18462 37716
rect 15092 37604 15148 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 2706 37548 2716 37604
rect 2772 37548 3612 37604
rect 3668 37548 3678 37604
rect 15092 37548 15932 37604
rect 15988 37548 18620 37604
rect 18676 37548 18686 37604
rect 33954 37548 33964 37604
rect 34020 37548 35532 37604
rect 35588 37548 37772 37604
rect 37828 37548 37838 37604
rect 1810 37436 1820 37492
rect 1876 37436 4620 37492
rect 4676 37436 5068 37492
rect 5124 37436 7868 37492
rect 7924 37436 7934 37492
rect 8978 37436 8988 37492
rect 9044 37436 9436 37492
rect 9492 37436 9996 37492
rect 10052 37436 10062 37492
rect 16706 37436 16716 37492
rect 16772 37436 18508 37492
rect 18564 37436 18574 37492
rect 25330 37436 25340 37492
rect 25396 37436 27580 37492
rect 27636 37436 27646 37492
rect 31266 37436 31276 37492
rect 31332 37436 37100 37492
rect 37156 37436 37166 37492
rect 3042 37324 3052 37380
rect 3108 37324 3948 37380
rect 4004 37324 4014 37380
rect 8418 37324 8428 37380
rect 8484 37324 9548 37380
rect 9604 37324 11340 37380
rect 11396 37324 12460 37380
rect 12516 37324 12526 37380
rect 26114 37324 26124 37380
rect 26180 37324 27132 37380
rect 27188 37324 27198 37380
rect 34626 37324 34636 37380
rect 34692 37324 35756 37380
rect 35812 37324 35822 37380
rect 38770 37324 38780 37380
rect 38836 37324 39564 37380
rect 39620 37324 39630 37380
rect 3154 37212 3164 37268
rect 3220 37212 3724 37268
rect 3780 37212 3790 37268
rect 10994 37212 11004 37268
rect 11060 37212 11900 37268
rect 11956 37212 11966 37268
rect 14914 37212 14924 37268
rect 14980 37212 16604 37268
rect 16660 37212 16670 37268
rect 17714 37212 17724 37268
rect 17780 37212 20300 37268
rect 20356 37212 21196 37268
rect 21252 37212 21262 37268
rect 24546 37212 24556 37268
rect 24612 37212 24892 37268
rect 24948 37212 24958 37268
rect 26786 37212 26796 37268
rect 26852 37212 29260 37268
rect 29316 37212 29326 37268
rect 30258 37212 30268 37268
rect 30324 37212 33068 37268
rect 33124 37212 33134 37268
rect 33394 37212 33404 37268
rect 33460 37212 34300 37268
rect 34356 37212 35644 37268
rect 35700 37212 35710 37268
rect 36194 37212 36204 37268
rect 36260 37212 36652 37268
rect 36708 37212 36718 37268
rect 41794 37212 41804 37268
rect 41860 37212 46172 37268
rect 46228 37212 46238 37268
rect 20402 37100 20412 37156
rect 20468 37100 20972 37156
rect 21028 37100 21038 37156
rect 22866 37100 22876 37156
rect 22932 37100 23884 37156
rect 23940 37100 25228 37156
rect 25284 37100 25294 37156
rect 31490 37100 31500 37156
rect 31556 37100 34076 37156
rect 34132 37100 34142 37156
rect 39218 37100 39228 37156
rect 39284 37100 39676 37156
rect 39732 37100 40908 37156
rect 40964 37100 40974 37156
rect 41234 37100 41244 37156
rect 41300 37100 43036 37156
rect 43092 37100 43102 37156
rect 7970 36988 7980 37044
rect 8036 36988 9660 37044
rect 9716 36988 9726 37044
rect 15138 36988 15148 37044
rect 15204 36988 20636 37044
rect 20692 36988 20702 37044
rect 32610 36988 32620 37044
rect 32676 36988 33628 37044
rect 33684 36988 33694 37044
rect 33852 36988 34412 37044
rect 34468 36988 36092 37044
rect 36148 36988 36158 37044
rect 45826 36988 45836 37044
rect 45892 36988 54012 37044
rect 54068 36988 54078 37044
rect 33852 36932 33908 36988
rect 22194 36876 22204 36932
rect 22260 36876 22876 36932
rect 22932 36876 23660 36932
rect 23716 36876 23726 36932
rect 33394 36876 33404 36932
rect 33460 36876 33908 36932
rect 35532 36876 35756 36932
rect 35812 36876 42700 36932
rect 42756 36876 42766 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 35532 36708 35588 36876
rect 36194 36764 36204 36820
rect 36260 36764 37100 36820
rect 37156 36764 37166 36820
rect 30940 36652 35588 36708
rect 36866 36652 36876 36708
rect 36932 36652 37548 36708
rect 37604 36652 37614 36708
rect 38612 36652 52332 36708
rect 52388 36652 52398 36708
rect 8194 36428 8204 36484
rect 8260 36428 8764 36484
rect 8820 36428 8830 36484
rect 12786 36428 12796 36484
rect 12852 36428 13468 36484
rect 13524 36428 13534 36484
rect 18274 36428 18284 36484
rect 18340 36428 20300 36484
rect 20356 36428 20366 36484
rect 22754 36428 22764 36484
rect 22820 36428 23324 36484
rect 23380 36428 27020 36484
rect 27076 36428 27086 36484
rect 8764 36316 11564 36372
rect 11620 36316 12236 36372
rect 12292 36316 12302 36372
rect 24322 36316 24332 36372
rect 24388 36316 26908 36372
rect 26964 36316 26974 36372
rect 8764 36260 8820 36316
rect 30940 36260 30996 36652
rect 33282 36540 33292 36596
rect 33348 36540 35196 36596
rect 35252 36540 35262 36596
rect 35410 36428 35420 36484
rect 35476 36428 37212 36484
rect 37268 36428 38332 36484
rect 38388 36428 38398 36484
rect 8418 36204 8428 36260
rect 8484 36204 8764 36260
rect 8820 36204 8830 36260
rect 10770 36204 10780 36260
rect 10836 36204 12684 36260
rect 12740 36204 12750 36260
rect 20738 36204 20748 36260
rect 20804 36204 21308 36260
rect 21364 36204 30996 36260
rect 31154 36204 31164 36260
rect 31220 36204 32060 36260
rect 32116 36204 32126 36260
rect 38612 36148 38668 36652
rect 9762 36092 9772 36148
rect 9828 36092 11004 36148
rect 11060 36092 11070 36148
rect 30146 36092 30156 36148
rect 30212 36092 38668 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 8866 35980 8876 36036
rect 8932 35980 9996 36036
rect 10052 35980 10062 36036
rect 10546 35868 10556 35924
rect 10612 35868 13580 35924
rect 13636 35868 13646 35924
rect 24210 35868 24220 35924
rect 24276 35868 25340 35924
rect 25396 35868 26012 35924
rect 26068 35868 26078 35924
rect 36530 35868 36540 35924
rect 36596 35868 37324 35924
rect 37380 35868 37390 35924
rect 38322 35868 38332 35924
rect 38388 35868 39004 35924
rect 39060 35868 39070 35924
rect 56914 35868 56924 35924
rect 56980 35868 57708 35924
rect 57764 35868 57774 35924
rect 2258 35756 2268 35812
rect 2324 35756 20748 35812
rect 20804 35756 20814 35812
rect 35186 35756 35196 35812
rect 35252 35756 36316 35812
rect 36372 35756 36382 35812
rect 7858 35644 7868 35700
rect 7924 35644 12572 35700
rect 12628 35644 12638 35700
rect 15698 35644 15708 35700
rect 15764 35644 17388 35700
rect 17444 35644 18508 35700
rect 18564 35644 18574 35700
rect 18834 35644 18844 35700
rect 18900 35644 19964 35700
rect 20020 35644 20030 35700
rect 21634 35644 21644 35700
rect 21700 35644 22540 35700
rect 22596 35644 22988 35700
rect 23044 35644 23054 35700
rect 29698 35644 29708 35700
rect 29764 35644 30492 35700
rect 30548 35644 30558 35700
rect 35522 35644 35532 35700
rect 35588 35644 35980 35700
rect 36036 35644 37436 35700
rect 37492 35644 37502 35700
rect 37986 35644 37996 35700
rect 38052 35644 39116 35700
rect 39172 35644 39182 35700
rect 42466 35644 42476 35700
rect 42532 35644 45500 35700
rect 45556 35644 45566 35700
rect 57026 35644 57036 35700
rect 57092 35644 57932 35700
rect 57988 35644 57998 35700
rect 10994 35532 11004 35588
rect 11060 35532 13580 35588
rect 13636 35532 13804 35588
rect 13860 35532 13870 35588
rect 14354 35532 14364 35588
rect 14420 35532 16044 35588
rect 16100 35532 16110 35588
rect 25442 35532 25452 35588
rect 25508 35532 27356 35588
rect 27412 35532 27422 35588
rect 31154 35532 31164 35588
rect 31220 35532 34188 35588
rect 34244 35532 34254 35588
rect 34962 35532 34972 35588
rect 35028 35532 36428 35588
rect 36484 35532 38108 35588
rect 38164 35532 38556 35588
rect 38612 35532 38622 35588
rect 55570 35532 55580 35588
rect 55636 35532 57148 35588
rect 57204 35532 57214 35588
rect 34188 35476 34244 35532
rect 8082 35420 8092 35476
rect 8148 35420 11340 35476
rect 11396 35420 11406 35476
rect 17042 35420 17052 35476
rect 17108 35420 21644 35476
rect 21700 35420 21710 35476
rect 34188 35420 36652 35476
rect 36708 35420 38220 35476
rect 38276 35420 38286 35476
rect 50306 35420 50316 35476
rect 50372 35420 51772 35476
rect 51828 35420 53116 35476
rect 53172 35420 53182 35476
rect 10210 35308 10220 35364
rect 10276 35308 12348 35364
rect 12404 35308 12414 35364
rect 23314 35308 23324 35364
rect 23380 35308 25676 35364
rect 25732 35308 25742 35364
rect 33282 35308 33292 35364
rect 33348 35308 34972 35364
rect 35028 35308 35038 35364
rect 36194 35308 36204 35364
rect 36260 35308 36988 35364
rect 37044 35308 37054 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 29586 35196 29596 35252
rect 29652 35196 31500 35252
rect 31556 35196 31566 35252
rect 40114 35196 40124 35252
rect 40180 35196 42588 35252
rect 42644 35196 42654 35252
rect 43698 35196 43708 35252
rect 43764 35196 44716 35252
rect 44772 35196 45500 35252
rect 45556 35196 45566 35252
rect 47730 35196 47740 35252
rect 47796 35196 50876 35252
rect 50932 35196 50942 35252
rect 10434 35084 10444 35140
rect 10500 35084 12796 35140
rect 12852 35084 14252 35140
rect 14308 35084 14318 35140
rect 0 35028 800 35056
rect 0 34972 1820 35028
rect 1876 34972 1886 35028
rect 28354 34972 28364 35028
rect 28420 34972 29148 35028
rect 29204 34972 29214 35028
rect 30930 34972 30940 35028
rect 30996 34972 31612 35028
rect 31668 34972 34748 35028
rect 34804 34972 35756 35028
rect 35812 34972 35822 35028
rect 38770 34972 38780 35028
rect 38836 34972 39340 35028
rect 39396 34972 40796 35028
rect 40852 34972 41244 35028
rect 41300 34972 41310 35028
rect 48850 34972 48860 35028
rect 48916 34972 49756 35028
rect 49812 34972 49822 35028
rect 0 34944 800 34972
rect 5842 34860 5852 34916
rect 5908 34860 29932 34916
rect 29988 34860 30268 34916
rect 30324 34860 30334 34916
rect 33842 34860 33852 34916
rect 33908 34860 34972 34916
rect 35028 34860 35038 34916
rect 36194 34860 36204 34916
rect 36260 34860 37884 34916
rect 37940 34860 37950 34916
rect 42354 34860 42364 34916
rect 42420 34860 43932 34916
rect 43988 34860 44268 34916
rect 44324 34860 44334 34916
rect 7522 34748 7532 34804
rect 7588 34748 10780 34804
rect 10836 34748 10846 34804
rect 29810 34748 29820 34804
rect 29876 34748 30716 34804
rect 30772 34748 30782 34804
rect 31042 34748 31052 34804
rect 31108 34748 35084 34804
rect 35140 34748 35150 34804
rect 39106 34748 39116 34804
rect 39172 34748 49420 34804
rect 49476 34748 49486 34804
rect 56242 34748 56252 34804
rect 56308 34748 57036 34804
rect 57092 34748 57102 34804
rect 15138 34636 15148 34692
rect 15204 34636 15820 34692
rect 15876 34636 16268 34692
rect 16324 34636 17948 34692
rect 18004 34636 18014 34692
rect 29586 34636 29596 34692
rect 29652 34636 30268 34692
rect 30324 34636 30334 34692
rect 37202 34636 37212 34692
rect 37268 34636 37660 34692
rect 37716 34636 37726 34692
rect 38658 34636 38668 34692
rect 38724 34636 39340 34692
rect 39396 34636 39406 34692
rect 53442 34636 53452 34692
rect 53508 34636 54012 34692
rect 54068 34636 55804 34692
rect 55860 34636 57260 34692
rect 57316 34636 57596 34692
rect 57652 34636 57662 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 38668 34356 38724 34636
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 40226 34412 40236 34468
rect 40292 34412 42700 34468
rect 42756 34412 43596 34468
rect 43652 34412 44492 34468
rect 44548 34412 44558 34468
rect 27906 34300 27916 34356
rect 27972 34300 38724 34356
rect 41458 34300 41468 34356
rect 41524 34300 42364 34356
rect 42420 34300 42430 34356
rect 47282 34300 47292 34356
rect 47348 34300 48188 34356
rect 48244 34300 48254 34356
rect 26852 34188 40124 34244
rect 40180 34188 40190 34244
rect 55010 34188 55020 34244
rect 55076 34188 56252 34244
rect 56308 34188 56318 34244
rect 21084 34076 21420 34132
rect 21476 34076 21486 34132
rect 21084 34020 21140 34076
rect 26852 34020 26908 34188
rect 30258 34076 30268 34132
rect 30324 34076 30940 34132
rect 30996 34076 31006 34132
rect 31826 34076 31836 34132
rect 31892 34076 33628 34132
rect 33684 34076 33694 34132
rect 36082 34076 36092 34132
rect 36148 34076 37100 34132
rect 37156 34076 37166 34132
rect 39218 34076 39228 34132
rect 39284 34076 39676 34132
rect 39732 34076 40460 34132
rect 40516 34076 40526 34132
rect 41234 34076 41244 34132
rect 41300 34076 42028 34132
rect 42084 34076 42094 34132
rect 44594 34076 44604 34132
rect 44660 34076 45052 34132
rect 45108 34076 45724 34132
rect 45780 34076 45790 34132
rect 15474 33964 15484 34020
rect 15540 33964 19180 34020
rect 19236 33964 21140 34020
rect 21298 33964 21308 34020
rect 21364 33964 26908 34020
rect 34860 33964 36652 34020
rect 36708 33964 37660 34020
rect 37716 33964 37726 34020
rect 34860 33908 34916 33964
rect 7410 33852 7420 33908
rect 7476 33852 7980 33908
rect 8036 33852 9884 33908
rect 9940 33852 9950 33908
rect 31826 33852 31836 33908
rect 31892 33852 34916 33908
rect 35074 33852 35084 33908
rect 35140 33852 36092 33908
rect 36148 33852 36158 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 28354 33628 28364 33684
rect 28420 33628 28812 33684
rect 28868 33628 28878 33684
rect 9538 33516 9548 33572
rect 9604 33516 10220 33572
rect 10276 33516 10286 33572
rect 13010 33516 13020 33572
rect 13076 33516 13916 33572
rect 13972 33516 15148 33572
rect 15204 33516 15214 33572
rect 22754 33516 22764 33572
rect 22820 33516 23548 33572
rect 23604 33516 23614 33572
rect 34850 33516 34860 33572
rect 34916 33516 37548 33572
rect 37604 33516 37614 33572
rect 38098 33516 38108 33572
rect 38164 33516 45948 33572
rect 46004 33516 46014 33572
rect 12450 33404 12460 33460
rect 12516 33404 14588 33460
rect 14644 33404 14654 33460
rect 15810 33404 15820 33460
rect 15876 33404 16716 33460
rect 16772 33404 16782 33460
rect 22530 33404 22540 33460
rect 22596 33404 25116 33460
rect 25172 33404 25182 33460
rect 12786 33292 12796 33348
rect 12852 33292 14812 33348
rect 14868 33292 14878 33348
rect 28130 33292 28140 33348
rect 28196 33292 28924 33348
rect 28980 33292 38892 33348
rect 38948 33292 38958 33348
rect 51874 33292 51884 33348
rect 51940 33292 53788 33348
rect 53844 33292 53854 33348
rect 55010 33292 55020 33348
rect 55076 33292 57484 33348
rect 57540 33292 57550 33348
rect 11442 33180 11452 33236
rect 11508 33180 13468 33236
rect 13524 33180 13534 33236
rect 16706 33180 16716 33236
rect 16772 33180 18620 33236
rect 18676 33180 18686 33236
rect 22054 33180 22092 33236
rect 22148 33180 22158 33236
rect 25778 33180 25788 33236
rect 25844 33180 27468 33236
rect 27524 33180 27534 33236
rect 30370 33180 30380 33236
rect 30436 33180 34524 33236
rect 34580 33180 34590 33236
rect 41794 33180 41804 33236
rect 41860 33180 42364 33236
rect 42420 33180 43372 33236
rect 43428 33180 43438 33236
rect 51986 33180 51996 33236
rect 52052 33180 53452 33236
rect 53508 33180 53518 33236
rect 19058 33068 19068 33124
rect 19124 33068 20076 33124
rect 20132 33068 20142 33124
rect 21410 33068 21420 33124
rect 21476 33068 23884 33124
rect 23940 33068 24668 33124
rect 24724 33068 24734 33124
rect 27794 33068 27804 33124
rect 27860 33068 28700 33124
rect 28756 33068 29372 33124
rect 29428 33068 29438 33124
rect 57026 33068 57036 33124
rect 57092 33068 57596 33124
rect 57652 33068 57662 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 11890 32732 11900 32788
rect 11956 32732 12796 32788
rect 12852 32732 12862 32788
rect 16818 32732 16828 32788
rect 16884 32732 17612 32788
rect 17668 32732 17678 32788
rect 18162 32732 18172 32788
rect 18228 32732 19404 32788
rect 19460 32732 19470 32788
rect 32162 32732 32172 32788
rect 32228 32732 33180 32788
rect 33236 32732 34748 32788
rect 34804 32732 35084 32788
rect 35140 32732 35150 32788
rect 53890 32732 53900 32788
rect 53956 32732 54908 32788
rect 54964 32732 55580 32788
rect 55636 32732 55646 32788
rect 13906 32620 13916 32676
rect 13972 32620 14588 32676
rect 14644 32620 14654 32676
rect 18834 32620 18844 32676
rect 18900 32620 19964 32676
rect 20020 32620 20030 32676
rect 31826 32620 31836 32676
rect 31892 32620 32284 32676
rect 32340 32620 32350 32676
rect 40450 32620 40460 32676
rect 40516 32620 41804 32676
rect 41860 32620 41870 32676
rect 52210 32620 52220 32676
rect 52276 32620 52668 32676
rect 52724 32620 54796 32676
rect 54852 32620 54862 32676
rect 7970 32508 7980 32564
rect 8036 32508 10332 32564
rect 10388 32508 10398 32564
rect 18498 32508 18508 32564
rect 18564 32508 19628 32564
rect 19684 32508 19694 32564
rect 37202 32508 37212 32564
rect 37268 32508 37996 32564
rect 38052 32508 40908 32564
rect 40964 32508 40974 32564
rect 41906 32508 41916 32564
rect 41972 32508 42252 32564
rect 42308 32508 42318 32564
rect 42700 32508 46732 32564
rect 46788 32508 46798 32564
rect 47394 32508 47404 32564
rect 47460 32508 48972 32564
rect 49028 32508 49038 32564
rect 49634 32508 49644 32564
rect 49700 32508 50428 32564
rect 50484 32508 50494 32564
rect 42700 32452 42756 32508
rect 11554 32396 11564 32452
rect 11620 32396 12236 32452
rect 12292 32396 14028 32452
rect 14084 32396 14094 32452
rect 37090 32396 37100 32452
rect 37156 32396 37660 32452
rect 37716 32396 42756 32452
rect 43586 32396 43596 32452
rect 43652 32396 44044 32452
rect 44100 32396 44110 32452
rect 13682 32284 13692 32340
rect 13748 32284 14812 32340
rect 14868 32284 14878 32340
rect 34850 32284 34860 32340
rect 34916 32284 37212 32340
rect 37268 32284 37278 32340
rect 39554 32284 39564 32340
rect 39620 32284 42028 32340
rect 42084 32284 42094 32340
rect 42242 32284 42252 32340
rect 42308 32284 42588 32340
rect 42644 32284 42654 32340
rect 12002 32172 12012 32228
rect 12068 32172 20636 32228
rect 20692 32172 20702 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 9202 32060 9212 32116
rect 9268 32060 10444 32116
rect 10500 32060 15372 32116
rect 15428 32060 15438 32116
rect 32274 32060 32284 32116
rect 32340 32060 34636 32116
rect 34692 32060 34702 32116
rect 51426 32060 51436 32116
rect 51492 32060 52780 32116
rect 52836 32060 55244 32116
rect 55300 32060 56028 32116
rect 56084 32060 58156 32116
rect 58212 32060 58222 32116
rect 34636 32004 34692 32060
rect 19842 31948 19852 32004
rect 19908 31948 21084 32004
rect 21140 31948 21150 32004
rect 34636 31948 36988 32004
rect 37044 31948 37054 32004
rect 7298 31836 7308 31892
rect 7364 31836 7868 31892
rect 7924 31836 7934 31892
rect 8642 31836 8652 31892
rect 8708 31836 9772 31892
rect 9828 31836 9838 31892
rect 12786 31836 12796 31892
rect 12852 31836 12862 31892
rect 14214 31836 14252 31892
rect 14308 31836 14318 31892
rect 17378 31836 17388 31892
rect 17444 31836 18620 31892
rect 18676 31836 18686 31892
rect 24098 31836 24108 31892
rect 24164 31836 26796 31892
rect 26852 31836 26862 31892
rect 30818 31836 30828 31892
rect 30884 31836 31276 31892
rect 31332 31836 32508 31892
rect 32564 31836 33852 31892
rect 33908 31836 33918 31892
rect 35186 31836 35196 31892
rect 35252 31836 37772 31892
rect 37828 31836 37838 31892
rect 38210 31836 38220 31892
rect 38276 31836 41468 31892
rect 41524 31836 45388 31892
rect 45444 31836 45454 31892
rect 50082 31836 50092 31892
rect 50148 31836 50876 31892
rect 50932 31836 51772 31892
rect 51828 31836 51838 31892
rect 12796 31332 12852 31836
rect 13570 31724 13580 31780
rect 13636 31724 14140 31780
rect 14196 31724 14206 31780
rect 18274 31724 18284 31780
rect 18340 31724 19404 31780
rect 19460 31724 20300 31780
rect 20356 31724 20366 31780
rect 32946 31724 32956 31780
rect 33012 31724 34524 31780
rect 34580 31724 34590 31780
rect 35410 31724 35420 31780
rect 35476 31724 37436 31780
rect 37492 31724 37884 31780
rect 37940 31724 38444 31780
rect 38500 31724 38510 31780
rect 44258 31724 44268 31780
rect 44324 31724 45164 31780
rect 45220 31724 45230 31780
rect 49298 31724 49308 31780
rect 49364 31724 50428 31780
rect 50484 31724 50494 31780
rect 28802 31612 28812 31668
rect 28868 31612 30604 31668
rect 30660 31612 35196 31668
rect 35252 31612 35262 31668
rect 47506 31612 47516 31668
rect 47572 31612 49420 31668
rect 49476 31612 49486 31668
rect 15026 31500 15036 31556
rect 15092 31500 15484 31556
rect 15540 31500 15550 31556
rect 34514 31500 34524 31556
rect 34580 31500 35084 31556
rect 35140 31500 36204 31556
rect 36260 31500 37100 31556
rect 37156 31500 48972 31556
rect 49028 31500 49532 31556
rect 49588 31500 49598 31556
rect 50754 31500 50764 31556
rect 50820 31500 53116 31556
rect 53172 31500 53182 31556
rect 59200 31444 60000 31472
rect 58146 31388 58156 31444
rect 58212 31388 60000 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 59200 31360 60000 31388
rect 7858 31276 7868 31332
rect 7924 31276 8428 31332
rect 12796 31276 13580 31332
rect 13636 31276 14476 31332
rect 14532 31276 14542 31332
rect 8372 30996 8428 31276
rect 21970 31164 21980 31220
rect 22036 31164 22540 31220
rect 22596 31164 22606 31220
rect 22082 31052 22092 31108
rect 22148 31052 22158 31108
rect 50372 31052 57820 31108
rect 57876 31052 57886 31108
rect 8372 30940 12908 30996
rect 12964 30940 13916 30996
rect 13972 30940 13982 30996
rect 22092 30884 22148 31052
rect 22866 30940 22876 30996
rect 22932 30940 23436 30996
rect 23492 30940 23996 30996
rect 24052 30940 24062 30996
rect 50372 30884 50428 31052
rect 55346 30940 55356 30996
rect 55412 30940 56588 30996
rect 56644 30940 56924 30996
rect 56980 30940 56990 30996
rect 11330 30828 11340 30884
rect 11396 30828 15708 30884
rect 15764 30828 15774 30884
rect 20290 30828 20300 30884
rect 20356 30828 21196 30884
rect 21252 30828 29708 30884
rect 29764 30828 29774 30884
rect 41682 30828 41692 30884
rect 41748 30828 50428 30884
rect 22054 30716 22092 30772
rect 22148 30716 22158 30772
rect 50194 30716 50204 30772
rect 50260 30716 50876 30772
rect 50932 30716 50942 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 22194 30380 22204 30436
rect 22260 30380 23100 30436
rect 23156 30380 23166 30436
rect 51538 30380 51548 30436
rect 51604 30380 55132 30436
rect 55188 30380 55198 30436
rect 29586 30268 29596 30324
rect 29652 30268 30044 30324
rect 30100 30268 30110 30324
rect 46946 30268 46956 30324
rect 47012 30268 49980 30324
rect 50036 30268 50046 30324
rect 51762 30268 51772 30324
rect 51828 30268 52668 30324
rect 52724 30268 52734 30324
rect 8418 30156 8428 30212
rect 8484 30156 14252 30212
rect 14308 30156 14318 30212
rect 19618 30156 19628 30212
rect 19684 30156 20524 30212
rect 20580 30156 20590 30212
rect 23986 30156 23996 30212
rect 24052 30156 25900 30212
rect 25956 30156 28140 30212
rect 28196 30156 28206 30212
rect 31266 30156 31276 30212
rect 31332 30156 33740 30212
rect 33796 30156 35084 30212
rect 35140 30156 35150 30212
rect 37090 30156 37100 30212
rect 37156 30156 38668 30212
rect 42354 30156 42364 30212
rect 42420 30156 45276 30212
rect 45332 30156 45612 30212
rect 45668 30156 45678 30212
rect 48738 30156 48748 30212
rect 48804 30156 49868 30212
rect 49924 30156 50876 30212
rect 50932 30156 50942 30212
rect 8372 30044 10108 30100
rect 10164 30044 10556 30100
rect 10612 30044 10622 30100
rect 16482 30044 16492 30100
rect 16548 30044 17052 30100
rect 17108 30044 17118 30100
rect 20962 30044 20972 30100
rect 21028 30044 21532 30100
rect 21588 30044 21598 30100
rect 21858 30044 21868 30100
rect 21924 30044 22316 30100
rect 22372 30044 24220 30100
rect 24276 30044 24286 30100
rect 30482 30044 30492 30100
rect 30548 30044 31164 30100
rect 31220 30044 31230 30100
rect 8372 29988 8428 30044
rect 7746 29932 7756 29988
rect 7812 29932 8428 29988
rect 8866 29932 8876 29988
rect 8932 29932 9660 29988
rect 9716 29932 9726 29988
rect 15810 29932 15820 29988
rect 15876 29932 16604 29988
rect 16660 29932 17836 29988
rect 17892 29932 20356 29988
rect 22194 29932 22204 29988
rect 22260 29932 22876 29988
rect 22932 29932 22942 29988
rect 24434 29932 24444 29988
rect 24500 29932 25452 29988
rect 25508 29932 25518 29988
rect 38612 29932 38668 30156
rect 38724 29932 40348 29988
rect 40404 29932 41916 29988
rect 41972 29932 41982 29988
rect 53218 29932 53228 29988
rect 53284 29932 54572 29988
rect 54628 29932 54638 29988
rect 54898 29932 54908 29988
rect 54964 29932 57036 29988
rect 57092 29932 57484 29988
rect 57540 29932 57550 29988
rect 20300 29876 20356 29932
rect 24444 29876 24500 29932
rect 9314 29820 9324 29876
rect 9380 29820 10892 29876
rect 10948 29820 11564 29876
rect 11620 29820 11630 29876
rect 20300 29820 24500 29876
rect 37762 29820 37772 29876
rect 37828 29820 39788 29876
rect 39844 29820 39854 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 8082 29708 8092 29764
rect 8148 29708 10780 29764
rect 10836 29708 10846 29764
rect 11330 29596 11340 29652
rect 11396 29596 12348 29652
rect 12404 29596 12414 29652
rect 23202 29596 23212 29652
rect 23268 29596 25564 29652
rect 25620 29596 25630 29652
rect 26898 29596 26908 29652
rect 26964 29596 27804 29652
rect 27860 29596 27870 29652
rect 28018 29596 28028 29652
rect 28084 29596 29036 29652
rect 29092 29596 29932 29652
rect 29988 29596 30604 29652
rect 30660 29596 30670 29652
rect 31602 29596 31612 29652
rect 31668 29596 34748 29652
rect 34804 29596 34814 29652
rect 49074 29596 49084 29652
rect 49140 29596 51100 29652
rect 51156 29596 51166 29652
rect 56914 29596 56924 29652
rect 56980 29596 57372 29652
rect 57428 29596 58156 29652
rect 58212 29596 58222 29652
rect 9090 29484 9100 29540
rect 9156 29484 9772 29540
rect 9828 29484 11116 29540
rect 11172 29484 11182 29540
rect 11442 29484 11452 29540
rect 11508 29484 13468 29540
rect 13524 29484 13534 29540
rect 21522 29484 21532 29540
rect 21588 29484 22092 29540
rect 22148 29484 22158 29540
rect 22418 29484 22428 29540
rect 22484 29484 23660 29540
rect 23716 29484 23726 29540
rect 27682 29484 27692 29540
rect 27748 29484 28476 29540
rect 28532 29484 28542 29540
rect 29474 29484 29484 29540
rect 29540 29484 31276 29540
rect 31332 29484 31342 29540
rect 51538 29484 51548 29540
rect 51604 29484 53004 29540
rect 53060 29484 53070 29540
rect 11452 29428 11508 29484
rect 29484 29428 29540 29484
rect 7186 29372 7196 29428
rect 7252 29372 9548 29428
rect 9604 29372 9614 29428
rect 10770 29372 10780 29428
rect 10836 29372 11508 29428
rect 13122 29372 13132 29428
rect 13188 29372 15148 29428
rect 15204 29372 15214 29428
rect 15474 29372 15484 29428
rect 15540 29372 16884 29428
rect 24770 29372 24780 29428
rect 24836 29372 25228 29428
rect 25284 29372 27580 29428
rect 27636 29372 29540 29428
rect 36866 29372 36876 29428
rect 36932 29372 37884 29428
rect 37940 29372 37950 29428
rect 50978 29372 50988 29428
rect 51044 29372 53228 29428
rect 53284 29372 53294 29428
rect 16828 29316 16884 29372
rect 12114 29260 12124 29316
rect 12180 29260 12796 29316
rect 12852 29260 15596 29316
rect 15652 29260 15662 29316
rect 16818 29260 16828 29316
rect 16884 29260 17388 29316
rect 17444 29260 17454 29316
rect 26450 29260 26460 29316
rect 26516 29260 27692 29316
rect 27748 29260 27758 29316
rect 28130 29260 28140 29316
rect 28196 29260 29708 29316
rect 29764 29260 29774 29316
rect 30930 29260 30940 29316
rect 30996 29260 31948 29316
rect 32004 29260 36540 29316
rect 36596 29260 36606 29316
rect 40226 29260 40236 29316
rect 40292 29260 41468 29316
rect 41524 29260 46508 29316
rect 46564 29260 46574 29316
rect 13430 29148 13468 29204
rect 13524 29148 13534 29204
rect 15362 29148 15372 29204
rect 15428 29148 21084 29204
rect 21140 29148 22876 29204
rect 22932 29148 22942 29204
rect 25554 29148 25564 29204
rect 25620 29148 35084 29204
rect 35140 29148 35150 29204
rect 39106 29148 39116 29204
rect 39172 29148 40124 29204
rect 40180 29148 40190 29204
rect 41794 29148 41804 29204
rect 41860 29148 42812 29204
rect 42868 29148 42878 29204
rect 12338 29036 12348 29092
rect 12404 29036 13580 29092
rect 13636 29036 13646 29092
rect 14802 29036 14812 29092
rect 14868 29036 15148 29092
rect 16370 29036 16380 29092
rect 16436 29036 18844 29092
rect 18900 29036 18910 29092
rect 20748 29036 26348 29092
rect 26404 29036 26414 29092
rect 30706 29036 30716 29092
rect 30772 29036 31388 29092
rect 31444 29036 31454 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 15092 28980 15148 29036
rect 20748 28980 20804 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 5058 28924 5068 28980
rect 5124 28924 8428 28980
rect 15092 28924 20804 28980
rect 21634 28924 21644 28980
rect 21700 28924 26908 28980
rect 26964 28924 26974 28980
rect 28140 28924 34580 28980
rect 8372 28756 8428 28924
rect 28140 28868 28196 28924
rect 34524 28868 34580 28924
rect 38612 28924 47964 28980
rect 48020 28924 48030 28980
rect 38612 28868 38668 28924
rect 14018 28812 14028 28868
rect 14084 28812 16380 28868
rect 16436 28812 16446 28868
rect 17602 28812 17612 28868
rect 17668 28812 18172 28868
rect 18228 28812 18238 28868
rect 19618 28812 19628 28868
rect 19684 28812 28196 28868
rect 28354 28812 28364 28868
rect 28420 28812 30604 28868
rect 30660 28812 30670 28868
rect 34524 28812 35308 28868
rect 35364 28812 35980 28868
rect 36036 28812 38668 28868
rect 49634 28812 49644 28868
rect 49700 28812 50652 28868
rect 50708 28812 50718 28868
rect 8372 28700 14924 28756
rect 14980 28700 14990 28756
rect 15092 28700 15820 28756
rect 15876 28700 15886 28756
rect 26852 28700 30380 28756
rect 30436 28700 30446 28756
rect 44370 28700 44380 28756
rect 44436 28700 45276 28756
rect 45332 28700 45342 28756
rect 48514 28700 48524 28756
rect 48580 28700 49756 28756
rect 49812 28700 49822 28756
rect 51426 28700 51436 28756
rect 51492 28700 55356 28756
rect 55412 28700 56588 28756
rect 56644 28700 58044 28756
rect 58100 28700 58110 28756
rect 15092 28644 15148 28700
rect 26852 28644 26908 28700
rect 4274 28588 4284 28644
rect 4340 28588 4732 28644
rect 4788 28588 6972 28644
rect 7028 28588 9660 28644
rect 9716 28588 9726 28644
rect 13692 28588 14028 28644
rect 14084 28588 14094 28644
rect 14802 28588 14812 28644
rect 14868 28588 15148 28644
rect 18162 28588 18172 28644
rect 18228 28588 18956 28644
rect 19012 28588 19022 28644
rect 25442 28588 25452 28644
rect 25508 28588 26908 28644
rect 29698 28588 29708 28644
rect 29764 28588 30268 28644
rect 30324 28588 31164 28644
rect 31220 28588 31230 28644
rect 35074 28588 35084 28644
rect 35140 28588 36092 28644
rect 36148 28588 37324 28644
rect 37380 28588 37390 28644
rect 45388 28588 53900 28644
rect 53956 28588 54236 28644
rect 54292 28588 54302 28644
rect 13692 28532 13748 28588
rect 45388 28532 45444 28588
rect 13682 28476 13692 28532
rect 13748 28476 13758 28532
rect 17490 28476 17500 28532
rect 17556 28476 18620 28532
rect 18676 28476 18686 28532
rect 40898 28476 40908 28532
rect 40964 28476 45444 28532
rect 52994 28476 53004 28532
rect 53060 28476 53564 28532
rect 53620 28476 53630 28532
rect 55122 28476 55132 28532
rect 55188 28476 56588 28532
rect 56644 28476 56654 28532
rect 14018 28364 14028 28420
rect 14084 28364 15708 28420
rect 15764 28364 15774 28420
rect 17042 28364 17052 28420
rect 17108 28364 18284 28420
rect 18340 28364 18350 28420
rect 37314 28364 37324 28420
rect 37380 28364 38108 28420
rect 38164 28364 38174 28420
rect 43362 28364 43372 28420
rect 43428 28364 44044 28420
rect 44100 28364 44110 28420
rect 50082 28364 50092 28420
rect 50148 28364 51660 28420
rect 51716 28364 51726 28420
rect 13906 28252 13916 28308
rect 13972 28252 13982 28308
rect 13916 28196 13972 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 9538 28140 9548 28196
rect 9604 28140 11004 28196
rect 11060 28140 11070 28196
rect 13916 28140 14364 28196
rect 14420 28140 14430 28196
rect 37426 28140 37436 28196
rect 37492 28140 38108 28196
rect 38164 28140 38174 28196
rect 55458 28140 55468 28196
rect 55524 28140 55534 28196
rect 55468 28084 55524 28140
rect 17154 28028 17164 28084
rect 17220 28028 18172 28084
rect 18228 28028 18238 28084
rect 26852 28028 28252 28084
rect 28308 28028 34972 28084
rect 35028 28028 38780 28084
rect 38836 28028 38846 28084
rect 39228 28028 55524 28084
rect 10994 27916 11004 27972
rect 11060 27916 15260 27972
rect 15316 27916 15326 27972
rect 7970 27804 7980 27860
rect 8036 27804 9548 27860
rect 9604 27804 9614 27860
rect 9874 27804 9884 27860
rect 9940 27804 14700 27860
rect 14756 27804 14766 27860
rect 19618 27804 19628 27860
rect 19684 27804 22876 27860
rect 22932 27804 22942 27860
rect 26852 27748 26908 28028
rect 30370 27916 30380 27972
rect 30436 27916 31052 27972
rect 31108 27916 32060 27972
rect 32116 27916 32126 27972
rect 38434 27916 38444 27972
rect 38500 27916 39004 27972
rect 39060 27916 39070 27972
rect 39228 27860 39284 28028
rect 52770 27916 52780 27972
rect 52836 27916 55188 27972
rect 55458 27916 55468 27972
rect 55524 27916 57260 27972
rect 57316 27916 57326 27972
rect 57922 27916 57932 27972
rect 57988 27916 58156 27972
rect 58212 27916 58222 27972
rect 55132 27860 55188 27916
rect 31490 27804 31500 27860
rect 31556 27804 32508 27860
rect 32564 27804 33404 27860
rect 33460 27804 34524 27860
rect 34580 27804 34590 27860
rect 34748 27804 39284 27860
rect 41122 27804 41132 27860
rect 41188 27804 41916 27860
rect 41972 27804 41982 27860
rect 50306 27804 50316 27860
rect 50372 27804 51436 27860
rect 51492 27804 51502 27860
rect 53330 27804 53340 27860
rect 53396 27804 53676 27860
rect 53732 27804 53742 27860
rect 55122 27804 55132 27860
rect 55188 27804 55198 27860
rect 34748 27748 34804 27804
rect 56812 27748 56868 27916
rect 5394 27692 5404 27748
rect 5460 27692 13356 27748
rect 13412 27692 13422 27748
rect 15698 27692 15708 27748
rect 15764 27692 25788 27748
rect 25844 27692 26908 27748
rect 30146 27692 30156 27748
rect 30212 27692 34804 27748
rect 38098 27692 38108 27748
rect 38164 27692 38668 27748
rect 38724 27692 38734 27748
rect 53442 27692 53452 27748
rect 53508 27692 54236 27748
rect 54292 27692 54302 27748
rect 56802 27692 56812 27748
rect 56868 27692 56878 27748
rect 8642 27580 8652 27636
rect 8708 27580 10108 27636
rect 10164 27580 10174 27636
rect 15810 27580 15820 27636
rect 15876 27580 17612 27636
rect 17668 27580 17678 27636
rect 18610 27580 18620 27636
rect 18676 27580 19292 27636
rect 19348 27580 34860 27636
rect 34916 27580 37772 27636
rect 37828 27580 39116 27636
rect 39172 27580 39182 27636
rect 56914 27580 56924 27636
rect 56980 27580 57932 27636
rect 57988 27580 57998 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 7298 27356 7308 27412
rect 7364 27356 11004 27412
rect 11060 27356 11070 27412
rect 7858 27244 7868 27300
rect 7924 27244 11564 27300
rect 11620 27244 12348 27300
rect 12404 27244 13132 27300
rect 13188 27244 13198 27300
rect 37090 27244 37100 27300
rect 37156 27244 38220 27300
rect 38276 27244 38668 27300
rect 38724 27244 55020 27300
rect 55076 27244 55086 27300
rect 12002 27132 12012 27188
rect 12068 27132 13916 27188
rect 13972 27132 13982 27188
rect 14476 27132 15148 27188
rect 15204 27132 15214 27188
rect 38882 27132 38892 27188
rect 38948 27132 40012 27188
rect 40068 27132 40908 27188
rect 40964 27132 40974 27188
rect 41906 27132 41916 27188
rect 41972 27132 42588 27188
rect 42644 27132 42654 27188
rect 56690 27132 56700 27188
rect 56756 27132 58156 27188
rect 58212 27132 58222 27188
rect 14476 27076 14532 27132
rect 5618 27020 5628 27076
rect 5684 27020 6748 27076
rect 6804 27020 7420 27076
rect 7476 27020 7486 27076
rect 12338 27020 12348 27076
rect 12404 27020 13580 27076
rect 13636 27020 14532 27076
rect 14690 27020 14700 27076
rect 14756 27020 15932 27076
rect 15988 27020 15998 27076
rect 26338 27020 26348 27076
rect 26404 27020 26414 27076
rect 26786 27020 26796 27076
rect 26852 27020 28028 27076
rect 28084 27020 28700 27076
rect 28756 27020 28766 27076
rect 26348 26964 26404 27020
rect 12226 26908 12236 26964
rect 12292 26908 14364 26964
rect 14420 26908 15260 26964
rect 15316 26908 15326 26964
rect 15698 26908 15708 26964
rect 15764 26908 15774 26964
rect 22866 26908 22876 26964
rect 22932 26908 23996 26964
rect 24052 26908 26404 26964
rect 36978 26908 36988 26964
rect 37044 26908 38108 26964
rect 38164 26908 38174 26964
rect 44258 26908 44268 26964
rect 44324 26908 45164 26964
rect 45220 26908 45230 26964
rect 52098 26908 52108 26964
rect 52164 26908 52780 26964
rect 52836 26908 52846 26964
rect 53676 26908 54236 26964
rect 54292 26908 54302 26964
rect 15708 26852 15764 26908
rect 53676 26852 53732 26908
rect 7074 26796 7084 26852
rect 7140 26796 7868 26852
rect 7924 26796 10668 26852
rect 10724 26796 10734 26852
rect 11218 26796 11228 26852
rect 11284 26796 11788 26852
rect 11844 26796 11854 26852
rect 13234 26796 13244 26852
rect 13300 26796 15764 26852
rect 24546 26796 24556 26852
rect 24612 26796 24780 26852
rect 24836 26796 25340 26852
rect 25396 26796 26572 26852
rect 26628 26796 26638 26852
rect 43922 26796 43932 26852
rect 43988 26796 44828 26852
rect 44884 26796 44894 26852
rect 53666 26796 53676 26852
rect 53732 26796 53742 26852
rect 25442 26684 25452 26740
rect 25508 26684 25564 26740
rect 25620 26684 25630 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 22866 26572 22876 26628
rect 22932 26572 35420 26628
rect 35476 26572 37660 26628
rect 37716 26572 37726 26628
rect 14578 26460 14588 26516
rect 14644 26460 14924 26516
rect 14980 26460 15596 26516
rect 15652 26460 15662 26516
rect 15922 26460 15932 26516
rect 15988 26460 25116 26516
rect 25172 26460 25182 26516
rect 25890 26460 25900 26516
rect 25956 26460 27020 26516
rect 27076 26460 27356 26516
rect 27412 26460 27422 26516
rect 27794 26460 27804 26516
rect 27860 26460 28476 26516
rect 28532 26460 29596 26516
rect 29652 26460 29662 26516
rect 34402 26460 34412 26516
rect 34468 26460 37100 26516
rect 37156 26460 37166 26516
rect 37986 26460 37996 26516
rect 38052 26460 38444 26516
rect 38500 26460 39228 26516
rect 39284 26460 39294 26516
rect 39442 26460 39452 26516
rect 39508 26460 40124 26516
rect 40180 26460 41916 26516
rect 41972 26460 41982 26516
rect 43698 26460 43708 26516
rect 43764 26460 47852 26516
rect 47908 26460 47918 26516
rect 56018 26460 56028 26516
rect 56084 26460 57036 26516
rect 57092 26460 57102 26516
rect 16594 26348 16604 26404
rect 16660 26348 17052 26404
rect 17108 26348 17118 26404
rect 17378 26348 17388 26404
rect 17444 26348 18060 26404
rect 18116 26348 18126 26404
rect 26226 26348 26236 26404
rect 26292 26348 27468 26404
rect 27524 26348 28812 26404
rect 28868 26348 28878 26404
rect 41458 26348 41468 26404
rect 41524 26348 46396 26404
rect 46452 26348 46462 26404
rect 2258 26236 2268 26292
rect 2324 26236 12516 26292
rect 16818 26236 16828 26292
rect 16884 26236 17724 26292
rect 17780 26236 17790 26292
rect 25554 26236 25564 26292
rect 25620 26236 26124 26292
rect 26180 26236 26190 26292
rect 26562 26236 26572 26292
rect 26628 26236 28252 26292
rect 28308 26236 28318 26292
rect 28578 26236 28588 26292
rect 28644 26236 29148 26292
rect 29204 26236 29372 26292
rect 29428 26236 29438 26292
rect 39442 26236 39452 26292
rect 39508 26236 40684 26292
rect 40740 26236 41132 26292
rect 41188 26236 41198 26292
rect 12460 26180 12516 26236
rect 8194 26124 8204 26180
rect 8260 26124 10556 26180
rect 10612 26124 10622 26180
rect 12460 26124 22316 26180
rect 22372 26124 22764 26180
rect 22820 26124 23324 26180
rect 23380 26124 23772 26180
rect 23828 26124 23838 26180
rect 24098 26124 24108 26180
rect 24164 26124 26908 26180
rect 26964 26124 26974 26180
rect 33282 26124 33292 26180
rect 33348 26124 39676 26180
rect 39732 26124 39742 26180
rect 24556 26012 26124 26068
rect 26180 26012 26190 26068
rect 26338 26012 26348 26068
rect 26404 26012 26908 26068
rect 30258 26012 30268 26068
rect 30324 26012 39116 26068
rect 39172 26012 39788 26068
rect 39844 26012 41020 26068
rect 41076 26012 41086 26068
rect 47618 26012 47628 26068
rect 47684 26012 49084 26068
rect 49140 26012 49150 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 24556 25844 24612 26012
rect 26852 25956 26908 26012
rect 26002 25900 26012 25956
rect 26068 25900 26572 25956
rect 26628 25900 26638 25956
rect 26852 25900 32396 25956
rect 32452 25900 32462 25956
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 23202 25788 23212 25844
rect 23268 25788 24556 25844
rect 24612 25788 24622 25844
rect 25900 25788 26684 25844
rect 26740 25788 26750 25844
rect 25900 25732 25956 25788
rect 17714 25676 17724 25732
rect 17780 25676 24108 25732
rect 24164 25676 24174 25732
rect 25554 25676 25564 25732
rect 25620 25676 25900 25732
rect 25956 25676 25966 25732
rect 26348 25676 27804 25732
rect 27860 25676 33180 25732
rect 33236 25676 33246 25732
rect 37314 25676 37324 25732
rect 37380 25676 40348 25732
rect 40404 25676 40414 25732
rect 43922 25676 43932 25732
rect 43988 25676 44940 25732
rect 44996 25676 45006 25732
rect 26348 25620 26404 25676
rect 19170 25564 19180 25620
rect 19236 25564 19964 25620
rect 20020 25564 20030 25620
rect 24658 25564 24668 25620
rect 24724 25564 26124 25620
rect 26180 25564 26190 25620
rect 26338 25564 26348 25620
rect 26404 25564 26414 25620
rect 26898 25564 26908 25620
rect 26964 25564 27692 25620
rect 27748 25564 27758 25620
rect 27906 25564 27916 25620
rect 27972 25564 28588 25620
rect 28644 25564 28654 25620
rect 34178 25564 34188 25620
rect 34244 25564 34972 25620
rect 35028 25564 36204 25620
rect 36260 25564 58268 25620
rect 58324 25564 58334 25620
rect 7634 25452 7644 25508
rect 7700 25452 8428 25508
rect 16594 25452 16604 25508
rect 16660 25452 17388 25508
rect 17444 25452 17454 25508
rect 24210 25452 24220 25508
rect 24276 25452 27244 25508
rect 27300 25452 27310 25508
rect 32610 25452 32620 25508
rect 32676 25452 33740 25508
rect 33796 25452 34636 25508
rect 34692 25452 40124 25508
rect 40180 25452 40684 25508
rect 40740 25452 40750 25508
rect 45042 25452 45052 25508
rect 45108 25452 45948 25508
rect 46004 25452 46014 25508
rect 46610 25452 46620 25508
rect 46676 25452 47292 25508
rect 47348 25452 47358 25508
rect 8372 25228 8428 25452
rect 45948 25396 46004 25452
rect 9314 25340 9324 25396
rect 9380 25340 13916 25396
rect 13972 25340 13982 25396
rect 16380 25340 16828 25396
rect 16884 25340 16894 25396
rect 24098 25340 24108 25396
rect 24164 25340 24668 25396
rect 24724 25340 24734 25396
rect 25890 25340 25900 25396
rect 25956 25340 27132 25396
rect 27188 25340 27198 25396
rect 35298 25340 35308 25396
rect 35364 25340 36764 25396
rect 36820 25340 37324 25396
rect 37380 25340 37390 25396
rect 37538 25340 37548 25396
rect 37604 25340 38332 25396
rect 38388 25340 38398 25396
rect 39218 25340 39228 25396
rect 39284 25340 40572 25396
rect 40628 25340 40638 25396
rect 41346 25340 41356 25396
rect 41412 25340 42476 25396
rect 42532 25340 43708 25396
rect 43764 25340 43774 25396
rect 45948 25340 46956 25396
rect 47012 25340 47022 25396
rect 52322 25340 52332 25396
rect 52388 25340 53676 25396
rect 53732 25340 53742 25396
rect 8484 25228 10444 25284
rect 10500 25228 12796 25284
rect 12852 25228 12862 25284
rect 16380 25172 16436 25340
rect 21746 25228 21756 25284
rect 21812 25228 22540 25284
rect 22596 25228 22606 25284
rect 24434 25228 24444 25284
rect 24500 25228 28028 25284
rect 28084 25228 29708 25284
rect 29764 25228 29774 25284
rect 33170 25228 33180 25284
rect 33236 25228 33740 25284
rect 33796 25228 34076 25284
rect 34132 25228 34142 25284
rect 36082 25228 36092 25284
rect 36148 25228 37100 25284
rect 37156 25228 37166 25284
rect 37426 25228 37436 25284
rect 37492 25228 37996 25284
rect 38052 25228 38062 25284
rect 41458 25228 41468 25284
rect 41524 25228 41916 25284
rect 41972 25228 44828 25284
rect 44884 25228 45836 25284
rect 45892 25228 45902 25284
rect 50194 25228 50204 25284
rect 50260 25228 52780 25284
rect 52836 25228 52846 25284
rect 57586 25228 57596 25284
rect 57652 25228 58156 25284
rect 58212 25228 58222 25284
rect 8866 25116 8876 25172
rect 8932 25116 9660 25172
rect 9716 25116 10220 25172
rect 10276 25116 13580 25172
rect 13636 25116 15036 25172
rect 15092 25116 15820 25172
rect 15876 25116 16436 25172
rect 21410 25116 21420 25172
rect 21476 25116 22204 25172
rect 22260 25116 22270 25172
rect 36530 25116 36540 25172
rect 36596 25116 39564 25172
rect 39620 25116 39630 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 14466 25004 14476 25060
rect 14532 25004 15148 25060
rect 15204 25004 18284 25060
rect 18340 25004 18350 25060
rect 29474 25004 29484 25060
rect 29540 25004 29932 25060
rect 29988 25004 33516 25060
rect 33572 25004 42140 25060
rect 42196 25004 43036 25060
rect 43092 25004 43102 25060
rect 16146 24892 16156 24948
rect 16212 24892 18172 24948
rect 18228 24892 19180 24948
rect 19236 24892 19246 24948
rect 25526 24892 25564 24948
rect 25620 24892 25630 24948
rect 27346 24892 27356 24948
rect 27412 24892 27692 24948
rect 27748 24892 29036 24948
rect 29092 24892 29102 24948
rect 12450 24780 12460 24836
rect 12516 24780 14252 24836
rect 14308 24780 14318 24836
rect 29138 24780 29148 24836
rect 29204 24780 29820 24836
rect 29876 24780 34188 24836
rect 34244 24780 41132 24836
rect 41188 24780 41198 24836
rect 13794 24668 13804 24724
rect 13860 24668 16492 24724
rect 16548 24668 16558 24724
rect 35410 24668 35420 24724
rect 35476 24668 38444 24724
rect 38500 24668 38510 24724
rect 38612 24668 41804 24724
rect 41860 24668 42700 24724
rect 42756 24668 43372 24724
rect 43428 24668 43438 24724
rect 52210 24668 52220 24724
rect 52276 24668 52892 24724
rect 52948 24668 54124 24724
rect 54180 24668 54190 24724
rect 56578 24668 56588 24724
rect 56644 24668 57148 24724
rect 57204 24668 57214 24724
rect 38612 24612 38668 24668
rect 10882 24556 10892 24612
rect 10948 24556 14364 24612
rect 14420 24556 14430 24612
rect 14578 24556 14588 24612
rect 14644 24556 15596 24612
rect 15652 24556 16380 24612
rect 16436 24556 16446 24612
rect 22642 24556 22652 24612
rect 22708 24556 23436 24612
rect 23492 24556 25228 24612
rect 25284 24556 25788 24612
rect 25844 24556 25854 24612
rect 31266 24556 31276 24612
rect 31332 24556 31836 24612
rect 31892 24556 35308 24612
rect 35364 24556 35374 24612
rect 35970 24556 35980 24612
rect 36036 24556 38668 24612
rect 43474 24556 43484 24612
rect 43540 24556 44828 24612
rect 44884 24556 48300 24612
rect 48356 24556 48366 24612
rect 48738 24556 48748 24612
rect 48804 24556 57484 24612
rect 57540 24556 57550 24612
rect 59200 24500 60000 24528
rect 26338 24444 26348 24500
rect 26404 24444 27020 24500
rect 27076 24444 27086 24500
rect 43586 24444 43596 24500
rect 43652 24444 45276 24500
rect 45332 24444 45342 24500
rect 58146 24444 58156 24500
rect 58212 24444 60000 24500
rect 59200 24416 60000 24444
rect 17602 24332 17612 24388
rect 17668 24332 18620 24388
rect 18676 24332 22988 24388
rect 23044 24332 28924 24388
rect 28980 24332 28990 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 18834 23996 18844 24052
rect 18900 23996 19404 24052
rect 19460 23996 20412 24052
rect 20468 23996 20478 24052
rect 40226 23996 40236 24052
rect 40292 23996 44604 24052
rect 44660 23996 45500 24052
rect 45556 23996 45566 24052
rect 52770 23996 52780 24052
rect 52836 23996 53452 24052
rect 53508 23996 53518 24052
rect 16370 23884 16380 23940
rect 16436 23884 18956 23940
rect 19012 23884 19022 23940
rect 22194 23884 22204 23940
rect 22260 23884 28252 23940
rect 28308 23884 28318 23940
rect 53218 23884 53228 23940
rect 53284 23884 54460 23940
rect 54516 23884 54526 23940
rect 24322 23772 24332 23828
rect 24388 23772 25340 23828
rect 25396 23772 25900 23828
rect 25956 23772 25966 23828
rect 43250 23772 43260 23828
rect 43316 23772 43708 23828
rect 43764 23772 44044 23828
rect 44100 23772 44110 23828
rect 52882 23772 52892 23828
rect 52948 23772 53452 23828
rect 53508 23772 53518 23828
rect 15810 23660 15820 23716
rect 15876 23660 16604 23716
rect 16660 23660 16670 23716
rect 18274 23660 18284 23716
rect 18340 23660 19852 23716
rect 19908 23660 20748 23716
rect 20804 23660 20814 23716
rect 40002 23660 40012 23716
rect 40068 23660 43596 23716
rect 43652 23660 43662 23716
rect 51426 23660 51436 23716
rect 51492 23660 53004 23716
rect 53060 23660 53070 23716
rect 22418 23548 22428 23604
rect 22484 23548 23100 23604
rect 23156 23548 24892 23604
rect 24948 23548 26908 23604
rect 26964 23548 26974 23604
rect 41916 23548 42924 23604
rect 42980 23548 44940 23604
rect 44996 23548 45388 23604
rect 45444 23548 45454 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41916 23492 41972 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 20188 23436 38668 23492
rect 41234 23436 41244 23492
rect 41300 23436 41972 23492
rect 45826 23436 45836 23492
rect 45892 23436 46844 23492
rect 46900 23436 46910 23492
rect 20188 23380 20244 23436
rect 38612 23380 38668 23436
rect 18946 23324 18956 23380
rect 19012 23324 19628 23380
rect 19684 23324 20244 23380
rect 21970 23324 21980 23380
rect 22036 23324 22876 23380
rect 22932 23324 23436 23380
rect 23492 23324 23502 23380
rect 23986 23324 23996 23380
rect 24052 23324 27580 23380
rect 27636 23324 30716 23380
rect 30772 23324 33180 23380
rect 33236 23324 33246 23380
rect 38612 23324 44156 23380
rect 44212 23324 45052 23380
rect 45108 23324 48748 23380
rect 48804 23324 48814 23380
rect 55122 23324 55132 23380
rect 55188 23324 56700 23380
rect 56756 23324 56766 23380
rect 20738 23212 20748 23268
rect 20804 23212 25508 23268
rect 26786 23212 26796 23268
rect 26852 23212 27356 23268
rect 27412 23212 27422 23268
rect 28802 23212 28812 23268
rect 28868 23212 38108 23268
rect 38164 23212 39228 23268
rect 39284 23212 39294 23268
rect 44930 23212 44940 23268
rect 44996 23212 45612 23268
rect 45668 23212 45678 23268
rect 52210 23212 52220 23268
rect 52276 23212 54124 23268
rect 54180 23212 54190 23268
rect 56578 23212 56588 23268
rect 56644 23212 57932 23268
rect 57988 23212 57998 23268
rect 25452 23156 25508 23212
rect 22978 23100 22988 23156
rect 23044 23100 24220 23156
rect 24276 23100 24286 23156
rect 24434 23100 24444 23156
rect 24500 23100 25228 23156
rect 25284 23100 25294 23156
rect 25452 23100 33628 23156
rect 33684 23100 34076 23156
rect 34132 23100 34142 23156
rect 37874 23100 37884 23156
rect 37940 23100 38444 23156
rect 38500 23100 41020 23156
rect 41076 23100 41086 23156
rect 42242 23100 42252 23156
rect 42308 23100 44156 23156
rect 44212 23100 44222 23156
rect 47954 23100 47964 23156
rect 48020 23100 50428 23156
rect 50484 23100 50494 23156
rect 50372 23044 50428 23100
rect 16706 22988 16716 23044
rect 16772 22988 17500 23044
rect 17556 22988 17566 23044
rect 46498 22988 46508 23044
rect 46564 22988 48188 23044
rect 48244 22988 48254 23044
rect 50372 22988 50764 23044
rect 50820 22988 51212 23044
rect 51268 22988 53340 23044
rect 53396 22988 54684 23044
rect 54740 22988 54750 23044
rect 22642 22764 22652 22820
rect 22708 22764 31948 22820
rect 32004 22764 33516 22820
rect 33572 22764 33582 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 35522 22540 35532 22596
rect 35588 22540 36428 22596
rect 36484 22540 38556 22596
rect 38612 22540 38622 22596
rect 33170 22428 33180 22484
rect 33236 22428 33516 22484
rect 33572 22428 33582 22484
rect 38770 22428 38780 22484
rect 38836 22428 40684 22484
rect 40740 22428 45724 22484
rect 45780 22428 45790 22484
rect 48178 22428 48188 22484
rect 48244 22428 50204 22484
rect 50260 22428 50270 22484
rect 45602 22316 45612 22372
rect 45668 22316 46732 22372
rect 46788 22316 46798 22372
rect 56802 22316 56812 22372
rect 56868 22316 57372 22372
rect 57428 22316 57438 22372
rect 23874 22204 23884 22260
rect 23940 22204 24108 22260
rect 24164 22204 25228 22260
rect 25284 22204 27804 22260
rect 27860 22204 27870 22260
rect 37314 22204 37324 22260
rect 37380 22204 38444 22260
rect 38500 22204 38510 22260
rect 41458 22204 41468 22260
rect 41524 22204 42028 22260
rect 42084 22204 42094 22260
rect 43698 22204 43708 22260
rect 43764 22204 45388 22260
rect 45444 22204 45948 22260
rect 46004 22204 46014 22260
rect 54562 22204 54572 22260
rect 54628 22204 57036 22260
rect 57092 22204 57102 22260
rect 33394 22092 33404 22148
rect 33460 22092 46396 22148
rect 46452 22092 47180 22148
rect 47236 22092 47246 22148
rect 56914 22092 56924 22148
rect 56980 22092 57596 22148
rect 57652 22092 57662 22148
rect 55122 21980 55132 22036
rect 55188 21980 57148 22036
rect 57204 21980 57214 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 44146 21868 44156 21924
rect 44212 21868 49084 21924
rect 49140 21868 49150 21924
rect 18610 21756 18620 21812
rect 18676 21756 19292 21812
rect 19348 21756 19964 21812
rect 20020 21756 25340 21812
rect 25396 21756 25406 21812
rect 28466 21756 28476 21812
rect 28532 21756 33628 21812
rect 33684 21756 36316 21812
rect 36372 21756 36764 21812
rect 36820 21756 36830 21812
rect 40338 21756 40348 21812
rect 40404 21756 41580 21812
rect 41636 21756 41646 21812
rect 46946 21756 46956 21812
rect 47012 21756 49644 21812
rect 49700 21756 49710 21812
rect 18946 21644 18956 21700
rect 19012 21644 20076 21700
rect 20132 21644 20142 21700
rect 31938 21644 31948 21700
rect 32004 21644 34524 21700
rect 34580 21644 34590 21700
rect 49746 21644 49756 21700
rect 49812 21644 50988 21700
rect 51044 21644 51054 21700
rect 21746 21532 21756 21588
rect 21812 21532 23996 21588
rect 24052 21532 24892 21588
rect 24948 21532 24958 21588
rect 34850 21532 34860 21588
rect 34916 21532 35644 21588
rect 35700 21532 35710 21588
rect 54786 21532 54796 21588
rect 54852 21532 55132 21588
rect 55188 21532 55198 21588
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 18722 20860 18732 20916
rect 18788 20860 19404 20916
rect 19460 20860 20300 20916
rect 20356 20860 29372 20916
rect 29428 20860 30156 20916
rect 30212 20860 30222 20916
rect 20514 20748 20524 20804
rect 20580 20748 22652 20804
rect 22708 20748 22718 20804
rect 30706 20748 30716 20804
rect 30772 20748 33964 20804
rect 34020 20748 34030 20804
rect 15922 20636 15932 20692
rect 15988 20636 18508 20692
rect 18564 20636 18574 20692
rect 20738 20636 20748 20692
rect 20804 20636 21868 20692
rect 21924 20636 21934 20692
rect 18386 20524 18396 20580
rect 18452 20524 19628 20580
rect 19684 20524 21756 20580
rect 21812 20524 21822 20580
rect 27570 20524 27580 20580
rect 27636 20524 31276 20580
rect 31332 20524 31342 20580
rect 28914 20412 28924 20468
rect 28980 20412 33740 20468
rect 33796 20412 33806 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 14802 20188 14812 20244
rect 14868 20188 15260 20244
rect 15316 20188 16884 20244
rect 16828 20020 16884 20188
rect 31388 20188 31948 20244
rect 32004 20188 32014 20244
rect 37202 20188 37212 20244
rect 37268 20188 37772 20244
rect 37828 20188 38556 20244
rect 38612 20188 38622 20244
rect 18162 20076 18172 20132
rect 18228 20076 18620 20132
rect 18676 20076 18686 20132
rect 26786 20076 26796 20132
rect 26852 20076 27132 20132
rect 27188 20076 27198 20132
rect 27458 20076 27468 20132
rect 27524 20076 28476 20132
rect 28532 20076 28542 20132
rect 31388 20020 31444 20188
rect 31602 20076 31612 20132
rect 31668 20076 32060 20132
rect 32116 20076 32126 20132
rect 40338 20076 40348 20132
rect 40404 20076 41244 20132
rect 41300 20076 46340 20132
rect 46284 20020 46340 20076
rect 16828 19964 18060 20020
rect 18116 19964 19404 20020
rect 19460 19964 19470 20020
rect 26562 19964 26572 20020
rect 26628 19964 27356 20020
rect 27412 19964 27422 20020
rect 28242 19964 28252 20020
rect 28308 19964 30492 20020
rect 30548 19964 31052 20020
rect 31108 19964 31118 20020
rect 31378 19964 31388 20020
rect 31444 19964 31454 20020
rect 41458 19964 41468 20020
rect 41524 19964 42140 20020
rect 42196 19964 42206 20020
rect 44594 19964 44604 20020
rect 44660 19964 45276 20020
rect 45332 19964 45342 20020
rect 46274 19964 46284 20020
rect 46340 19964 46844 20020
rect 46900 19964 46910 20020
rect 47282 19964 47292 20020
rect 47348 19964 47964 20020
rect 48020 19964 48030 20020
rect 21970 19852 21980 19908
rect 22036 19852 22876 19908
rect 22932 19852 22942 19908
rect 27122 19852 27132 19908
rect 27188 19852 27692 19908
rect 27748 19852 29148 19908
rect 29204 19852 29214 19908
rect 41010 19852 41020 19908
rect 41076 19852 42588 19908
rect 42644 19852 42654 19908
rect 46722 19852 46732 19908
rect 46788 19852 47852 19908
rect 47908 19852 47918 19908
rect 46946 19740 46956 19796
rect 47012 19740 47516 19796
rect 47572 19740 47582 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 38658 19516 38668 19572
rect 38724 19516 38780 19572
rect 38836 19516 40908 19572
rect 40964 19516 40974 19572
rect 34290 19404 34300 19460
rect 34356 19404 36988 19460
rect 37044 19404 42252 19460
rect 42308 19404 42318 19460
rect 46162 19404 46172 19460
rect 46228 19404 47628 19460
rect 47684 19404 47694 19460
rect 19058 19292 19068 19348
rect 19124 19292 26236 19348
rect 26292 19292 26796 19348
rect 26852 19292 26862 19348
rect 34178 19292 34188 19348
rect 34244 19292 34636 19348
rect 34692 19292 39060 19348
rect 39330 19292 39340 19348
rect 39396 19292 39788 19348
rect 39844 19292 44604 19348
rect 44660 19292 44670 19348
rect 23202 19180 23212 19236
rect 23268 19180 23660 19236
rect 23716 19180 24332 19236
rect 24388 19180 25004 19236
rect 25060 19180 25070 19236
rect 34066 19180 34076 19236
rect 34132 19180 35420 19236
rect 35476 19180 35486 19236
rect 37090 19180 37100 19236
rect 37156 19180 38668 19236
rect 38724 19180 38734 19236
rect 39004 19124 39060 19292
rect 40338 19180 40348 19236
rect 40404 19180 40414 19236
rect 47170 19180 47180 19236
rect 47236 19180 50092 19236
rect 50148 19180 50158 19236
rect 40348 19124 40404 19180
rect 29932 19068 31500 19124
rect 31556 19068 31948 19124
rect 32004 19068 32014 19124
rect 39004 19068 40404 19124
rect 47730 19068 47740 19124
rect 47796 19068 50876 19124
rect 50932 19068 50942 19124
rect 29932 19012 29988 19068
rect 17154 18956 17164 19012
rect 17220 18956 17836 19012
rect 17892 18956 18508 19012
rect 18564 18956 18574 19012
rect 28466 18956 28476 19012
rect 28532 18956 29932 19012
rect 29988 18956 29998 19012
rect 30146 18956 30156 19012
rect 30212 18956 30716 19012
rect 30772 18956 31052 19012
rect 31108 18956 31118 19012
rect 34962 18956 34972 19012
rect 35028 18956 38332 19012
rect 38388 18956 38398 19012
rect 38546 18956 38556 19012
rect 38612 18956 38892 19012
rect 38948 18956 38958 19012
rect 42018 18956 42028 19012
rect 42084 18956 44716 19012
rect 44772 18956 44782 19012
rect 50754 18956 50764 19012
rect 50820 18956 50988 19012
rect 51044 18956 51054 19012
rect 51202 18956 51212 19012
rect 51268 18956 51436 19012
rect 51492 18956 51884 19012
rect 51940 18956 51950 19012
rect 38332 18900 38388 18956
rect 38332 18844 40236 18900
rect 40292 18844 40302 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 33058 18732 33068 18788
rect 33124 18732 35364 18788
rect 36306 18732 36316 18788
rect 36372 18732 37884 18788
rect 37940 18732 39564 18788
rect 39620 18732 41244 18788
rect 41300 18732 41310 18788
rect 35308 18676 35364 18732
rect 29362 18620 29372 18676
rect 29428 18620 30604 18676
rect 30660 18620 33852 18676
rect 33908 18620 35084 18676
rect 35140 18620 35150 18676
rect 35308 18620 42364 18676
rect 42420 18620 43148 18676
rect 43204 18620 45276 18676
rect 45332 18620 45948 18676
rect 46004 18620 46014 18676
rect 24210 18508 24220 18564
rect 24276 18508 33628 18564
rect 33684 18508 34636 18564
rect 34692 18508 34702 18564
rect 35970 18508 35980 18564
rect 36036 18508 37100 18564
rect 37156 18508 37166 18564
rect 40898 18508 40908 18564
rect 40964 18508 42140 18564
rect 42196 18508 42206 18564
rect 44706 18508 44716 18564
rect 44772 18508 46732 18564
rect 46788 18508 46798 18564
rect 51090 18508 51100 18564
rect 51156 18508 52500 18564
rect 24220 18452 24276 18508
rect 52444 18452 52500 18508
rect 15026 18396 15036 18452
rect 15092 18396 18060 18452
rect 18116 18396 18126 18452
rect 18274 18396 18284 18452
rect 18340 18396 19068 18452
rect 19124 18396 19134 18452
rect 23090 18396 23100 18452
rect 23156 18396 24276 18452
rect 27122 18396 27132 18452
rect 27188 18396 28588 18452
rect 28644 18396 28654 18452
rect 32162 18396 32172 18452
rect 32228 18396 33516 18452
rect 33572 18396 33582 18452
rect 35522 18396 35532 18452
rect 35588 18396 36876 18452
rect 36932 18396 36942 18452
rect 41346 18396 41356 18452
rect 41412 18396 42588 18452
rect 42644 18396 42654 18452
rect 44482 18396 44492 18452
rect 44548 18396 44558 18452
rect 51538 18396 51548 18452
rect 51604 18396 52220 18452
rect 52276 18396 52286 18452
rect 52444 18396 53452 18452
rect 53508 18396 53518 18452
rect 44492 18340 44548 18396
rect 17378 18284 17388 18340
rect 17444 18284 17948 18340
rect 18004 18284 18014 18340
rect 23762 18284 23772 18340
rect 23828 18284 23838 18340
rect 24434 18284 24444 18340
rect 24500 18284 27916 18340
rect 27972 18284 27982 18340
rect 28130 18284 28140 18340
rect 28196 18284 28700 18340
rect 28756 18284 28766 18340
rect 29138 18284 29148 18340
rect 29204 18284 32284 18340
rect 32340 18284 32350 18340
rect 35298 18284 35308 18340
rect 35364 18284 37884 18340
rect 37940 18284 38556 18340
rect 38612 18284 38622 18340
rect 40226 18284 40236 18340
rect 40292 18284 41804 18340
rect 41860 18284 41870 18340
rect 44492 18284 52556 18340
rect 52612 18284 52622 18340
rect 53218 18284 53228 18340
rect 53284 18284 54460 18340
rect 54516 18284 54526 18340
rect 23772 18228 23828 18284
rect 23772 18172 25004 18228
rect 25060 18172 43036 18228
rect 43092 18172 43596 18228
rect 43652 18172 43932 18228
rect 43988 18172 43998 18228
rect 51314 18172 51324 18228
rect 51380 18172 51772 18228
rect 51828 18172 51838 18228
rect 52322 18172 52332 18228
rect 52388 18172 53564 18228
rect 53620 18172 53630 18228
rect 54562 18172 54572 18228
rect 54628 18172 56476 18228
rect 56532 18172 56542 18228
rect 19842 18060 19852 18116
rect 19908 18060 24444 18116
rect 24500 18060 24510 18116
rect 27906 18060 27916 18116
rect 27972 18060 29148 18116
rect 29204 18060 29214 18116
rect 30818 18060 30828 18116
rect 30884 18060 31388 18116
rect 31444 18060 31454 18116
rect 45714 18060 45724 18116
rect 45780 18060 47852 18116
rect 47908 18060 47918 18116
rect 52108 18060 53788 18116
rect 53844 18060 53854 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 50642 17948 50652 18004
rect 50708 17948 51436 18004
rect 51492 17948 51502 18004
rect 52108 17892 52164 18060
rect 52556 17948 53116 18004
rect 53172 17948 53182 18004
rect 41458 17836 41468 17892
rect 41524 17836 44268 17892
rect 44324 17836 45276 17892
rect 45332 17836 45342 17892
rect 50978 17836 50988 17892
rect 51044 17836 52108 17892
rect 52164 17836 52174 17892
rect 52556 17780 52612 17948
rect 52770 17836 52780 17892
rect 52836 17836 54124 17892
rect 54180 17836 54190 17892
rect 21522 17724 21532 17780
rect 21588 17724 22316 17780
rect 22372 17724 30828 17780
rect 30884 17724 37212 17780
rect 37268 17724 37278 17780
rect 39778 17724 39788 17780
rect 39844 17724 40684 17780
rect 40740 17724 40750 17780
rect 50978 17724 50988 17780
rect 51044 17724 53620 17780
rect 53564 17668 53620 17724
rect 18946 17612 18956 17668
rect 19012 17612 22428 17668
rect 22484 17612 22494 17668
rect 28914 17612 28924 17668
rect 28980 17612 30492 17668
rect 30548 17612 30558 17668
rect 41682 17612 41692 17668
rect 41748 17612 44940 17668
rect 44996 17612 45006 17668
rect 47170 17612 47180 17668
rect 47236 17612 49868 17668
rect 49924 17612 50652 17668
rect 50708 17612 50718 17668
rect 53564 17612 54348 17668
rect 54404 17612 54414 17668
rect 49298 17500 49308 17556
rect 49364 17500 50428 17556
rect 50484 17500 50494 17556
rect 52882 17500 52892 17556
rect 52948 17500 53228 17556
rect 53284 17500 53294 17556
rect 14690 17388 14700 17444
rect 14756 17388 17500 17444
rect 17556 17388 17566 17444
rect 18274 17388 18284 17444
rect 18340 17388 19180 17444
rect 19236 17388 21196 17444
rect 21252 17388 21262 17444
rect 25330 17388 25340 17444
rect 25396 17388 28028 17444
rect 28084 17388 28094 17444
rect 35074 17388 35084 17444
rect 35140 17388 35980 17444
rect 36036 17388 36046 17444
rect 44258 17388 44268 17444
rect 44324 17388 46620 17444
rect 46676 17388 47404 17444
rect 47460 17388 47470 17444
rect 51090 17388 51100 17444
rect 51156 17388 51324 17444
rect 51380 17388 51390 17444
rect 52322 17388 52332 17444
rect 52388 17388 52556 17444
rect 52612 17388 53116 17444
rect 53172 17388 53182 17444
rect 53564 17332 53620 17612
rect 59200 17556 60000 17584
rect 55010 17500 55020 17556
rect 55076 17500 57820 17556
rect 57876 17500 57886 17556
rect 58146 17500 58156 17556
rect 58212 17500 60000 17556
rect 59200 17472 60000 17500
rect 17378 17276 17388 17332
rect 17444 17276 18396 17332
rect 18452 17276 18462 17332
rect 53554 17276 53564 17332
rect 53620 17276 53630 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 17714 17164 17724 17220
rect 17780 17164 18284 17220
rect 18340 17164 19684 17220
rect 28690 17164 28700 17220
rect 28756 17164 31500 17220
rect 31556 17164 31566 17220
rect 53442 17164 53452 17220
rect 53508 17164 55132 17220
rect 55188 17164 55198 17220
rect 19628 17108 19684 17164
rect 16818 17052 16828 17108
rect 16884 17052 18060 17108
rect 18116 17052 18508 17108
rect 18564 17052 18574 17108
rect 18722 17052 18732 17108
rect 18788 17052 18798 17108
rect 19628 17052 26908 17108
rect 28354 17052 28364 17108
rect 28420 17052 29708 17108
rect 29764 17052 30940 17108
rect 30996 17052 33180 17108
rect 33236 17052 33246 17108
rect 51986 17052 51996 17108
rect 52052 17052 52668 17108
rect 52724 17052 52734 17108
rect 18732 16996 18788 17052
rect 16706 16940 16716 16996
rect 16772 16940 18788 16996
rect 26852 16996 26908 17052
rect 26852 16940 27580 16996
rect 27636 16940 28140 16996
rect 28196 16940 35532 16996
rect 35588 16940 35598 16996
rect 35970 16940 35980 16996
rect 36036 16940 57036 16996
rect 57092 16940 57102 16996
rect 16828 16828 17612 16884
rect 17668 16828 19628 16884
rect 19684 16828 19694 16884
rect 51398 16828 51436 16884
rect 51492 16828 51502 16884
rect 51650 16828 51660 16884
rect 51716 16828 52892 16884
rect 52948 16828 52958 16884
rect 53778 16828 53788 16884
rect 53844 16828 55132 16884
rect 55188 16828 55198 16884
rect 16828 16772 16884 16828
rect 15922 16716 15932 16772
rect 15988 16716 16884 16772
rect 28242 16716 28252 16772
rect 28308 16716 28812 16772
rect 28868 16716 28878 16772
rect 31714 16716 31724 16772
rect 31780 16716 32508 16772
rect 32564 16716 32574 16772
rect 51762 16716 51772 16772
rect 51828 16716 52332 16772
rect 52388 16716 53340 16772
rect 53396 16716 53406 16772
rect 55234 16716 55244 16772
rect 55300 16716 57372 16772
rect 57428 16716 57438 16772
rect 38098 16604 38108 16660
rect 38164 16604 39116 16660
rect 39172 16604 39182 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 12898 16268 12908 16324
rect 12964 16268 21028 16324
rect 34962 16268 34972 16324
rect 35028 16268 37884 16324
rect 37940 16268 38332 16324
rect 38388 16268 41020 16324
rect 41076 16268 41086 16324
rect 14018 16156 14028 16212
rect 14084 16156 15932 16212
rect 15988 16156 15998 16212
rect 20972 16100 21028 16268
rect 21746 16156 21756 16212
rect 21812 16156 22428 16212
rect 22484 16156 22764 16212
rect 22820 16156 22830 16212
rect 24658 16156 24668 16212
rect 24724 16156 25228 16212
rect 25284 16156 35588 16212
rect 35532 16100 35588 16156
rect 20972 16044 32060 16100
rect 32116 16044 33628 16100
rect 33684 16044 33694 16100
rect 35522 16044 35532 16100
rect 35588 16044 36092 16100
rect 36148 16044 36158 16100
rect 18498 15932 18508 15988
rect 18564 15932 19292 15988
rect 19348 15932 27468 15988
rect 27524 15932 28140 15988
rect 28196 15932 28206 15988
rect 28354 15932 28364 15988
rect 28420 15932 29372 15988
rect 29428 15932 29438 15988
rect 34290 15932 34300 15988
rect 34356 15932 37772 15988
rect 37828 15932 37838 15988
rect 47730 15932 47740 15988
rect 47796 15932 50540 15988
rect 50596 15932 50606 15988
rect 22978 15820 22988 15876
rect 23044 15820 23660 15876
rect 23716 15820 23726 15876
rect 32498 15820 32508 15876
rect 32564 15820 33852 15876
rect 33908 15820 33918 15876
rect 37874 15820 37884 15876
rect 37940 15820 38556 15876
rect 38612 15820 38622 15876
rect 39554 15820 39564 15876
rect 39620 15820 41132 15876
rect 41188 15820 45052 15876
rect 45108 15820 45388 15876
rect 45444 15820 45454 15876
rect 45714 15820 45724 15876
rect 45780 15820 47180 15876
rect 47236 15820 48972 15876
rect 49028 15820 49420 15876
rect 49476 15820 50092 15876
rect 50148 15820 50158 15876
rect 32610 15708 32620 15764
rect 32676 15708 33068 15764
rect 33124 15708 37548 15764
rect 37604 15708 41916 15764
rect 41972 15708 41982 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 47282 15484 47292 15540
rect 47348 15484 48972 15540
rect 49028 15484 52108 15540
rect 52164 15484 52174 15540
rect 51762 15372 51772 15428
rect 51828 15372 52444 15428
rect 52500 15372 52510 15428
rect 38434 15260 38444 15316
rect 38500 15260 39564 15316
rect 39620 15260 39630 15316
rect 41010 15260 41020 15316
rect 41076 15260 41916 15316
rect 41972 15260 41982 15316
rect 45714 15260 45724 15316
rect 45780 15260 46844 15316
rect 46900 15260 46910 15316
rect 31714 15148 31724 15204
rect 31780 15148 32396 15204
rect 32452 15148 33740 15204
rect 33796 15148 33806 15204
rect 43652 15148 44716 15204
rect 44772 15148 46620 15204
rect 46676 15148 46686 15204
rect 50194 15148 50204 15204
rect 50260 15148 51548 15204
rect 51604 15148 52668 15204
rect 52724 15148 52734 15204
rect 43652 15092 43708 15148
rect 41682 15036 41692 15092
rect 41748 15036 42812 15092
rect 42868 15036 43708 15092
rect 50642 15036 50652 15092
rect 50708 15036 53564 15092
rect 53620 15036 54012 15092
rect 54068 15036 54460 15092
rect 54516 15036 54526 15092
rect 38612 14924 51100 14980
rect 51156 14924 51996 14980
rect 52052 14924 52062 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 38612 14756 38668 14924
rect 28466 14700 28476 14756
rect 28532 14700 38332 14756
rect 38388 14700 38668 14756
rect 49298 14700 49308 14756
rect 49364 14700 50540 14756
rect 50596 14700 50606 14756
rect 51202 14700 51212 14756
rect 51268 14700 52780 14756
rect 52836 14700 52846 14756
rect 23314 14588 23324 14644
rect 23380 14588 25788 14644
rect 25844 14588 26460 14644
rect 26516 14588 26526 14644
rect 26852 14588 27580 14644
rect 27636 14588 32620 14644
rect 32676 14588 32686 14644
rect 37090 14588 37100 14644
rect 37156 14588 40460 14644
rect 40516 14588 40526 14644
rect 41458 14588 41468 14644
rect 41524 14588 42588 14644
rect 42644 14588 42654 14644
rect 50418 14588 50428 14644
rect 50484 14588 50764 14644
rect 50820 14588 50830 14644
rect 18498 14476 18508 14532
rect 18564 14476 22204 14532
rect 22260 14476 22270 14532
rect 22642 14364 22652 14420
rect 22708 14364 26796 14420
rect 26852 14364 26908 14588
rect 41906 14476 41916 14532
rect 41972 14476 43036 14532
rect 43092 14476 44044 14532
rect 44100 14476 44716 14532
rect 44772 14476 44782 14532
rect 48066 14476 48076 14532
rect 48132 14476 50204 14532
rect 50260 14476 51212 14532
rect 51268 14476 51278 14532
rect 39554 14364 39564 14420
rect 39620 14364 40908 14420
rect 40964 14364 40974 14420
rect 48076 14308 48132 14476
rect 48290 14364 48300 14420
rect 48356 14364 51604 14420
rect 51762 14364 51772 14420
rect 51828 14364 53340 14420
rect 53396 14364 53406 14420
rect 54114 14364 54124 14420
rect 54180 14364 56588 14420
rect 56644 14364 56654 14420
rect 57250 14364 57260 14420
rect 57316 14364 57820 14420
rect 57876 14364 57886 14420
rect 51548 14308 51604 14364
rect 24322 14252 24332 14308
rect 24388 14252 27132 14308
rect 27188 14252 27198 14308
rect 41458 14252 41468 14308
rect 41524 14252 42700 14308
rect 42756 14252 42766 14308
rect 47618 14252 47628 14308
rect 47684 14252 48132 14308
rect 50530 14252 50540 14308
rect 50596 14252 50988 14308
rect 51044 14252 51054 14308
rect 51538 14252 51548 14308
rect 51604 14252 53116 14308
rect 53172 14252 53182 14308
rect 34066 14140 34076 14196
rect 34132 14140 34860 14196
rect 34916 14140 34926 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 18498 14028 18508 14084
rect 18564 14028 18732 14084
rect 18788 14028 18798 14084
rect 14690 13916 14700 13972
rect 14756 13916 20748 13972
rect 20804 13916 20814 13972
rect 21298 13916 21308 13972
rect 21364 13916 22204 13972
rect 22260 13916 22876 13972
rect 22932 13916 22942 13972
rect 28914 13916 28924 13972
rect 28980 13916 30044 13972
rect 30100 13916 35868 13972
rect 35924 13916 35934 13972
rect 41906 13916 41916 13972
rect 41972 13916 43260 13972
rect 43316 13916 43326 13972
rect 21074 13804 21084 13860
rect 21140 13804 22092 13860
rect 22148 13804 29372 13860
rect 29428 13804 29438 13860
rect 33740 13804 41132 13860
rect 41188 13804 41198 13860
rect 44930 13804 44940 13860
rect 44996 13804 47516 13860
rect 47572 13804 47582 13860
rect 52770 13804 52780 13860
rect 52836 13804 55244 13860
rect 55300 13804 55310 13860
rect 33740 13748 33796 13804
rect 18834 13692 18844 13748
rect 18900 13692 21756 13748
rect 21812 13692 21822 13748
rect 22642 13692 22652 13748
rect 22708 13692 23324 13748
rect 23380 13692 23390 13748
rect 30146 13692 30156 13748
rect 30212 13692 33068 13748
rect 33124 13692 33740 13748
rect 33796 13692 33806 13748
rect 38612 13692 39004 13748
rect 39060 13692 39070 13748
rect 47282 13692 47292 13748
rect 47348 13692 50204 13748
rect 50260 13692 50270 13748
rect 51874 13692 51884 13748
rect 51940 13692 52668 13748
rect 52724 13692 52734 13748
rect 16818 13580 16828 13636
rect 16884 13580 18732 13636
rect 18788 13580 19852 13636
rect 19908 13580 19918 13636
rect 20402 13580 20412 13636
rect 20468 13580 21196 13636
rect 21252 13580 23548 13636
rect 23604 13580 23614 13636
rect 30482 13580 30492 13636
rect 30548 13580 32060 13636
rect 32116 13580 32126 13636
rect 38612 13524 38668 13692
rect 42130 13580 42140 13636
rect 42196 13580 43708 13636
rect 43764 13580 50316 13636
rect 50372 13580 50382 13636
rect 52210 13580 52220 13636
rect 52276 13580 53116 13636
rect 53172 13580 53182 13636
rect 54450 13580 54460 13636
rect 54516 13580 55916 13636
rect 55972 13580 56700 13636
rect 56756 13580 57260 13636
rect 57316 13580 57326 13636
rect 17490 13468 17500 13524
rect 17556 13468 19516 13524
rect 19572 13468 23212 13524
rect 23268 13468 23278 13524
rect 24546 13468 24556 13524
rect 24612 13468 35308 13524
rect 35364 13468 35756 13524
rect 35812 13468 37212 13524
rect 37268 13468 37548 13524
rect 37604 13468 37884 13524
rect 37940 13468 38444 13524
rect 38500 13468 38668 13524
rect 40562 13468 40572 13524
rect 40628 13468 42476 13524
rect 42532 13468 42542 13524
rect 44594 13468 44604 13524
rect 44660 13468 44670 13524
rect 50866 13468 50876 13524
rect 50932 13468 51324 13524
rect 51380 13468 51390 13524
rect 44604 13412 44660 13468
rect 18274 13356 18284 13412
rect 18340 13356 19628 13412
rect 19684 13356 19694 13412
rect 38612 13356 39116 13412
rect 39172 13356 40012 13412
rect 40068 13356 40078 13412
rect 44146 13356 44156 13412
rect 44212 13356 44660 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 17826 13132 17836 13188
rect 17892 13132 18284 13188
rect 18340 13132 18350 13188
rect 19628 12964 19684 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 34962 13132 34972 13188
rect 35028 13132 35644 13188
rect 35700 13132 35710 13188
rect 29474 13020 29484 13076
rect 29540 13020 29932 13076
rect 29988 13020 29998 13076
rect 32162 13020 32172 13076
rect 32228 13020 33068 13076
rect 33124 13020 33134 13076
rect 33394 13020 33404 13076
rect 33460 13020 33964 13076
rect 34020 13020 34636 13076
rect 34692 13020 35084 13076
rect 35140 13020 35150 13076
rect 35858 13020 35868 13076
rect 35924 13020 37100 13076
rect 37156 13020 37166 13076
rect 38612 12964 38668 13356
rect 39218 13244 39228 13300
rect 39284 13244 39900 13300
rect 39956 13244 42364 13300
rect 42420 13244 49532 13300
rect 49588 13244 49598 13300
rect 17938 12908 17948 12964
rect 18004 12908 18732 12964
rect 18788 12908 18798 12964
rect 19628 12908 19852 12964
rect 19908 12908 19918 12964
rect 23762 12908 23772 12964
rect 23828 12908 34860 12964
rect 34916 12908 36316 12964
rect 36372 12908 38668 12964
rect 43362 12908 43372 12964
rect 43428 12908 43708 12964
rect 43764 12908 43774 12964
rect 22530 12796 22540 12852
rect 22596 12796 24108 12852
rect 24164 12796 24174 12852
rect 30370 12796 30380 12852
rect 30436 12796 31500 12852
rect 31556 12796 31566 12852
rect 32386 12796 32396 12852
rect 32452 12796 33292 12852
rect 33348 12796 33358 12852
rect 41122 12796 41132 12852
rect 41188 12796 42028 12852
rect 42084 12796 42588 12852
rect 42644 12796 42654 12852
rect 45490 12796 45500 12852
rect 45556 12796 47516 12852
rect 47572 12796 50204 12852
rect 50260 12796 50270 12852
rect 17826 12684 17836 12740
rect 17892 12684 19404 12740
rect 19460 12684 19470 12740
rect 24770 12684 24780 12740
rect 24836 12684 25228 12740
rect 25284 12684 27020 12740
rect 27076 12684 32228 12740
rect 33394 12684 33404 12740
rect 33460 12684 38780 12740
rect 38836 12684 39676 12740
rect 39732 12684 53004 12740
rect 53060 12684 53070 12740
rect 32172 12628 32228 12684
rect 20178 12572 20188 12628
rect 20244 12572 20860 12628
rect 20916 12572 28476 12628
rect 28532 12572 28542 12628
rect 32172 12572 35868 12628
rect 35924 12572 35934 12628
rect 44034 12572 44044 12628
rect 44100 12572 45276 12628
rect 45332 12572 47852 12628
rect 47908 12572 47918 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 18470 12460 18508 12516
rect 18564 12460 18574 12516
rect 26852 12460 30156 12516
rect 30212 12460 30222 12516
rect 35522 12460 35532 12516
rect 35588 12460 35980 12516
rect 36036 12460 36046 12516
rect 39666 12460 39676 12516
rect 39732 12460 42140 12516
rect 42196 12460 42206 12516
rect 26852 12404 26908 12460
rect 22418 12348 22428 12404
rect 22484 12348 23324 12404
rect 23380 12348 26908 12404
rect 27122 12348 27132 12404
rect 27188 12348 27580 12404
rect 27636 12348 28364 12404
rect 28420 12348 29484 12404
rect 29540 12348 30380 12404
rect 30436 12348 30446 12404
rect 31602 12348 31612 12404
rect 31668 12348 32508 12404
rect 32564 12348 32574 12404
rect 34514 12348 34524 12404
rect 34580 12348 35196 12404
rect 35252 12348 35262 12404
rect 38994 12348 39004 12404
rect 39060 12348 39340 12404
rect 39396 12348 39406 12404
rect 42354 12348 42364 12404
rect 42420 12348 42812 12404
rect 42868 12348 43484 12404
rect 43540 12348 49868 12404
rect 49924 12348 50652 12404
rect 50708 12348 51436 12404
rect 51492 12348 51502 12404
rect 44706 12236 44716 12292
rect 44772 12236 45612 12292
rect 45668 12236 45678 12292
rect 50306 12236 50316 12292
rect 50372 12236 52220 12292
rect 52276 12236 52668 12292
rect 52724 12236 52734 12292
rect 26852 12124 30156 12180
rect 30212 12124 33404 12180
rect 33460 12124 33470 12180
rect 26852 12068 26908 12124
rect 18274 12012 18284 12068
rect 18340 12012 21196 12068
rect 21252 12012 26908 12068
rect 27458 12012 27468 12068
rect 27524 12012 27916 12068
rect 27972 12012 34300 12068
rect 34356 12012 35084 12068
rect 35140 12012 38668 12068
rect 40226 12012 40236 12068
rect 40292 12012 42140 12068
rect 42196 12012 42206 12068
rect 38612 11956 38668 12012
rect 34626 11900 34636 11956
rect 34692 11900 37660 11956
rect 37716 11900 38108 11956
rect 38164 11900 38174 11956
rect 38612 11900 38836 11956
rect 38780 11844 38836 11900
rect 18722 11788 18732 11844
rect 18788 11788 20188 11844
rect 20244 11788 20254 11844
rect 38770 11788 38780 11844
rect 38836 11788 41692 11844
rect 41748 11788 50764 11844
rect 50820 11788 50988 11844
rect 51044 11788 51054 11844
rect 0 11732 800 11760
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 0 11676 2996 11732
rect 5842 11676 5852 11732
rect 5908 11676 5918 11732
rect 14466 11676 14476 11732
rect 14532 11676 17724 11732
rect 17780 11676 19516 11732
rect 19572 11676 19582 11732
rect 50082 11676 50092 11732
rect 50148 11676 54460 11732
rect 54516 11676 55580 11732
rect 55636 11676 55646 11732
rect 0 11648 800 11676
rect 2940 11620 2996 11676
rect 5852 11620 5908 11676
rect 2940 11564 5908 11620
rect 22642 11564 22652 11620
rect 22708 11564 32060 11620
rect 32116 11564 33964 11620
rect 34020 11564 34030 11620
rect 17266 11452 17276 11508
rect 17332 11452 18284 11508
rect 18340 11452 18732 11508
rect 18788 11452 18798 11508
rect 19170 11452 19180 11508
rect 19236 11452 21308 11508
rect 21364 11452 21374 11508
rect 29362 11452 29372 11508
rect 29428 11452 31836 11508
rect 31892 11452 31902 11508
rect 35522 11452 35532 11508
rect 35588 11452 38332 11508
rect 38388 11452 39452 11508
rect 39508 11452 39518 11508
rect 41010 11452 41020 11508
rect 41076 11452 43036 11508
rect 43092 11452 43102 11508
rect 47842 11452 47852 11508
rect 47908 11452 48860 11508
rect 48916 11452 48926 11508
rect 51650 11452 51660 11508
rect 51716 11452 54796 11508
rect 54852 11452 54862 11508
rect 27234 11340 27244 11396
rect 27300 11340 28252 11396
rect 28308 11340 29260 11396
rect 29316 11340 37940 11396
rect 52098 11340 52108 11396
rect 52164 11340 52892 11396
rect 52948 11340 52958 11396
rect 37884 11284 37940 11340
rect 33282 11228 33292 11284
rect 33348 11228 35532 11284
rect 35588 11228 35598 11284
rect 37874 11228 37884 11284
rect 37940 11228 38668 11284
rect 38724 11228 38734 11284
rect 15810 11116 15820 11172
rect 15876 11116 18844 11172
rect 18900 11116 18910 11172
rect 31826 11116 31836 11172
rect 31892 11116 33516 11172
rect 33572 11116 33582 11172
rect 20290 11004 20300 11060
rect 20356 11004 42252 11060
rect 42308 11004 42318 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 33506 10892 33516 10948
rect 33572 10892 39676 10948
rect 39732 10892 39742 10948
rect 26226 10780 26236 10836
rect 26292 10780 32620 10836
rect 32676 10780 32686 10836
rect 18386 10668 18396 10724
rect 18452 10668 21532 10724
rect 21588 10668 21598 10724
rect 26852 10668 27580 10724
rect 27636 10668 27646 10724
rect 31154 10668 31164 10724
rect 31220 10668 31724 10724
rect 31780 10668 46620 10724
rect 46676 10668 48300 10724
rect 48356 10668 48366 10724
rect 50866 10668 50876 10724
rect 50932 10668 51324 10724
rect 51380 10668 52444 10724
rect 52500 10668 52510 10724
rect 26852 10612 26908 10668
rect 59200 10612 60000 10640
rect 24546 10556 24556 10612
rect 24612 10556 25340 10612
rect 25396 10556 26908 10612
rect 43138 10556 43148 10612
rect 43204 10556 44268 10612
rect 44324 10556 44334 10612
rect 49858 10556 49868 10612
rect 49924 10556 51212 10612
rect 51268 10556 51278 10612
rect 58146 10556 58156 10612
rect 58212 10556 60000 10612
rect 59200 10528 60000 10556
rect 42242 10444 42252 10500
rect 42308 10444 50652 10500
rect 50708 10444 50718 10500
rect 18834 10332 18844 10388
rect 18900 10332 20076 10388
rect 20132 10332 20142 10388
rect 21634 10332 21644 10388
rect 21700 10332 22764 10388
rect 22820 10332 25340 10388
rect 25396 10332 25406 10388
rect 42130 10332 42140 10388
rect 42196 10332 51996 10388
rect 52052 10332 52062 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 24658 10108 24668 10164
rect 24724 10108 27356 10164
rect 27412 10108 27422 10164
rect 38994 10108 39004 10164
rect 39060 10108 40236 10164
rect 40292 10108 41804 10164
rect 41860 10108 43036 10164
rect 43092 10108 46844 10164
rect 46900 10108 46910 10164
rect 17826 9996 17836 10052
rect 17892 9996 19516 10052
rect 19572 9996 19582 10052
rect 31042 9996 31052 10052
rect 31108 9996 33404 10052
rect 33460 9996 33470 10052
rect 50194 9996 50204 10052
rect 50260 9996 50988 10052
rect 51044 9996 51054 10052
rect 21746 9884 21756 9940
rect 21812 9884 22204 9940
rect 22260 9884 25004 9940
rect 25060 9884 25070 9940
rect 29698 9884 29708 9940
rect 29764 9884 30492 9940
rect 30548 9884 30558 9940
rect 31154 9884 31164 9940
rect 31220 9884 32284 9940
rect 32340 9884 33292 9940
rect 33348 9884 33358 9940
rect 33730 9884 33740 9940
rect 33796 9884 34580 9940
rect 42242 9884 42252 9940
rect 42308 9884 42588 9940
rect 42644 9884 42654 9940
rect 51538 9884 51548 9940
rect 51604 9884 52668 9940
rect 52724 9884 52734 9940
rect 34524 9828 34580 9884
rect 42588 9828 42644 9884
rect 17266 9772 17276 9828
rect 17332 9772 17948 9828
rect 18004 9772 18732 9828
rect 18788 9772 19180 9828
rect 19236 9772 19246 9828
rect 26562 9772 26572 9828
rect 26628 9772 27020 9828
rect 27076 9772 28028 9828
rect 28084 9772 28094 9828
rect 31378 9772 31388 9828
rect 31444 9772 31836 9828
rect 31892 9772 31902 9828
rect 33170 9772 33180 9828
rect 33236 9772 34076 9828
rect 34132 9772 34142 9828
rect 34514 9772 34524 9828
rect 34580 9772 35644 9828
rect 35700 9772 35710 9828
rect 36082 9772 36092 9828
rect 36148 9772 37100 9828
rect 37156 9772 37166 9828
rect 42588 9772 43820 9828
rect 43876 9772 43886 9828
rect 19282 9660 19292 9716
rect 19348 9660 19358 9716
rect 19842 9660 19852 9716
rect 19908 9660 23436 9716
rect 23492 9660 23502 9716
rect 27682 9660 27692 9716
rect 27748 9660 28588 9716
rect 28644 9660 29932 9716
rect 29988 9660 29998 9716
rect 32722 9660 32732 9716
rect 32788 9660 33292 9716
rect 33348 9660 33358 9716
rect 36530 9660 36540 9716
rect 36596 9660 40348 9716
rect 40404 9660 40414 9716
rect 42438 9660 42476 9716
rect 42532 9660 42542 9716
rect 51650 9660 51660 9716
rect 51716 9660 54796 9716
rect 54852 9660 54862 9716
rect 19292 9604 19348 9660
rect 15810 9548 15820 9604
rect 15876 9548 18844 9604
rect 18900 9548 18910 9604
rect 19292 9548 20412 9604
rect 20468 9548 21420 9604
rect 21476 9548 21486 9604
rect 26674 9548 26684 9604
rect 26740 9548 27580 9604
rect 27636 9548 27646 9604
rect 30034 9548 30044 9604
rect 30100 9548 30604 9604
rect 30660 9548 30670 9604
rect 29698 9436 29708 9492
rect 29764 9436 37324 9492
rect 37380 9436 37390 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 33282 9324 33292 9380
rect 33348 9324 38668 9380
rect 38612 9268 38668 9324
rect 18162 9212 18172 9268
rect 18228 9212 18732 9268
rect 18788 9212 18798 9268
rect 18946 9212 18956 9268
rect 19012 9212 19628 9268
rect 19684 9212 19694 9268
rect 32834 9212 32844 9268
rect 32900 9212 33852 9268
rect 33908 9212 33918 9268
rect 38612 9212 43596 9268
rect 43652 9212 43662 9268
rect 51314 9212 51324 9268
rect 51380 9212 51996 9268
rect 52052 9212 52062 9268
rect 34402 9100 34412 9156
rect 34468 9100 35532 9156
rect 35588 9100 37660 9156
rect 37716 9100 39228 9156
rect 39284 9100 39788 9156
rect 39844 9100 39854 9156
rect 42466 9100 42476 9156
rect 42532 9100 42812 9156
rect 42868 9100 43484 9156
rect 43540 9100 43550 9156
rect 47170 9100 47180 9156
rect 47236 9100 49980 9156
rect 50036 9100 50046 9156
rect 18274 8988 18284 9044
rect 18340 8988 18956 9044
rect 19012 8988 19516 9044
rect 19572 8988 19582 9044
rect 35074 8988 35084 9044
rect 35140 8988 35868 9044
rect 35924 8988 35934 9044
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 22418 8428 22428 8484
rect 22484 8428 25452 8484
rect 25508 8428 26572 8484
rect 26628 8428 26638 8484
rect 31948 8428 34188 8484
rect 34244 8428 34254 8484
rect 50418 8428 50428 8484
rect 50484 8428 50494 8484
rect 31948 8372 32004 8428
rect 50428 8372 50484 8428
rect 30930 8316 30940 8372
rect 30996 8316 32004 8372
rect 32498 8316 32508 8372
rect 32564 8316 38668 8372
rect 44930 8316 44940 8372
rect 44996 8316 45612 8372
rect 45668 8316 45678 8372
rect 47394 8316 47404 8372
rect 47460 8316 51212 8372
rect 51268 8316 51278 8372
rect 38612 8260 38668 8316
rect 26852 8036 26908 8260
rect 26964 8204 26974 8260
rect 27346 8204 27356 8260
rect 27412 8204 36316 8260
rect 36372 8204 36382 8260
rect 38612 8204 42140 8260
rect 42196 8204 45724 8260
rect 45780 8204 45790 8260
rect 46386 8204 46396 8260
rect 46452 8204 47516 8260
rect 47572 8204 47582 8260
rect 48850 8204 48860 8260
rect 48916 8204 50428 8260
rect 50484 8204 51324 8260
rect 51380 8204 51390 8260
rect 31154 8092 31164 8148
rect 31220 8092 31612 8148
rect 31668 8092 31678 8148
rect 19282 7980 19292 8036
rect 19348 7980 20300 8036
rect 20356 7980 20366 8036
rect 26338 7980 26348 8036
rect 26404 7980 26908 8036
rect 29810 7980 29820 8036
rect 29876 7980 30716 8036
rect 30772 7980 30782 8036
rect 33954 7980 33964 8036
rect 34020 7980 34972 8036
rect 35028 7980 35038 8036
rect 36316 7924 36372 8204
rect 45724 8148 45780 8204
rect 36754 8092 36764 8148
rect 36820 8092 42924 8148
rect 42980 8092 42990 8148
rect 45724 8092 46620 8148
rect 46676 8092 46686 8148
rect 47842 8092 47852 8148
rect 47908 8092 48636 8148
rect 48692 8092 48702 8148
rect 49830 8092 49868 8148
rect 49924 8092 49934 8148
rect 38994 7980 39004 8036
rect 39060 7980 39676 8036
rect 39732 7980 39742 8036
rect 43698 7980 43708 8036
rect 43764 7980 46172 8036
rect 46228 7980 46238 8036
rect 47170 7980 47180 8036
rect 47236 7980 48524 8036
rect 48580 7980 49532 8036
rect 49588 7980 49598 8036
rect 18834 7868 18844 7924
rect 18900 7868 19404 7924
rect 19460 7868 19470 7924
rect 36316 7868 39172 7924
rect 41458 7868 41468 7924
rect 41524 7868 49308 7924
rect 49364 7868 49374 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 28018 7756 28028 7812
rect 28084 7756 38668 7812
rect 38612 7700 38668 7756
rect 30930 7644 30940 7700
rect 30996 7644 31500 7700
rect 31556 7644 31566 7700
rect 35522 7644 35532 7700
rect 35588 7644 36092 7700
rect 36148 7644 37436 7700
rect 37492 7644 37502 7700
rect 38612 7644 38892 7700
rect 38948 7644 38958 7700
rect 19058 7532 19068 7588
rect 19124 7532 19628 7588
rect 19684 7532 19694 7588
rect 33842 7532 33852 7588
rect 33908 7532 35644 7588
rect 35700 7532 36428 7588
rect 36484 7532 36494 7588
rect 39116 7476 39172 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 39554 7756 39564 7812
rect 39620 7756 47180 7812
rect 47236 7756 47246 7812
rect 40002 7644 40012 7700
rect 40068 7644 41468 7700
rect 41524 7644 41534 7700
rect 40114 7532 40124 7588
rect 40180 7532 41692 7588
rect 41748 7532 43820 7588
rect 43876 7532 43886 7588
rect 49868 7532 50652 7588
rect 50708 7532 51548 7588
rect 51604 7532 51614 7588
rect 49868 7476 49924 7532
rect 19394 7420 19404 7476
rect 19460 7420 21532 7476
rect 21588 7420 21598 7476
rect 24098 7420 24108 7476
rect 24164 7420 27244 7476
rect 27300 7420 28140 7476
rect 28196 7420 28206 7476
rect 34178 7420 34188 7476
rect 34244 7420 35420 7476
rect 35476 7420 35486 7476
rect 38098 7420 38108 7476
rect 38164 7420 38668 7476
rect 38724 7420 38734 7476
rect 39106 7420 39116 7476
rect 39172 7420 39900 7476
rect 39956 7420 40796 7476
rect 40852 7420 40862 7476
rect 41234 7420 41244 7476
rect 41300 7420 41804 7476
rect 41860 7420 41870 7476
rect 49858 7420 49868 7476
rect 49924 7420 49934 7476
rect 50092 7420 51436 7476
rect 51492 7420 51502 7476
rect 35420 7364 35476 7420
rect 50092 7364 50148 7420
rect 27010 7308 27020 7364
rect 27076 7308 27692 7364
rect 27748 7308 31724 7364
rect 31780 7308 31790 7364
rect 35420 7308 38220 7364
rect 38276 7308 39340 7364
rect 39396 7308 39406 7364
rect 48626 7308 48636 7364
rect 48692 7308 50148 7364
rect 50204 7308 50876 7364
rect 50932 7308 50942 7364
rect 51538 7308 51548 7364
rect 51604 7308 52444 7364
rect 52500 7308 52510 7364
rect 19282 7196 19292 7252
rect 19348 7196 19852 7252
rect 19908 7196 20748 7252
rect 20804 7196 21420 7252
rect 21476 7196 21486 7252
rect 23762 7196 23772 7252
rect 23828 7196 25788 7252
rect 25844 7196 26796 7252
rect 26852 7196 26862 7252
rect 34962 7196 34972 7252
rect 35028 7196 35980 7252
rect 36036 7196 36046 7252
rect 39666 7196 39676 7252
rect 39732 7196 49420 7252
rect 49476 7196 49486 7252
rect 50204 7140 50260 7308
rect 43250 7084 43260 7140
rect 43316 7084 50260 7140
rect 50372 7196 50652 7252
rect 50708 7196 50718 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 20514 6972 20524 7028
rect 20580 6972 21308 7028
rect 21364 6972 22764 7028
rect 22820 6972 23548 7028
rect 23604 6972 23614 7028
rect 37986 6972 37996 7028
rect 38052 6972 38780 7028
rect 38836 6972 38846 7028
rect 23874 6860 23884 6916
rect 23940 6860 24444 6916
rect 24500 6860 24510 6916
rect 38994 6860 39004 6916
rect 39060 6860 40796 6916
rect 40852 6860 41300 6916
rect 41244 6804 41300 6860
rect 50372 6804 50428 7196
rect 17714 6748 17724 6804
rect 17780 6748 18620 6804
rect 18676 6748 18686 6804
rect 20178 6748 20188 6804
rect 20244 6748 22204 6804
rect 22260 6748 22270 6804
rect 23202 6748 23212 6804
rect 23268 6748 24332 6804
rect 24388 6748 24398 6804
rect 41234 6748 41244 6804
rect 41300 6748 41310 6804
rect 42028 6748 43260 6804
rect 43316 6748 43326 6804
rect 48738 6748 48748 6804
rect 48804 6748 49812 6804
rect 49970 6748 49980 6804
rect 50036 6748 50428 6804
rect 51538 6748 51548 6804
rect 51604 6748 52668 6804
rect 52724 6748 52734 6804
rect 42028 6692 42084 6748
rect 49756 6692 49812 6748
rect 15474 6636 15484 6692
rect 15540 6636 17500 6692
rect 17556 6636 17566 6692
rect 20626 6636 20636 6692
rect 20692 6636 21308 6692
rect 21364 6636 21374 6692
rect 21980 6636 24108 6692
rect 24164 6636 26236 6692
rect 26292 6636 27244 6692
rect 27300 6636 27310 6692
rect 30482 6636 30492 6692
rect 30548 6636 31836 6692
rect 31892 6636 32396 6692
rect 32452 6636 32462 6692
rect 39330 6636 39340 6692
rect 39396 6636 40236 6692
rect 40292 6636 40302 6692
rect 40562 6636 40572 6692
rect 40628 6636 42084 6692
rect 43026 6636 43036 6692
rect 43092 6636 45164 6692
rect 45220 6636 45230 6692
rect 46498 6636 46508 6692
rect 46564 6636 47292 6692
rect 47348 6636 47358 6692
rect 49746 6636 49756 6692
rect 49812 6636 49822 6692
rect 52546 6636 52556 6692
rect 52612 6636 54796 6692
rect 54852 6636 54862 6692
rect 21980 6580 22036 6636
rect 40572 6580 40628 6636
rect 16146 6524 16156 6580
rect 16212 6524 17388 6580
rect 17444 6524 17454 6580
rect 18946 6524 18956 6580
rect 19012 6524 21980 6580
rect 22036 6524 22046 6580
rect 23314 6524 23324 6580
rect 23380 6524 25228 6580
rect 25284 6524 25294 6580
rect 26562 6524 26572 6580
rect 26628 6524 27188 6580
rect 30258 6524 30268 6580
rect 30324 6524 31948 6580
rect 32004 6524 32014 6580
rect 32274 6524 32284 6580
rect 32340 6524 32620 6580
rect 32676 6524 32686 6580
rect 38546 6524 38556 6580
rect 38612 6524 40628 6580
rect 41794 6524 41804 6580
rect 41860 6524 49420 6580
rect 49476 6524 50428 6580
rect 50484 6524 50494 6580
rect 26572 6468 26628 6524
rect 19170 6412 19180 6468
rect 19236 6412 20412 6468
rect 20468 6412 21756 6468
rect 21812 6412 21822 6468
rect 22194 6412 22204 6468
rect 22260 6412 23660 6468
rect 23716 6412 23726 6468
rect 23874 6412 23884 6468
rect 23940 6412 26628 6468
rect 27132 6468 27188 6524
rect 27132 6412 27524 6468
rect 43810 6412 43820 6468
rect 43876 6412 48188 6468
rect 48244 6412 48254 6468
rect 50372 6412 54012 6468
rect 54068 6412 54078 6468
rect 27468 6356 27524 6412
rect 43820 6356 43876 6412
rect 50372 6356 50428 6412
rect 20290 6300 20300 6356
rect 20356 6300 24220 6356
rect 24276 6300 24286 6356
rect 26002 6300 26012 6356
rect 26068 6300 27300 6356
rect 27468 6300 33628 6356
rect 33684 6300 33694 6356
rect 40002 6300 40012 6356
rect 40068 6300 40348 6356
rect 40404 6300 43876 6356
rect 46610 6300 46620 6356
rect 46676 6300 50428 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 27244 6244 27300 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 25106 6188 25116 6244
rect 25172 6188 26908 6244
rect 27244 6188 28140 6244
rect 28196 6188 28206 6244
rect 31266 6188 31276 6244
rect 31332 6188 32060 6244
rect 32116 6188 43932 6244
rect 43988 6188 43998 6244
rect 26852 6132 26908 6188
rect 17490 6076 17500 6132
rect 17556 6076 18396 6132
rect 18452 6076 18462 6132
rect 26852 6076 27580 6132
rect 27636 6076 30716 6132
rect 30772 6076 30782 6132
rect 45042 6076 45052 6132
rect 45108 6076 46732 6132
rect 46788 6076 46798 6132
rect 48402 6076 48412 6132
rect 48468 6076 50428 6132
rect 50484 6076 51212 6132
rect 51268 6076 51278 6132
rect 30818 5964 30828 6020
rect 30884 5964 30894 6020
rect 46498 5964 46508 6020
rect 46564 5964 47068 6020
rect 47124 5964 47134 6020
rect 21186 5852 21196 5908
rect 21252 5852 21980 5908
rect 22036 5852 22046 5908
rect 30828 5572 30884 5964
rect 49830 5852 49868 5908
rect 49924 5852 49934 5908
rect 32162 5628 32172 5684
rect 32228 5628 44940 5684
rect 44996 5628 45276 5684
rect 45332 5628 45342 5684
rect 21746 5516 21756 5572
rect 21812 5516 26908 5572
rect 30818 5516 30828 5572
rect 30884 5516 30894 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 26852 5460 26908 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 26852 5404 29372 5460
rect 29428 5404 31500 5460
rect 31556 5404 31566 5460
rect 37650 5292 37660 5348
rect 37716 5292 39452 5348
rect 39508 5292 39900 5348
rect 39956 5292 40908 5348
rect 40964 5292 41244 5348
rect 41300 5292 41310 5348
rect 18386 5180 18396 5236
rect 18452 5180 21420 5236
rect 21476 5180 21486 5236
rect 29698 5180 29708 5236
rect 29764 5180 30940 5236
rect 30996 5180 31006 5236
rect 34514 5180 34524 5236
rect 34580 5180 35644 5236
rect 35700 5180 35710 5236
rect 44594 5180 44604 5236
rect 44660 5180 45500 5236
rect 45556 5180 46508 5236
rect 46564 5180 46574 5236
rect 48850 5180 48860 5236
rect 48916 5180 49868 5236
rect 49924 5180 49934 5236
rect 30818 5068 30828 5124
rect 30884 5068 32060 5124
rect 32116 5068 32126 5124
rect 38210 5068 38220 5124
rect 38276 5068 39116 5124
rect 39172 5068 39182 5124
rect 47058 5068 47068 5124
rect 47124 5068 50316 5124
rect 50372 5012 50428 5124
rect 50372 4956 53340 5012
rect 53396 4956 55468 5012
rect 55524 4956 55534 5012
rect 51314 4844 51324 4900
rect 51380 4844 52668 4900
rect 52724 4844 52734 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 28578 4508 28588 4564
rect 28644 4508 30492 4564
rect 30548 4508 30558 4564
rect 46946 4508 46956 4564
rect 47012 4508 48748 4564
rect 48804 4508 48814 4564
rect 28588 4340 28644 4508
rect 40786 4396 40796 4452
rect 40852 4396 41692 4452
rect 41748 4396 41758 4452
rect 25330 4284 25340 4340
rect 25396 4284 28644 4340
rect 54002 4284 54012 4340
rect 54068 4284 57596 4340
rect 57652 4284 57662 4340
rect 46050 4172 46060 4228
rect 46116 4172 47068 4228
rect 47124 4172 48524 4228
rect 48580 4172 48590 4228
rect 57362 4172 57372 4228
rect 57428 4172 58156 4228
rect 58212 4172 58222 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 59200 3668 60000 3696
rect 58146 3612 58156 3668
rect 58212 3612 60000 3668
rect 59200 3584 60000 3612
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 49084 63084 49140 63140
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 49084 60956 49140 61012
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4284 51100 4340 51156
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 4284 50316 4340 50372
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 14252 45164 14308 45220
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 14924 42588 14980 42644
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 13468 40348 13524 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 14924 39900 14980 39956
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 46060 38668 46116 38724
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 46060 37996 46116 38052
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 22092 33180 22148 33236
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 14252 31836 14308 31892
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 22092 30716 22148 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 13468 29148 13524 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 25564 26684 25620 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 25564 26236 25620 26292
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 25564 24892 25620 24948
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 38668 19516 38724 19572
rect 38668 19180 38724 19236
rect 50988 18956 51044 19012
rect 51436 18956 51492 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 50988 17836 51044 17892
rect 51324 17388 51380 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 51436 16828 51492 16884
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 18508 14028 18564 14084
rect 51324 13468 51380 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 18508 12460 18564 12516
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 42476 9660 42532 9716
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 42476 9100 42532 9156
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 49868 8092 49924 8148
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 49868 5852 49924 5908
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 66668 4768 66700
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4284 51156 4340 51166
rect 4284 50372 4340 51100
rect 4284 50306 4340 50316
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 19808 65884 20128 66700
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 14252 45220 14308 45230
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 13468 40404 13524 40414
rect 13468 29204 13524 40348
rect 14252 31892 14308 45164
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 14924 42644 14980 42654
rect 14924 39956 14980 42588
rect 14924 39890 14980 39900
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 14252 31826 14308 31836
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 35168 66668 35488 66700
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 50528 65884 50848 66700
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 49084 63140 49140 63150
rect 49084 61012 49140 63084
rect 49084 60946 49140 60956
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 46060 38724 46116 38734
rect 46060 38052 46116 38668
rect 46060 37986 46116 37996
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 13468 29138 13524 29148
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 22092 33236 22148 33246
rect 22092 30772 22148 33180
rect 22092 30706 22148 30716
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 25564 26740 25620 26750
rect 25564 26292 25620 26684
rect 25564 24948 25620 26236
rect 25564 24882 25620 24892
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 18508 14084 18564 14094
rect 18508 12516 18564 14028
rect 18508 12450 18564 12460
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 35168 18060 35488 19572
rect 38668 19572 38724 19582
rect 38668 19236 38724 19516
rect 38668 19170 38724 19180
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50988 19012 51044 19022
rect 50988 17892 51044 18956
rect 50988 17826 51044 17836
rect 51436 19012 51492 19022
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 51324 17444 51380 17454
rect 51324 13524 51380 17388
rect 51436 16884 51492 18956
rect 51436 16818 51492 16828
rect 51324 13458 51380 13468
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 42476 9716 42532 9726
rect 42476 9156 42532 9660
rect 42476 9090 42532 9100
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 49868 8148 49924 8158
rect 49868 5908 49924 8092
rect 49868 5842 49924 5852
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1260_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1261_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23744 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1263_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1264_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1265_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26992 0 -1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1266_
timestamp 1698431365
transform -1 0 24192 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1267_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1268_
timestamp 1698431365
transform -1 0 23520 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1269_
timestamp 1698431365
transform 1 0 21952 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1270_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25760 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1271_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22400 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1272_
timestamp 1698431365
transform 1 0 27328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1273_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28336 0 -1 40768
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1274_
timestamp 1698431365
transform 1 0 23968 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1275_
timestamp 1698431365
transform -1 0 24864 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1276_
timestamp 1698431365
transform -1 0 24864 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1277_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1278_
timestamp 1698431365
transform 1 0 22848 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1279_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28336 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1280_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1281_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1282_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31472 0 1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1283_
timestamp 1698431365
transform -1 0 31472 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1284_
timestamp 1698431365
transform 1 0 34496 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1285_
timestamp 1698431365
transform -1 0 37744 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1286_
timestamp 1698431365
transform -1 0 35840 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1287_
timestamp 1698431365
transform 1 0 38080 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1288_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1289_
timestamp 1698431365
transform -1 0 41664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1290_
timestamp 1698431365
transform -1 0 38304 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1291_
timestamp 1698431365
transform -1 0 36288 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1292_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35056 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1293_
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1294_
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1295_
timestamp 1698431365
transform 1 0 34384 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1296_
timestamp 1698431365
transform -1 0 34496 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1297_
timestamp 1698431365
transform -1 0 38304 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1298_
timestamp 1698431365
transform -1 0 36512 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1299_
timestamp 1698431365
transform -1 0 35280 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1300_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33936 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1301_
timestamp 1698431365
transform -1 0 21056 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1302_
timestamp 1698431365
transform 1 0 20944 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1303_
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1304_
timestamp 1698431365
transform -1 0 19152 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1305_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19600 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1306_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18368 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1307_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16352 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1308_
timestamp 1698431365
transform 1 0 15344 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1309_
timestamp 1698431365
transform 1 0 20944 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1310_
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1311_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16352 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1312_
timestamp 1698431365
transform 1 0 16912 0 1 37632
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1313_
timestamp 1698431365
transform 1 0 20160 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1314_
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1315_
timestamp 1698431365
transform 1 0 19376 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1316_
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1317_
timestamp 1698431365
transform -1 0 16576 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1318_
timestamp 1698431365
transform 1 0 7056 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1319_
timestamp 1698431365
transform 1 0 7168 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1320_
timestamp 1698431365
transform -1 0 8512 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1321_
timestamp 1698431365
transform -1 0 10976 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1322_
timestamp 1698431365
transform 1 0 7728 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1323_
timestamp 1698431365
transform 1 0 9408 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1324_
timestamp 1698431365
transform -1 0 11424 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1325_
timestamp 1698431365
transform 1 0 10864 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1326_
timestamp 1698431365
transform 1 0 7616 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1327_
timestamp 1698431365
transform -1 0 12432 0 -1 31360
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1328_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1329_
timestamp 1698431365
transform -1 0 12768 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1330_
timestamp 1698431365
transform -1 0 11536 0 1 31360
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1331_
timestamp 1698431365
transform 1 0 6720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1332_
timestamp 1698431365
transform 1 0 11424 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1333_
timestamp 1698431365
transform 1 0 13776 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1334_
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1335_
timestamp 1698431365
transform -1 0 13104 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1336_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11984 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1337_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1338_
timestamp 1698431365
transform 1 0 33264 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1339_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35392 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1340_
timestamp 1698431365
transform 1 0 34496 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1341_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38192 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37408 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1343_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24416 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1344_
timestamp 1698431365
transform 1 0 23856 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1345_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27664 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1346_
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1347_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1348_
timestamp 1698431365
transform -1 0 39312 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1349_
timestamp 1698431365
transform -1 0 38080 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1350_
timestamp 1698431365
transform -1 0 36624 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1351_
timestamp 1698431365
transform -1 0 35840 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1352_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1353_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37520 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1354_
timestamp 1698431365
transform -1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1355_
timestamp 1698431365
transform -1 0 19376 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1356_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20720 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1358_
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1359_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1360_
timestamp 1698431365
transform 1 0 16016 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1361_
timestamp 1698431365
transform 1 0 17360 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1362_
timestamp 1698431365
transform -1 0 12768 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1363_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1364_
timestamp 1698431365
transform -1 0 14224 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1365_
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1366_
timestamp 1698431365
transform 1 0 11648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1367_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14784 0 -1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1368_
timestamp 1698431365
transform 1 0 11536 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1369_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1370_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10752 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1371_
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1372_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37968 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1373_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37408 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1374_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38080 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1375_
timestamp 1698431365
transform 1 0 37408 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1376_
timestamp 1698431365
transform -1 0 11200 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1377_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1378_
timestamp 1698431365
transform -1 0 14000 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1379_
timestamp 1698431365
transform -1 0 14896 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1380_
timestamp 1698431365
transform -1 0 15120 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1381_
timestamp 1698431365
transform -1 0 14784 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1382_
timestamp 1698431365
transform -1 0 10864 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1383_
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1384_
timestamp 1698431365
transform 1 0 6496 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1385_
timestamp 1698431365
transform 1 0 7168 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1386_
timestamp 1698431365
transform -1 0 8400 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1387_
timestamp 1698431365
transform -1 0 11536 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1388_
timestamp 1698431365
transform -1 0 11312 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1389_
timestamp 1698431365
transform 1 0 12208 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1390_
timestamp 1698431365
transform -1 0 13104 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1391_
timestamp 1698431365
transform 1 0 18704 0 1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1392_
timestamp 1698431365
transform -1 0 20944 0 -1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1393_
timestamp 1698431365
transform 1 0 19264 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1394_
timestamp 1698431365
transform -1 0 20272 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1395_
timestamp 1698431365
transform -1 0 15344 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1396_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1397_
timestamp 1698431365
transform 1 0 15792 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1398_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15344 0 1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1399_
timestamp 1698431365
transform 1 0 15120 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1400_
timestamp 1698431365
transform -1 0 37296 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1401_
timestamp 1698431365
transform 1 0 34384 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1402_
timestamp 1698431365
transform -1 0 33264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1403_
timestamp 1698431365
transform 1 0 36848 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1404_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1405_
timestamp 1698431365
transform 1 0 31360 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1406_
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1407_
timestamp 1698431365
transform 1 0 22848 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1408_
timestamp 1698431365
transform -1 0 28000 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1409_
timestamp 1698431365
transform 1 0 25760 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1410_
timestamp 1698431365
transform -1 0 25984 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1411_
timestamp 1698431365
transform -1 0 28784 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1412_
timestamp 1698431365
transform -1 0 27888 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1413_
timestamp 1698431365
transform 1 0 24640 0 1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1414_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27104 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1415_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17360 0 -1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1416_
timestamp 1698431365
transform 1 0 35616 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1417_
timestamp 1698431365
transform 1 0 36176 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1418_
timestamp 1698431365
transform 1 0 38304 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1419_
timestamp 1698431365
transform 1 0 17136 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1420_
timestamp 1698431365
transform -1 0 26096 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1421_
timestamp 1698431365
transform -1 0 24976 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1422_
timestamp 1698431365
transform -1 0 24864 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1423_
timestamp 1698431365
transform -1 0 24864 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1424_
timestamp 1698431365
transform -1 0 36960 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1426_
timestamp 1698431365
transform -1 0 36176 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1427_
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1428_
timestamp 1698431365
transform -1 0 24416 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1429_
timestamp 1698431365
transform 1 0 23744 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1698431365
transform -1 0 26320 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1431_
timestamp 1698431365
transform -1 0 28224 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1432_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1433_
timestamp 1698431365
transform -1 0 28336 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1434_
timestamp 1698431365
transform -1 0 15568 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1435_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1436_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1437_
timestamp 1698431365
transform 1 0 14112 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1438_
timestamp 1698431365
transform 1 0 15568 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1439_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1440_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 42336
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1441_
timestamp 1698431365
transform 1 0 14224 0 -1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1442_
timestamp 1698431365
transform -1 0 14000 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1443_
timestamp 1698431365
transform -1 0 15344 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1444_
timestamp 1698431365
transform 1 0 15344 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1445_
timestamp 1698431365
transform 1 0 17024 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1446_
timestamp 1698431365
transform 1 0 25536 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1447_
timestamp 1698431365
transform 1 0 34272 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1448_
timestamp 1698431365
transform 1 0 34608 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1449_
timestamp 1698431365
transform 1 0 35952 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1450_
timestamp 1698431365
transform 1 0 25648 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1451_
timestamp 1698431365
transform 1 0 28224 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1452_
timestamp 1698431365
transform -1 0 27776 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698431365
transform 1 0 28112 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1454_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1455_
timestamp 1698431365
transform 1 0 26768 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1456_
timestamp 1698431365
transform 1 0 29568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1457_
timestamp 1698431365
transform -1 0 31360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1458_
timestamp 1698431365
transform -1 0 33264 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1459_
timestamp 1698431365
transform 1 0 31136 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1460_
timestamp 1698431365
transform 1 0 14112 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1461_
timestamp 1698431365
transform 1 0 9632 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1462_
timestamp 1698431365
transform 1 0 13552 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1463_
timestamp 1698431365
transform 1 0 14224 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1464_
timestamp 1698431365
transform -1 0 14224 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1465_
timestamp 1698431365
transform -1 0 13104 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1466_
timestamp 1698431365
transform 1 0 13216 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1467_
timestamp 1698431365
transform 1 0 16016 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1468_
timestamp 1698431365
transform 1 0 14448 0 1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1469_
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1470_
timestamp 1698431365
transform 1 0 34496 0 1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1471_
timestamp 1698431365
transform 1 0 37520 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1472_
timestamp 1698431365
transform 1 0 38752 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1473_
timestamp 1698431365
transform 1 0 34720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1474_
timestamp 1698431365
transform 1 0 36064 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1475_
timestamp 1698431365
transform -1 0 31808 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1476_
timestamp 1698431365
transform 1 0 31808 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1477_
timestamp 1698431365
transform 1 0 32592 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1478_
timestamp 1698431365
transform -1 0 33712 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28336 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1480_
timestamp 1698431365
transform 1 0 29232 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1481_
timestamp 1698431365
transform 1 0 29680 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1482_
timestamp 1698431365
transform 1 0 31024 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1483_
timestamp 1698431365
transform 1 0 31248 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1698431365
transform 1 0 13888 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1485_
timestamp 1698431365
transform -1 0 16240 0 -1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1486_
timestamp 1698431365
transform -1 0 15568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1487_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1488_
timestamp 1698431365
transform 1 0 8512 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1489_
timestamp 1698431365
transform -1 0 10080 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1490_
timestamp 1698431365
transform -1 0 9072 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1491_
timestamp 1698431365
transform -1 0 10080 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1492_
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1493_
timestamp 1698431365
transform -1 0 15456 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1494_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14672 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1495_
timestamp 1698431365
transform 1 0 15792 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1496_
timestamp 1698431365
transform 1 0 33264 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1497_
timestamp 1698431365
transform 1 0 35056 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1498_
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_
timestamp 1698431365
transform -1 0 42672 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1500_
timestamp 1698431365
transform -1 0 31472 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1501_
timestamp 1698431365
transform -1 0 30576 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1502_
timestamp 1698431365
transform -1 0 30016 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1503_
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1504_
timestamp 1698431365
transform -1 0 31808 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1505_
timestamp 1698431365
transform 1 0 26320 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1506_
timestamp 1698431365
transform -1 0 29568 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1507_
timestamp 1698431365
transform -1 0 29568 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1508_
timestamp 1698431365
transform 1 0 28336 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1509_
timestamp 1698431365
transform 1 0 28224 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1510_
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1511_
timestamp 1698431365
transform 1 0 30352 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1512_
timestamp 1698431365
transform -1 0 20944 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1698431365
transform 1 0 21056 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1514_
timestamp 1698431365
transform -1 0 22176 0 -1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1515_
timestamp 1698431365
transform -1 0 18816 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1516_
timestamp 1698431365
transform -1 0 9968 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1517_
timestamp 1698431365
transform 1 0 7616 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1518_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1519_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1520_
timestamp 1698431365
transform 1 0 10864 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1521_
timestamp 1698431365
transform -1 0 13664 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1522_
timestamp 1698431365
transform -1 0 15120 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1523_
timestamp 1698431365
transform 1 0 14896 0 -1 54880
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1524_
timestamp 1698431365
transform 1 0 32592 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1525_
timestamp 1698431365
transform -1 0 31248 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1698431365
transform -1 0 31808 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1527_
timestamp 1698431365
transform 1 0 31808 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1528_
timestamp 1698431365
transform 1 0 32592 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1529_
timestamp 1698431365
transform 1 0 33376 0 -1 56448
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1530_
timestamp 1698431365
transform 1 0 35280 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1698431365
transform -1 0 36960 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1532_
timestamp 1698431365
transform -1 0 36624 0 1 53312
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1533_
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1534_
timestamp 1698431365
transform 1 0 41888 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1535_
timestamp 1698431365
transform 1 0 34384 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1536_
timestamp 1698431365
transform -1 0 36624 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform -1 0 31248 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1538_
timestamp 1698431365
transform 1 0 29904 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1539_
timestamp 1698431365
transform 1 0 31248 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1540_
timestamp 1698431365
transform -1 0 32592 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1541_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31696 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1542_
timestamp 1698431365
transform 1 0 11312 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1543_
timestamp 1698431365
transform -1 0 12096 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1544_
timestamp 1698431365
transform -1 0 14672 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1545_
timestamp 1698431365
transform 1 0 14896 0 -1 40768
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1546_
timestamp 1698431365
transform 1 0 12656 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1547_
timestamp 1698431365
transform -1 0 11760 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1548_
timestamp 1698431365
transform -1 0 12656 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1549_
timestamp 1698431365
transform 1 0 11872 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1550_
timestamp 1698431365
transform 1 0 13776 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1551_
timestamp 1698431365
transform -1 0 11536 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1552_
timestamp 1698431365
transform -1 0 10864 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1698431365
transform 1 0 10864 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1554_
timestamp 1698431365
transform 1 0 14336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1555_
timestamp 1698431365
transform -1 0 14896 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1556_
timestamp 1698431365
transform 1 0 14784 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1698431365
transform -1 0 23968 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1558_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1559_
timestamp 1698431365
transform -1 0 30800 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1560_
timestamp 1698431365
transform 1 0 30576 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1561_
timestamp 1698431365
transform 1 0 25648 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1562_
timestamp 1698431365
transform 1 0 26992 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1563_
timestamp 1698431365
transform 1 0 25872 0 -1 58016
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1564_
timestamp 1698431365
transform 1 0 35952 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1565_
timestamp 1698431365
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1566_
timestamp 1698431365
transform -1 0 36512 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1567_
timestamp 1698431365
transform 1 0 35392 0 -1 56448
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1568_
timestamp 1698431365
transform -1 0 36176 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1569_
timestamp 1698431365
transform -1 0 25648 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1570_
timestamp 1698431365
transform -1 0 25872 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1571_
timestamp 1698431365
transform 1 0 25200 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1572_
timestamp 1698431365
transform 1 0 26656 0 1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1573_
timestamp 1698431365
transform -1 0 31472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1574_
timestamp 1698431365
transform -1 0 30240 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1575_
timestamp 1698431365
transform -1 0 28112 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1576_
timestamp 1698431365
transform 1 0 27664 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform -1 0 27552 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1698431365
transform 1 0 26992 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1698431365
transform -1 0 29568 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1580_
timestamp 1698431365
transform -1 0 15680 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1698431365
transform -1 0 14000 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1582_
timestamp 1698431365
transform -1 0 13216 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1583_
timestamp 1698431365
transform -1 0 11984 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1584_
timestamp 1698431365
transform -1 0 10528 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1585_
timestamp 1698431365
transform 1 0 9968 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1586_
timestamp 1698431365
transform -1 0 13440 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1587_
timestamp 1698431365
transform 1 0 10976 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1588_
timestamp 1698431365
transform 1 0 12096 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1589_
timestamp 1698431365
transform 1 0 12208 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1590_
timestamp 1698431365
transform 1 0 13216 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1591_
timestamp 1698431365
transform -1 0 15344 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1592_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1593_
timestamp 1698431365
transform 1 0 28448 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1594_
timestamp 1698431365
transform 1 0 35616 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1595_
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1596_
timestamp 1698431365
transform 1 0 42784 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform 1 0 34832 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1598_
timestamp 1698431365
transform 1 0 34272 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1599_
timestamp 1698431365
transform -1 0 37520 0 -1 59584
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1600_
timestamp 1698431365
transform 1 0 27552 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1601_
timestamp 1698431365
transform -1 0 34384 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1602_
timestamp 1698431365
transform -1 0 31472 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1603_
timestamp 1698431365
transform 1 0 30912 0 1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1604_
timestamp 1698431365
transform -1 0 14896 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1605_
timestamp 1698431365
transform 1 0 15456 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1606_
timestamp 1698431365
transform 1 0 16016 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1607_
timestamp 1698431365
transform 1 0 16240 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1608_
timestamp 1698431365
transform -1 0 16240 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1698431365
transform 1 0 17808 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1698431365
transform 1 0 16016 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1611_
timestamp 1698431365
transform 1 0 12208 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1698431365
transform -1 0 14112 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1613_
timestamp 1698431365
transform -1 0 14448 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1614_
timestamp 1698431365
transform -1 0 15344 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1615_
timestamp 1698431365
transform 1 0 16576 0 1 59584
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1616_
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1617_
timestamp 1698431365
transform 1 0 34272 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1618_
timestamp 1698431365
transform 1 0 36736 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1619_
timestamp 1698431365
transform 1 0 47040 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1620_
timestamp 1698431365
transform 1 0 31808 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1621_
timestamp 1698431365
transform -1 0 30912 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1698431365
transform 1 0 32256 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform -1 0 33376 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1698431365
transform -1 0 32928 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1626_
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1627_
timestamp 1698431365
transform 1 0 37408 0 -1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1628_
timestamp 1698431365
transform 1 0 34048 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1629_
timestamp 1698431365
transform -1 0 37744 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1698431365
transform 1 0 38304 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1631_
timestamp 1698431365
transform 1 0 52304 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1632_
timestamp 1698431365
transform 1 0 38080 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1633_
timestamp 1698431365
transform -1 0 40320 0 -1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1634_
timestamp 1698431365
transform 1 0 52864 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1635_
timestamp 1698431365
transform -1 0 53424 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1636_
timestamp 1698431365
transform -1 0 55104 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform 1 0 50624 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1638_
timestamp 1698431365
transform 1 0 51632 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1639_
timestamp 1698431365
transform -1 0 50512 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1640_
timestamp 1698431365
transform 1 0 29792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1641_
timestamp 1698431365
transform -1 0 35168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1642_
timestamp 1698431365
transform -1 0 40320 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1643_
timestamp 1698431365
transform -1 0 29792 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1644_
timestamp 1698431365
transform -1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1645_
timestamp 1698431365
transform 1 0 23408 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1646_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1647_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1648_
timestamp 1698431365
transform -1 0 31584 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1649_
timestamp 1698431365
transform -1 0 32032 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1650_
timestamp 1698431365
transform -1 0 31472 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1698431365
transform -1 0 36064 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1652_
timestamp 1698431365
transform 1 0 35616 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1653_
timestamp 1698431365
transform -1 0 35280 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1654_
timestamp 1698431365
transform 1 0 30240 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1655_
timestamp 1698431365
transform -1 0 57568 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1656_
timestamp 1698431365
transform -1 0 34944 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1657_
timestamp 1698431365
transform 1 0 33600 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1658_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1659_
timestamp 1698431365
transform 1 0 23072 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1660_
timestamp 1698431365
transform -1 0 42672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1661_
timestamp 1698431365
transform 1 0 31360 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1662_
timestamp 1698431365
transform 1 0 30464 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1663_
timestamp 1698431365
transform -1 0 34160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1664_
timestamp 1698431365
transform -1 0 33824 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1665_
timestamp 1698431365
transform -1 0 31136 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1666_
timestamp 1698431365
transform -1 0 31360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1667_
timestamp 1698431365
transform -1 0 58016 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1668_
timestamp 1698431365
transform -1 0 44352 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1669_
timestamp 1698431365
transform 1 0 31136 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1670_
timestamp 1698431365
transform 1 0 30800 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1671_
timestamp 1698431365
transform -1 0 49056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1672_
timestamp 1698431365
transform -1 0 39536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1673_
timestamp 1698431365
transform 1 0 40432 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1675_
timestamp 1698431365
transform 1 0 42672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1676_
timestamp 1698431365
transform 1 0 43344 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1698431365
transform 1 0 46032 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1678_
timestamp 1698431365
transform 1 0 46592 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1679_
timestamp 1698431365
transform 1 0 46032 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1680_
timestamp 1698431365
transform 1 0 45136 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1681_
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1682_
timestamp 1698431365
transform 1 0 45696 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1683_
timestamp 1698431365
transform 1 0 44912 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1684_
timestamp 1698431365
transform 1 0 43456 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1685_
timestamp 1698431365
transform 1 0 42784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1686_
timestamp 1698431365
transform -1 0 49952 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1687_
timestamp 1698431365
transform 1 0 30016 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1688_
timestamp 1698431365
transform 1 0 39536 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform 1 0 44464 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1690_
timestamp 1698431365
transform 1 0 45360 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1691_
timestamp 1698431365
transform -1 0 47600 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1692_
timestamp 1698431365
transform 1 0 46592 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1693_
timestamp 1698431365
transform 1 0 46816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1694_
timestamp 1698431365
transform 1 0 46480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1695_
timestamp 1698431365
transform 1 0 47376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1696_
timestamp 1698431365
transform 1 0 45472 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1697_
timestamp 1698431365
transform -1 0 23296 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1698_
timestamp 1698431365
transform 1 0 20160 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1699_
timestamp 1698431365
transform -1 0 46928 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1700_
timestamp 1698431365
transform 1 0 45584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1701_
timestamp 1698431365
transform 1 0 40992 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1702_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1703_
timestamp 1698431365
transform 1 0 49952 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1704_
timestamp 1698431365
transform -1 0 49504 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1705_
timestamp 1698431365
transform -1 0 42336 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1707_
timestamp 1698431365
transform 1 0 38528 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1708_
timestamp 1698431365
transform 1 0 40768 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1709_
timestamp 1698431365
transform 1 0 38752 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1710_
timestamp 1698431365
transform 1 0 39424 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1711_
timestamp 1698431365
transform -1 0 40544 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1712_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1713_
timestamp 1698431365
transform 1 0 22512 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1714_
timestamp 1698431365
transform 1 0 22064 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1715_
timestamp 1698431365
transform 1 0 49056 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1716_
timestamp 1698431365
transform -1 0 49504 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1717_
timestamp 1698431365
transform -1 0 24528 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform 1 0 21504 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1719_
timestamp 1698431365
transform 1 0 22064 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1720_
timestamp 1698431365
transform 1 0 22960 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1721_
timestamp 1698431365
transform -1 0 24192 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1698431365
transform 1 0 23296 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1723_
timestamp 1698431365
transform -1 0 24864 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1724_
timestamp 1698431365
transform -1 0 25088 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1725_
timestamp 1698431365
transform -1 0 23856 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1726_
timestamp 1698431365
transform 1 0 19488 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1727_
timestamp 1698431365
transform 1 0 19264 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1728_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1729_
timestamp 1698431365
transform 1 0 19936 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1730_
timestamp 1698431365
transform 1 0 19040 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1698431365
transform 1 0 21280 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1732_
timestamp 1698431365
transform -1 0 21280 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1733_
timestamp 1698431365
transform -1 0 19712 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1734_
timestamp 1698431365
transform 1 0 6832 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1735_
timestamp 1698431365
transform 1 0 18480 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1736_
timestamp 1698431365
transform -1 0 18480 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1737_
timestamp 1698431365
transform -1 0 20832 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1738_
timestamp 1698431365
transform -1 0 20272 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1739_
timestamp 1698431365
transform 1 0 20048 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1740_
timestamp 1698431365
transform -1 0 24864 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1741_
timestamp 1698431365
transform -1 0 22848 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1742_
timestamp 1698431365
transform -1 0 23520 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1743_
timestamp 1698431365
transform 1 0 23744 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1744_
timestamp 1698431365
transform 1 0 23520 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1745_
timestamp 1698431365
transform -1 0 24752 0 -1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1746_
timestamp 1698431365
transform 1 0 22512 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1747_
timestamp 1698431365
transform 1 0 23408 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1748_
timestamp 1698431365
transform -1 0 24976 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1749_
timestamp 1698431365
transform -1 0 24864 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1750_
timestamp 1698431365
transform -1 0 25760 0 1 59584
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1751_
timestamp 1698431365
transform -1 0 23184 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1752_
timestamp 1698431365
transform -1 0 22064 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1753_
timestamp 1698431365
transform 1 0 24752 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1754_
timestamp 1698431365
transform 1 0 25760 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1755_
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1756_
timestamp 1698431365
transform 1 0 25760 0 1 59584
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1757_
timestamp 1698431365
transform -1 0 21168 0 -1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1758_
timestamp 1698431365
transform -1 0 18368 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1759_
timestamp 1698431365
transform -1 0 19936 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1760_
timestamp 1698431365
transform -1 0 20496 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1761_
timestamp 1698431365
transform -1 0 20832 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1698431365
transform -1 0 11760 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1763_
timestamp 1698431365
transform 1 0 3472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1764_
timestamp 1698431365
transform 1 0 2576 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform -1 0 4256 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1766_
timestamp 1698431365
transform -1 0 4928 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1767_
timestamp 1698431365
transform -1 0 3248 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1768_
timestamp 1698431365
transform -1 0 6160 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1698431365
transform -1 0 6048 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1770_
timestamp 1698431365
transform -1 0 5264 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1771_
timestamp 1698431365
transform -1 0 6384 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1698431365
transform -1 0 5264 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1773_
timestamp 1698431365
transform -1 0 3808 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1774_
timestamp 1698431365
transform -1 0 4144 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1775_
timestamp 1698431365
transform -1 0 3024 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1776_
timestamp 1698431365
transform -1 0 5264 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1777_
timestamp 1698431365
transform -1 0 5264 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1778_
timestamp 1698431365
transform -1 0 5936 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1779_
timestamp 1698431365
transform -1 0 2912 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1698431365
transform -1 0 6160 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1698431365
transform -1 0 6496 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1782_
timestamp 1698431365
transform -1 0 5936 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1783_
timestamp 1698431365
transform 1 0 4816 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1698431365
transform 1 0 2912 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1785_
timestamp 1698431365
transform -1 0 4592 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1786_
timestamp 1698431365
transform 1 0 4256 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1698431365
transform 1 0 3136 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1788_
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1789_
timestamp 1698431365
transform -1 0 6272 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1790_
timestamp 1698431365
transform -1 0 4144 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1791_
timestamp 1698431365
transform -1 0 7504 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1792_
timestamp 1698431365
transform 1 0 3696 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1793_
timestamp 1698431365
transform 1 0 2800 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1794_
timestamp 1698431365
transform 1 0 4144 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1795_
timestamp 1698431365
transform 1 0 4816 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1796_
timestamp 1698431365
transform -1 0 5152 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1797_
timestamp 1698431365
transform -1 0 6160 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1798_
timestamp 1698431365
transform 1 0 4256 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1698431365
transform 1 0 3696 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1800_
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1801_
timestamp 1698431365
transform -1 0 20944 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1803_
timestamp 1698431365
transform -1 0 6384 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1804_
timestamp 1698431365
transform 1 0 6160 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1805_
timestamp 1698431365
transform 1 0 5824 0 -1 61152
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1806_
timestamp 1698431365
transform -1 0 7952 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1807_
timestamp 1698431365
transform -1 0 6608 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform 1 0 6608 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1809_
timestamp 1698431365
transform -1 0 7952 0 1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1810_
timestamp 1698431365
transform -1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1811_
timestamp 1698431365
transform -1 0 8848 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1812_
timestamp 1698431365
transform -1 0 7504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1813_
timestamp 1698431365
transform 1 0 6384 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1814_
timestamp 1698431365
transform 1 0 7728 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1815_
timestamp 1698431365
transform 1 0 8288 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1816_
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1817_
timestamp 1698431365
transform -1 0 20944 0 1 59584
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1818_
timestamp 1698431365
transform 1 0 19824 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1819_
timestamp 1698431365
transform -1 0 19712 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1820_
timestamp 1698431365
transform 1 0 35504 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1821_
timestamp 1698431365
transform -1 0 42896 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1822_
timestamp 1698431365
transform 1 0 19712 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1823_
timestamp 1698431365
transform -1 0 20160 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1824_
timestamp 1698431365
transform -1 0 12992 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1825_
timestamp 1698431365
transform -1 0 6832 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1826_
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1827_
timestamp 1698431365
transform 1 0 7728 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1828_
timestamp 1698431365
transform -1 0 10416 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1829_
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1830_
timestamp 1698431365
transform 1 0 8624 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1831_
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1832_
timestamp 1698431365
transform -1 0 11088 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1833_
timestamp 1698431365
transform -1 0 9296 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1834_
timestamp 1698431365
transform 1 0 7616 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1835_
timestamp 1698431365
transform 1 0 7952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1698431365
transform 1 0 7056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1698431365
transform 1 0 8624 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1838_
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1839_
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1840_
timestamp 1698431365
transform 1 0 10080 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1841_
timestamp 1698431365
transform 1 0 12432 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1842_
timestamp 1698431365
transform 1 0 10976 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 13888 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1844_
timestamp 1698431365
transform -1 0 12320 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1845_
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1846_
timestamp 1698431365
transform -1 0 9184 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1847_
timestamp 1698431365
transform -1 0 8736 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1848_
timestamp 1698431365
transform 1 0 9072 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1849_
timestamp 1698431365
transform -1 0 10528 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1850_
timestamp 1698431365
transform -1 0 9968 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1851_
timestamp 1698431365
transform -1 0 10416 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1852_
timestamp 1698431365
transform -1 0 8512 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1698431365
transform 1 0 8288 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 6944 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1855_
timestamp 1698431365
transform 1 0 8512 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1856_
timestamp 1698431365
transform -1 0 8736 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1857_
timestamp 1698431365
transform 1 0 8736 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1858_
timestamp 1698431365
transform -1 0 11088 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1859_
timestamp 1698431365
transform -1 0 8960 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1860_
timestamp 1698431365
transform 1 0 7840 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1861_
timestamp 1698431365
transform -1 0 48384 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1862_
timestamp 1698431365
transform -1 0 10864 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1863_
timestamp 1698431365
transform -1 0 10304 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1864_
timestamp 1698431365
transform 1 0 10080 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1865_
timestamp 1698431365
transform 1 0 9968 0 1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1866_
timestamp 1698431365
transform -1 0 12208 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1867_
timestamp 1698431365
transform 1 0 10640 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1868_
timestamp 1698431365
transform -1 0 13552 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1869_
timestamp 1698431365
transform -1 0 12992 0 -1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1870_
timestamp 1698431365
transform 1 0 10752 0 -1 64288
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform -1 0 12880 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1872_
timestamp 1698431365
transform 1 0 11760 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1873_
timestamp 1698431365
transform 1 0 12544 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1874_
timestamp 1698431365
transform -1 0 14000 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1875_
timestamp 1698431365
transform -1 0 14224 0 -1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1876_
timestamp 1698431365
transform -1 0 17248 0 1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1877_
timestamp 1698431365
transform 1 0 14672 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1698431365
transform 1 0 16240 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1879_
timestamp 1698431365
transform 1 0 25312 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1880_
timestamp 1698431365
transform -1 0 39424 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1881_
timestamp 1698431365
transform 1 0 17248 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1882_
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1883_
timestamp 1698431365
transform -1 0 57344 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1884_
timestamp 1698431365
transform 1 0 48720 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1885_
timestamp 1698431365
transform 1 0 53760 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1886_
timestamp 1698431365
transform -1 0 55440 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1887_
timestamp 1698431365
transform -1 0 53872 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1888_
timestamp 1698431365
transform 1 0 50400 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1889_
timestamp 1698431365
transform -1 0 56224 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1890_
timestamp 1698431365
transform -1 0 57120 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1891_
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1892_
timestamp 1698431365
transform -1 0 54768 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1893_
timestamp 1698431365
transform -1 0 55664 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1894_
timestamp 1698431365
transform 1 0 53312 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1895_
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1896_
timestamp 1698431365
transform -1 0 52304 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1698431365
transform -1 0 51408 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1898_
timestamp 1698431365
transform 1 0 51408 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1899_
timestamp 1698431365
transform 1 0 35392 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1900_
timestamp 1698431365
transform 1 0 49056 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1901_
timestamp 1698431365
transform 1 0 51408 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1698431365
transform -1 0 50400 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1903_
timestamp 1698431365
transform 1 0 50176 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1904_
timestamp 1698431365
transform -1 0 52192 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1698431365
transform -1 0 51520 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1906_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1907_
timestamp 1698431365
transform 1 0 49280 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1908_
timestamp 1698431365
transform 1 0 52752 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1909_
timestamp 1698431365
transform -1 0 53424 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1910_
timestamp 1698431365
transform -1 0 50960 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1911_
timestamp 1698431365
transform -1 0 50400 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1912_
timestamp 1698431365
transform 1 0 49392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1913_
timestamp 1698431365
transform 1 0 51296 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1914_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49168 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1915_
timestamp 1698431365
transform 1 0 50064 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1916_
timestamp 1698431365
transform 1 0 51632 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1917_
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1918_
timestamp 1698431365
transform -1 0 53760 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1919_
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1920_
timestamp 1698431365
transform 1 0 50848 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1921_
timestamp 1698431365
transform 1 0 52976 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1922_
timestamp 1698431365
transform -1 0 53984 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1698431365
transform -1 0 52864 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1924_
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1925_
timestamp 1698431365
transform -1 0 53984 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform -1 0 53088 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1927_
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1928_
timestamp 1698431365
transform -1 0 53984 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1698431365
transform 1 0 53984 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1930_
timestamp 1698431365
transform -1 0 53424 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1931_
timestamp 1698431365
transform 1 0 53872 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1932_
timestamp 1698431365
transform 1 0 54992 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1933_
timestamp 1698431365
transform -1 0 57568 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1934_
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1935_
timestamp 1698431365
transform 1 0 54432 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1936_
timestamp 1698431365
transform 1 0 54432 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1937_
timestamp 1698431365
transform -1 0 58128 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698431365
transform -1 0 57008 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1939_
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1698431365
transform -1 0 56896 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1942_
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1698431365
transform 1 0 57680 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1698431365
transform 1 0 57120 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1698431365
transform -1 0 57344 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1698431365
transform -1 0 57232 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1947_
timestamp 1698431365
transform 1 0 54656 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1948_
timestamp 1698431365
transform 1 0 57344 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1949_
timestamp 1698431365
transform 1 0 54880 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1950_
timestamp 1698431365
transform -1 0 57344 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1951_
timestamp 1698431365
transform 1 0 52976 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform -1 0 57344 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1953_
timestamp 1698431365
transform -1 0 57232 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1954_
timestamp 1698431365
transform 1 0 56560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1698431365
transform 1 0 57456 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1698431365
transform 1 0 56112 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform 1 0 56560 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1958_
timestamp 1698431365
transform -1 0 56000 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform -1 0 55216 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1960_
timestamp 1698431365
transform 1 0 54880 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1698431365
transform -1 0 54208 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1962_
timestamp 1698431365
transform -1 0 52304 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1963_
timestamp 1698431365
transform -1 0 52304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1964_
timestamp 1698431365
transform -1 0 46816 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1965_
timestamp 1698431365
transform 1 0 46256 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1966_
timestamp 1698431365
transform 1 0 50176 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1967_
timestamp 1698431365
transform 1 0 48832 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1968_
timestamp 1698431365
transform -1 0 57568 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1969_
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1970_
timestamp 1698431365
transform -1 0 58016 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1698431365
transform -1 0 56224 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1972_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 54208 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1973_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 54768 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1974_
timestamp 1698431365
transform 1 0 42896 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1975_
timestamp 1698431365
transform 1 0 45472 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1698431365
transform 1 0 47152 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1977_
timestamp 1698431365
transform 1 0 49504 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1978_
timestamp 1698431365
transform -1 0 57792 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1979_
timestamp 1698431365
transform -1 0 57904 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1980_
timestamp 1698431365
transform -1 0 42224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1981_
timestamp 1698431365
transform 1 0 26656 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1982_
timestamp 1698431365
transform 1 0 38528 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1983_
timestamp 1698431365
transform 1 0 42784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1984_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1985_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1986_
timestamp 1698431365
transform -1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1987_
timestamp 1698431365
transform -1 0 44352 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1988_
timestamp 1698431365
transform -1 0 44240 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1989_
timestamp 1698431365
transform -1 0 43792 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1990_
timestamp 1698431365
transform -1 0 43344 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1991_
timestamp 1698431365
transform -1 0 44464 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1992_
timestamp 1698431365
transform -1 0 44240 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1993_
timestamp 1698431365
transform 1 0 43792 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1698431365
transform 1 0 43792 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1995_
timestamp 1698431365
transform -1 0 43792 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1996_
timestamp 1698431365
transform 1 0 41888 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1997_
timestamp 1698431365
transform -1 0 41888 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1998_
timestamp 1698431365
transform -1 0 42448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform -1 0 44352 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2000_
timestamp 1698431365
transform 1 0 43904 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2001_
timestamp 1698431365
transform -1 0 45248 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1698431365
transform -1 0 44240 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2003_
timestamp 1698431365
transform 1 0 45472 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2004_
timestamp 1698431365
transform 1 0 46816 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2005_
timestamp 1698431365
transform 1 0 45808 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2006_
timestamp 1698431365
transform -1 0 46256 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2007_
timestamp 1698431365
transform 1 0 46256 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2008_
timestamp 1698431365
transform -1 0 47712 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2009_
timestamp 1698431365
transform 1 0 43120 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2010_
timestamp 1698431365
transform 1 0 44912 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2011_
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2012_
timestamp 1698431365
transform -1 0 44464 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2013_
timestamp 1698431365
transform 1 0 45024 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2014_
timestamp 1698431365
transform -1 0 45024 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2015_
timestamp 1698431365
transform 1 0 31920 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2016_
timestamp 1698431365
transform 1 0 34496 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2017_
timestamp 1698431365
transform 1 0 33600 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2018_
timestamp 1698431365
transform -1 0 38304 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2019_
timestamp 1698431365
transform 1 0 31024 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2020_
timestamp 1698431365
transform 1 0 31696 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2021_
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2022_
timestamp 1698431365
transform 1 0 29008 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2023_
timestamp 1698431365
transform 1 0 31584 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2024_
timestamp 1698431365
transform 1 0 29232 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2025_
timestamp 1698431365
transform 1 0 28448 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2026_
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2027_
timestamp 1698431365
transform 1 0 28336 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2028_
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2029_
timestamp 1698431365
transform -1 0 29680 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2030_
timestamp 1698431365
transform 1 0 30352 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2031_
timestamp 1698431365
transform 1 0 28224 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2032_
timestamp 1698431365
transform 1 0 29680 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2033_
timestamp 1698431365
transform -1 0 30464 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2034_
timestamp 1698431365
transform -1 0 28784 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2035_
timestamp 1698431365
transform 1 0 27664 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2036_
timestamp 1698431365
transform 1 0 27552 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2037_
timestamp 1698431365
transform 1 0 26544 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2038_
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2039_
timestamp 1698431365
transform 1 0 28784 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2040_
timestamp 1698431365
transform -1 0 30576 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2041_
timestamp 1698431365
transform 1 0 29232 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2042_
timestamp 1698431365
transform 1 0 31920 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2043_
timestamp 1698431365
transform 1 0 29680 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2044_
timestamp 1698431365
transform 1 0 30352 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2045_
timestamp 1698431365
transform -1 0 31024 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2046_
timestamp 1698431365
transform 1 0 25984 0 -1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1698431365
transform 1 0 26880 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2048_
timestamp 1698431365
transform 1 0 25984 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2049_
timestamp 1698431365
transform -1 0 28336 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2050_
timestamp 1698431365
transform 1 0 27104 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2051_
timestamp 1698431365
transform 1 0 27328 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2052_
timestamp 1698431365
transform -1 0 30688 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2053_
timestamp 1698431365
transform -1 0 29904 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2054_
timestamp 1698431365
transform 1 0 28784 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2055_
timestamp 1698431365
transform 1 0 31024 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2056_
timestamp 1698431365
transform -1 0 31248 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2057_
timestamp 1698431365
transform 1 0 32816 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2058_
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2059_
timestamp 1698431365
transform -1 0 35280 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2060_
timestamp 1698431365
transform -1 0 32816 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2061_
timestamp 1698431365
transform -1 0 32592 0 1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2062_
timestamp 1698431365
transform -1 0 32704 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2063_
timestamp 1698431365
transform -1 0 23856 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2064_
timestamp 1698431365
transform 1 0 49616 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2065_
timestamp 1698431365
transform -1 0 52416 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2066_
timestamp 1698431365
transform 1 0 41552 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2067_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 54208 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2068_
timestamp 1698431365
transform 1 0 46480 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2069_
timestamp 1698431365
transform -1 0 51856 0 1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2070_
timestamp 1698431365
transform -1 0 51744 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2071_
timestamp 1698431365
transform 1 0 50848 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2072_
timestamp 1698431365
transform 1 0 51408 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2073_
timestamp 1698431365
transform -1 0 28448 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2074_
timestamp 1698431365
transform 1 0 51184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2075_
timestamp 1698431365
transform 1 0 50288 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2076_
timestamp 1698431365
transform 1 0 51184 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2077_
timestamp 1698431365
transform -1 0 37744 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2078_
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2079_
timestamp 1698431365
transform 1 0 51296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2080_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 52080 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2081_
timestamp 1698431365
transform 1 0 54320 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2082_
timestamp 1698431365
transform 1 0 50400 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2083_
timestamp 1698431365
transform 1 0 53424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1698431365
transform -1 0 52304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2085_
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2086_
timestamp 1698431365
transform 1 0 54992 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2087_
timestamp 1698431365
transform -1 0 49504 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2088_
timestamp 1698431365
transform 1 0 49952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2089_
timestamp 1698431365
transform -1 0 51968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2090_
timestamp 1698431365
transform -1 0 52864 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2091_
timestamp 1698431365
transform 1 0 43568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2092_
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2093_
timestamp 1698431365
transform 1 0 53872 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2094_
timestamp 1698431365
transform -1 0 49616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2095_
timestamp 1698431365
transform -1 0 50960 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2096_
timestamp 1698431365
transform 1 0 46704 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2097_
timestamp 1698431365
transform -1 0 51072 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2098_
timestamp 1698431365
transform 1 0 50960 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2099_
timestamp 1698431365
transform 1 0 52528 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2100_
timestamp 1698431365
transform 1 0 49728 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2101_
timestamp 1698431365
transform -1 0 47376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2102_
timestamp 1698431365
transform -1 0 48272 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2103_
timestamp 1698431365
transform -1 0 48048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2104_
timestamp 1698431365
transform -1 0 48384 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2105_
timestamp 1698431365
transform 1 0 47600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2106_
timestamp 1698431365
transform -1 0 45920 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2107_
timestamp 1698431365
transform 1 0 44912 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2108_
timestamp 1698431365
transform -1 0 45360 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2109_
timestamp 1698431365
transform -1 0 45248 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2110_
timestamp 1698431365
transform 1 0 43904 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2111_
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2112_
timestamp 1698431365
transform -1 0 44912 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2113_
timestamp 1698431365
transform -1 0 43008 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2114_
timestamp 1698431365
transform -1 0 42560 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2115_
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2116_
timestamp 1698431365
transform 1 0 40880 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2117_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2118_
timestamp 1698431365
transform 1 0 42448 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2119_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41328 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2120_
timestamp 1698431365
transform -1 0 40320 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2121_
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2122_
timestamp 1698431365
transform 1 0 50512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2123_
timestamp 1698431365
transform -1 0 39760 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2124_
timestamp 1698431365
transform 1 0 38640 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2125_
timestamp 1698431365
transform 1 0 39536 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2126_
timestamp 1698431365
transform -1 0 38864 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2127_
timestamp 1698431365
transform 1 0 38080 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2128_
timestamp 1698431365
transform -1 0 39424 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2129_
timestamp 1698431365
transform -1 0 37632 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2130_
timestamp 1698431365
transform 1 0 28560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2131_
timestamp 1698431365
transform 1 0 27664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform 1 0 51184 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2133_
timestamp 1698431365
transform 1 0 48048 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2134_
timestamp 1698431365
transform 1 0 35280 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2135_
timestamp 1698431365
transform -1 0 41664 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2136_
timestamp 1698431365
transform -1 0 50848 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2137_
timestamp 1698431365
transform 1 0 50624 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2138_
timestamp 1698431365
transform 1 0 51408 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2139_
timestamp 1698431365
transform 1 0 47152 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2140_
timestamp 1698431365
transform 1 0 50848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2141_
timestamp 1698431365
transform -1 0 50624 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2142_
timestamp 1698431365
transform 1 0 42784 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2143_
timestamp 1698431365
transform 1 0 50400 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2144_
timestamp 1698431365
transform 1 0 52304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2145_
timestamp 1698431365
transform -1 0 49056 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2146_
timestamp 1698431365
transform -1 0 50176 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2147_
timestamp 1698431365
transform 1 0 49504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2148_
timestamp 1698431365
transform 1 0 50176 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2149_
timestamp 1698431365
transform 1 0 51072 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2150_
timestamp 1698431365
transform -1 0 39872 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2151_
timestamp 1698431365
transform -1 0 39760 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2152_
timestamp 1698431365
transform 1 0 39648 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2153_
timestamp 1698431365
transform -1 0 42000 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2154_
timestamp 1698431365
transform -1 0 40432 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2155_
timestamp 1698431365
transform -1 0 41664 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2156_
timestamp 1698431365
transform -1 0 41104 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2157_
timestamp 1698431365
transform 1 0 40544 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2158_
timestamp 1698431365
transform -1 0 37856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2159_
timestamp 1698431365
transform -1 0 38304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2160_
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2161_
timestamp 1698431365
transform -1 0 39088 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2162_
timestamp 1698431365
transform 1 0 37968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2163_
timestamp 1698431365
transform -1 0 35728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2164_
timestamp 1698431365
transform -1 0 35728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2165_
timestamp 1698431365
transform 1 0 35728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2166_
timestamp 1698431365
transform -1 0 36960 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2167_
timestamp 1698431365
transform -1 0 36288 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2168_
timestamp 1698431365
transform 1 0 35280 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2169_
timestamp 1698431365
transform -1 0 34608 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2170_
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2171_
timestamp 1698431365
transform 1 0 33488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2172_
timestamp 1698431365
transform 1 0 33376 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2173_
timestamp 1698431365
transform -1 0 33040 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2174_
timestamp 1698431365
transform 1 0 33376 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2175_
timestamp 1698431365
transform -1 0 34048 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2176_
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2177_
timestamp 1698431365
transform 1 0 31360 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2178_
timestamp 1698431365
transform 1 0 32592 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2179_
timestamp 1698431365
transform -1 0 33600 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2180_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2181_
timestamp 1698431365
transform -1 0 32704 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2182_
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2183_
timestamp 1698431365
transform 1 0 34720 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2184_
timestamp 1698431365
transform 1 0 34272 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2185_
timestamp 1698431365
transform 1 0 34160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2186_
timestamp 1698431365
transform 1 0 35168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2187_
timestamp 1698431365
transform -1 0 42448 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2188_
timestamp 1698431365
transform -1 0 32816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2189_
timestamp 1698431365
transform 1 0 33600 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2190_
timestamp 1698431365
transform 1 0 34160 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2191_
timestamp 1698431365
transform 1 0 35168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2192_
timestamp 1698431365
transform 1 0 39424 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2194_
timestamp 1698431365
transform 1 0 7504 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2195_
timestamp 1698431365
transform -1 0 27664 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2196_
timestamp 1698431365
transform 1 0 23520 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2197_
timestamp 1698431365
transform 1 0 18592 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2198_
timestamp 1698431365
transform 1 0 23184 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2199_
timestamp 1698431365
transform 1 0 27328 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2200_
timestamp 1698431365
transform -1 0 26544 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2201_
timestamp 1698431365
transform 1 0 26544 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2202_
timestamp 1698431365
transform -1 0 27776 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2203_
timestamp 1698431365
transform 1 0 26544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2204_
timestamp 1698431365
transform -1 0 26544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2205_
timestamp 1698431365
transform 1 0 26544 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2206_
timestamp 1698431365
transform -1 0 27104 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2207_
timestamp 1698431365
transform 1 0 25760 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2208_
timestamp 1698431365
transform -1 0 25536 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2209_
timestamp 1698431365
transform -1 0 23520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2210_
timestamp 1698431365
transform -1 0 24528 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2211_
timestamp 1698431365
transform 1 0 23408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2212_
timestamp 1698431365
transform 1 0 23296 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2213_
timestamp 1698431365
transform -1 0 23408 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2214_
timestamp 1698431365
transform -1 0 22624 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2215_
timestamp 1698431365
transform 1 0 21392 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2216_
timestamp 1698431365
transform -1 0 21504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2217_
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1698431365
transform -1 0 21952 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2219_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2220_
timestamp 1698431365
transform -1 0 20384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2221_
timestamp 1698431365
transform -1 0 19488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2222_
timestamp 1698431365
transform -1 0 19488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2223_
timestamp 1698431365
transform 1 0 19488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2224_
timestamp 1698431365
transform -1 0 19824 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2225_
timestamp 1698431365
transform -1 0 17696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2226_
timestamp 1698431365
transform -1 0 18592 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2227_
timestamp 1698431365
transform -1 0 18480 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2228_
timestamp 1698431365
transform 1 0 18592 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2229_
timestamp 1698431365
transform -1 0 19824 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2230_
timestamp 1698431365
transform -1 0 16016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2231_
timestamp 1698431365
transform -1 0 21840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2232_
timestamp 1698431365
transform -1 0 19040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2233_
timestamp 1698431365
transform 1 0 19040 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2234_
timestamp 1698431365
transform -1 0 18144 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2235_
timestamp 1698431365
transform 1 0 19712 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2236_
timestamp 1698431365
transform -1 0 19824 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2237_
timestamp 1698431365
transform -1 0 16016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2238_
timestamp 1698431365
transform 1 0 20272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2239_
timestamp 1698431365
transform 1 0 18144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2240_
timestamp 1698431365
transform -1 0 20720 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2242_
timestamp 1698431365
transform -1 0 19152 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2243_
timestamp 1698431365
transform -1 0 21952 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2244_
timestamp 1698431365
transform 1 0 22400 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2245_
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2246_
timestamp 1698431365
transform 1 0 23184 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2247_
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2248_
timestamp 1698431365
transform 1 0 24080 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2249_
timestamp 1698431365
transform -1 0 22624 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2250_
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2251_
timestamp 1698431365
transform 1 0 22960 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2252_
timestamp 1698431365
transform 1 0 24304 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2253_
timestamp 1698431365
transform 1 0 19824 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2254_
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2255_
timestamp 1698431365
transform 1 0 36288 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2256_
timestamp 1698431365
transform -1 0 47040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2257_
timestamp 1698431365
transform 1 0 46368 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2258_
timestamp 1698431365
transform -1 0 45920 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34384 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2260_
timestamp 1698431365
transform -1 0 36064 0 -1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2261_
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2262_
timestamp 1698431365
transform -1 0 44464 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2263_
timestamp 1698431365
transform -1 0 41888 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2264_
timestamp 1698431365
transform 1 0 43344 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2265_
timestamp 1698431365
transform 1 0 43792 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2266_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2267_
timestamp 1698431365
transform 1 0 36848 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2268_
timestamp 1698431365
transform 1 0 44240 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2269_
timestamp 1698431365
transform 1 0 45584 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2270_
timestamp 1698431365
transform -1 0 45696 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2271_
timestamp 1698431365
transform -1 0 43344 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2272_
timestamp 1698431365
transform 1 0 43120 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1698431365
transform 1 0 42224 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2274_
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2275_
timestamp 1698431365
transform -1 0 43456 0 1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2276_
timestamp 1698431365
transform -1 0 41440 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2277_
timestamp 1698431365
transform 1 0 41440 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2278_
timestamp 1698431365
transform -1 0 42336 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2279_
timestamp 1698431365
transform 1 0 36960 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2280_
timestamp 1698431365
transform 1 0 41664 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2281_
timestamp 1698431365
transform -1 0 42560 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2282_
timestamp 1698431365
transform -1 0 41664 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1698431365
transform 1 0 41440 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2284_
timestamp 1698431365
transform -1 0 41440 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2285_
timestamp 1698431365
transform 1 0 40768 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2286_
timestamp 1698431365
transform -1 0 41888 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2287_
timestamp 1698431365
transform -1 0 42000 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2288_
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2289_
timestamp 1698431365
transform 1 0 39760 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2290_
timestamp 1698431365
transform 1 0 39312 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2291_
timestamp 1698431365
transform -1 0 49504 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2292_
timestamp 1698431365
transform 1 0 42224 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2293_
timestamp 1698431365
transform 1 0 42672 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2294_
timestamp 1698431365
transform 1 0 41216 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2295_
timestamp 1698431365
transform 1 0 43120 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2296_
timestamp 1698431365
transform 1 0 42784 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2297_
timestamp 1698431365
transform 1 0 44800 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2298_
timestamp 1698431365
transform -1 0 43456 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2299_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43120 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2300_
timestamp 1698431365
transform 1 0 42784 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2301_
timestamp 1698431365
transform 1 0 41216 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2302_
timestamp 1698431365
transform 1 0 39200 0 -1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2303_
timestamp 1698431365
transform -1 0 41104 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2304_
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1698431365
transform -1 0 43008 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2306_
timestamp 1698431365
transform -1 0 42784 0 -1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2307_
timestamp 1698431365
transform -1 0 43904 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2308_
timestamp 1698431365
transform 1 0 40208 0 1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2309_
timestamp 1698431365
transform 1 0 42112 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2310_
timestamp 1698431365
transform 1 0 42896 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2311_
timestamp 1698431365
transform -1 0 47040 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1698431365
transform 1 0 43904 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2313_
timestamp 1698431365
transform -1 0 44352 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2314_
timestamp 1698431365
transform 1 0 44464 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2315_
timestamp 1698431365
transform -1 0 45920 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2316_
timestamp 1698431365
transform 1 0 45920 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2317_
timestamp 1698431365
transform -1 0 45696 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2318_
timestamp 1698431365
transform -1 0 47488 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2319_
timestamp 1698431365
transform 1 0 46368 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2320_
timestamp 1698431365
transform 1 0 52528 0 1 61152
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2321_
timestamp 1698431365
transform 1 0 56448 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2322_
timestamp 1698431365
transform 1 0 53760 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2323_
timestamp 1698431365
transform 1 0 52864 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2324_
timestamp 1698431365
transform -1 0 54992 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2325_
timestamp 1698431365
transform 1 0 53648 0 -1 61152
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2326_
timestamp 1698431365
transform -1 0 57120 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2327_
timestamp 1698431365
transform -1 0 57680 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2328_
timestamp 1698431365
transform 1 0 57568 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2329_
timestamp 1698431365
transform -1 0 57568 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2330_
timestamp 1698431365
transform 1 0 52304 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2331_
timestamp 1698431365
transform -1 0 53200 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2332_
timestamp 1698431365
transform 1 0 51408 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2333_
timestamp 1698431365
transform 1 0 53984 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2334_
timestamp 1698431365
transform -1 0 55104 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2335_
timestamp 1698431365
transform -1 0 56224 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2336_
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2337_
timestamp 1698431365
transform 1 0 54992 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2338_
timestamp 1698431365
transform -1 0 56560 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2339_
timestamp 1698431365
transform 1 0 54544 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2340_
timestamp 1698431365
transform -1 0 55776 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2341_
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2342_
timestamp 1698431365
transform -1 0 56224 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2343_
timestamp 1698431365
transform -1 0 51296 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2344_
timestamp 1698431365
transform 1 0 50736 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2345_
timestamp 1698431365
transform -1 0 52752 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2346_
timestamp 1698431365
transform -1 0 55328 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2347_
timestamp 1698431365
transform -1 0 54768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2348_
timestamp 1698431365
transform -1 0 53424 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2349_
timestamp 1698431365
transform -1 0 49728 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2350_
timestamp 1698431365
transform 1 0 46592 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2351_
timestamp 1698431365
transform 1 0 47152 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2352_
timestamp 1698431365
transform 1 0 39088 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2353_
timestamp 1698431365
transform -1 0 47488 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2354_
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2355_
timestamp 1698431365
transform 1 0 51184 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2356_
timestamp 1698431365
transform 1 0 50736 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46816 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2358_
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2359_
timestamp 1698431365
transform -1 0 47264 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2360_
timestamp 1698431365
transform 1 0 43008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2361_
timestamp 1698431365
transform -1 0 50512 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2362_
timestamp 1698431365
transform 1 0 45696 0 -1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2363_
timestamp 1698431365
transform 1 0 45360 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2364_
timestamp 1698431365
transform 1 0 46704 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2365_
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2366_
timestamp 1698431365
transform -1 0 51520 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2367_
timestamp 1698431365
transform -1 0 50736 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2368_
timestamp 1698431365
transform 1 0 48608 0 -1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2369_
timestamp 1698431365
transform -1 0 48384 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2370_
timestamp 1698431365
transform 1 0 48720 0 -1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2371_
timestamp 1698431365
transform 1 0 48944 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2372_
timestamp 1698431365
transform 1 0 49280 0 -1 64288
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2373_
timestamp 1698431365
transform -1 0 50512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2374_
timestamp 1698431365
transform 1 0 50400 0 1 62720
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2375_
timestamp 1698431365
transform 1 0 51520 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2376_
timestamp 1698431365
transform 1 0 50736 0 1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2377_
timestamp 1698431365
transform 1 0 51856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2378_
timestamp 1698431365
transform -1 0 53536 0 1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2379_
timestamp 1698431365
transform 1 0 51296 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2380_
timestamp 1698431365
transform 1 0 50176 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2381_
timestamp 1698431365
transform -1 0 31808 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2382_
timestamp 1698431365
transform 1 0 31248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2383_
timestamp 1698431365
transform -1 0 24640 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2384_
timestamp 1698431365
transform -1 0 23744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2385_
timestamp 1698431365
transform 1 0 22512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2386_
timestamp 1698431365
transform -1 0 27552 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2387_
timestamp 1698431365
transform 1 0 24640 0 1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2388_
timestamp 1698431365
transform 1 0 36624 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2389_
timestamp 1698431365
transform 1 0 33488 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2390_
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2391_
timestamp 1698431365
transform 1 0 41104 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2392_
timestamp 1698431365
transform -1 0 24528 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2393_
timestamp 1698431365
transform 1 0 34496 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2394_
timestamp 1698431365
transform -1 0 42448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2395_
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2396_
timestamp 1698431365
transform -1 0 36624 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2397_
timestamp 1698431365
transform 1 0 41104 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2398_
timestamp 1698431365
transform 1 0 42000 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2399_
timestamp 1698431365
transform 1 0 39424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2400_
timestamp 1698431365
transform 1 0 38640 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2401_
timestamp 1698431365
transform -1 0 39424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2402_
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2403_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2404_
timestamp 1698431365
transform -1 0 34384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2405_
timestamp 1698431365
transform -1 0 34048 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2406_
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2407_
timestamp 1698431365
transform -1 0 35952 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2408_
timestamp 1698431365
transform 1 0 34160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2409_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2410_
timestamp 1698431365
transform -1 0 27888 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2411_
timestamp 1698431365
transform -1 0 27104 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2412_
timestamp 1698431365
transform 1 0 26320 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2413_
timestamp 1698431365
transform 1 0 27776 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2414_
timestamp 1698431365
transform 1 0 29120 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2415_
timestamp 1698431365
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2416_
timestamp 1698431365
transform 1 0 34832 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2417_
timestamp 1698431365
transform 1 0 28560 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2418_
timestamp 1698431365
transform 1 0 27664 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2419_
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2420_
timestamp 1698431365
transform 1 0 26992 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2421_
timestamp 1698431365
transform 1 0 29792 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2422_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2423_
timestamp 1698431365
transform 1 0 18704 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2424_
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2425_
timestamp 1698431365
transform 1 0 28336 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2426_
timestamp 1698431365
transform 1 0 26432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2427_
timestamp 1698431365
transform 1 0 31360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2428_
timestamp 1698431365
transform 1 0 30464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2429_
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2430_
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2431_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2432_
timestamp 1698431365
transform -1 0 18816 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2433_
timestamp 1698431365
transform -1 0 19488 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2434_
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2435_
timestamp 1698431365
transform 1 0 18368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2436_
timestamp 1698431365
transform -1 0 23296 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2437_
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2438_
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2439_
timestamp 1698431365
transform -1 0 20160 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2440_
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2441_
timestamp 1698431365
transform 1 0 18256 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2442_
timestamp 1698431365
transform 1 0 18144 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2443_
timestamp 1698431365
transform 1 0 17808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1698431365
transform 1 0 21616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2445_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2446_
timestamp 1698431365
transform -1 0 35952 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2447_
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2448_
timestamp 1698431365
transform 1 0 20048 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2449_
timestamp 1698431365
transform -1 0 31472 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2450_
timestamp 1698431365
transform 1 0 24416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2451_
timestamp 1698431365
transform -1 0 32928 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2452_
timestamp 1698431365
transform -1 0 28784 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2453_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2454_
timestamp 1698431365
transform 1 0 25760 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2455_
timestamp 1698431365
transform 1 0 26320 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2456_
timestamp 1698431365
transform 1 0 28560 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2457_
timestamp 1698431365
transform 1 0 27888 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2458_
timestamp 1698431365
transform 1 0 30464 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2459_
timestamp 1698431365
transform 1 0 30688 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2461_
timestamp 1698431365
transform -1 0 25760 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2462_
timestamp 1698431365
transform 1 0 30576 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2463_
timestamp 1698431365
transform -1 0 30688 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2464_
timestamp 1698431365
transform -1 0 30128 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2465_
timestamp 1698431365
transform -1 0 29008 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2466_
timestamp 1698431365
transform -1 0 28224 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1698431365
transform -1 0 33488 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2468_
timestamp 1698431365
transform 1 0 25648 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2469_
timestamp 1698431365
transform 1 0 25424 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2470_
timestamp 1698431365
transform -1 0 24864 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2471_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2472_
timestamp 1698431365
transform -1 0 24192 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2474_
timestamp 1698431365
transform 1 0 24080 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2475_
timestamp 1698431365
transform -1 0 23632 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2476_
timestamp 1698431365
transform -1 0 23408 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2477_
timestamp 1698431365
transform -1 0 22512 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2478_
timestamp 1698431365
transform -1 0 23072 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2479_
timestamp 1698431365
transform -1 0 22512 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2480_
timestamp 1698431365
transform -1 0 22624 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2481_
timestamp 1698431365
transform -1 0 22064 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2482_
timestamp 1698431365
transform -1 0 29344 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2483_
timestamp 1698431365
transform -1 0 26320 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2484_
timestamp 1698431365
transform -1 0 25648 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2485_
timestamp 1698431365
transform -1 0 16128 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2486_
timestamp 1698431365
transform -1 0 14896 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2487_
timestamp 1698431365
transform -1 0 15568 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2488_
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2489_
timestamp 1698431365
transform -1 0 15008 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2490_
timestamp 1698431365
transform -1 0 19376 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2491_
timestamp 1698431365
transform -1 0 14448 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2492_
timestamp 1698431365
transform -1 0 15456 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2493_
timestamp 1698431365
transform -1 0 14896 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2494_
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2495_
timestamp 1698431365
transform -1 0 14896 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2496_
timestamp 1698431365
transform -1 0 28000 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2497_
timestamp 1698431365
transform -1 0 24416 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2498_
timestamp 1698431365
transform -1 0 17024 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2499_
timestamp 1698431365
transform -1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1698431365
transform -1 0 17584 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2501_
timestamp 1698431365
transform -1 0 17024 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2502_
timestamp 1698431365
transform 1 0 17920 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2503_
timestamp 1698431365
transform -1 0 35616 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2504_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2505_
timestamp 1698431365
transform 1 0 17920 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2506_
timestamp 1698431365
transform 1 0 16800 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2507_
timestamp 1698431365
transform -1 0 16800 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2508_
timestamp 1698431365
transform -1 0 16800 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2509_
timestamp 1698431365
transform 1 0 27776 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2510_
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2511_
timestamp 1698431365
transform 1 0 21280 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1698431365
transform -1 0 24528 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2513_
timestamp 1698431365
transform 1 0 22288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2514_
timestamp 1698431365
transform 1 0 28560 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2515_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2516_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2517_
timestamp 1698431365
transform 1 0 38976 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2518_
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2519_
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2520_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2521_
timestamp 1698431365
transform -1 0 38192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2522_
timestamp 1698431365
transform -1 0 37520 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2523_
timestamp 1698431365
transform -1 0 40432 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2524_
timestamp 1698431365
transform 1 0 37968 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2525_
timestamp 1698431365
transform 1 0 38528 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2526_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2527_
timestamp 1698431365
transform -1 0 30688 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2528_
timestamp 1698431365
transform -1 0 30800 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2529_
timestamp 1698431365
transform -1 0 30688 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2530_
timestamp 1698431365
transform -1 0 32480 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2531_
timestamp 1698431365
transform 1 0 46816 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2532_
timestamp 1698431365
transform 1 0 44464 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2533_
timestamp 1698431365
transform 1 0 44016 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2534_
timestamp 1698431365
transform -1 0 44688 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2535_
timestamp 1698431365
transform 1 0 47712 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2536_
timestamp 1698431365
transform 1 0 46928 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2537_
timestamp 1698431365
transform 1 0 44912 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2538_
timestamp 1698431365
transform 1 0 45136 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2539_
timestamp 1698431365
transform -1 0 43232 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2540_
timestamp 1698431365
transform -1 0 44016 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2541_
timestamp 1698431365
transform 1 0 18816 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2542_
timestamp 1698431365
transform 1 0 22736 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2543_
timestamp 1698431365
transform 1 0 16464 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2544_
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2545_
timestamp 1698431365
transform 1 0 20496 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2546_
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2547_
timestamp 1698431365
transform 1 0 21504 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2548_
timestamp 1698431365
transform 1 0 16352 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2549_
timestamp 1698431365
transform 1 0 19936 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2550_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2551_
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2552_
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2553_
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2554_
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2555_
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2556_
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2557_
timestamp 1698431365
transform 1 0 2576 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2558_
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2559_
timestamp 1698431365
transform -1 0 21952 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2560_
timestamp 1698431365
transform 1 0 17696 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2561_
timestamp 1698431365
transform 1 0 4368 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2562_
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2563_
timestamp 1698431365
transform 1 0 5824 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2564_
timestamp 1698431365
transform -1 0 13104 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2565_
timestamp 1698431365
transform 1 0 5824 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2566_
timestamp 1698431365
transform 1 0 5040 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2567_
timestamp 1698431365
transform 1 0 6496 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2568_
timestamp 1698431365
transform 1 0 8176 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2569_
timestamp 1698431365
transform 1 0 9072 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2570_
timestamp 1698431365
transform 1 0 13328 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2571_
timestamp 1698431365
transform -1 0 20496 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2572_
timestamp 1698431365
transform 1 0 53424 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2573_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2574_
timestamp 1698431365
transform -1 0 58352 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2575_
timestamp 1698431365
transform 1 0 52864 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2576_
timestamp 1698431365
transform 1 0 49840 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2577_
timestamp 1698431365
transform 1 0 48944 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2578_
timestamp 1698431365
transform 1 0 50064 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2579_
timestamp 1698431365
transform -1 0 48496 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2580_
timestamp 1698431365
transform -1 0 50064 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2581_
timestamp 1698431365
transform 1 0 51184 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2582_
timestamp 1698431365
transform 1 0 49280 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2583_
timestamp 1698431365
transform 1 0 50512 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2584_
timestamp 1698431365
transform -1 0 55328 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2585_
timestamp 1698431365
transform 1 0 55104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2586_
timestamp 1698431365
transform -1 0 58240 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2587_
timestamp 1698431365
transform 1 0 55104 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2588_
timestamp 1698431365
transform 1 0 55104 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2589_
timestamp 1698431365
transform 1 0 55104 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2590_
timestamp 1698431365
transform 1 0 55104 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2591_
timestamp 1698431365
transform 1 0 53088 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2592_
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2593_
timestamp 1698431365
transform 1 0 48160 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2594_
timestamp 1698431365
transform -1 0 50064 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2595_
timestamp 1698431365
transform 1 0 42336 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2596_
timestamp 1698431365
transform 1 0 40880 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2597_
timestamp 1698431365
transform 1 0 42112 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2598_
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2599_
timestamp 1698431365
transform -1 0 45808 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2600_
timestamp 1698431365
transform -1 0 49168 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2601_
timestamp 1698431365
transform -1 0 49504 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2602_
timestamp 1698431365
transform 1 0 45024 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2603_
timestamp 1698431365
transform -1 0 36400 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2604_
timestamp 1698431365
transform -1 0 34160 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2605_
timestamp 1698431365
transform 1 0 25312 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2606_
timestamp 1698431365
transform 1 0 25088 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2607_
timestamp 1698431365
transform -1 0 34720 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2608_
timestamp 1698431365
transform 1 0 23856 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2609_
timestamp 1698431365
transform 1 0 27888 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2610_
timestamp 1698431365
transform -1 0 36624 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2611_
timestamp 1698431365
transform 1 0 21616 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2612_
timestamp 1698431365
transform -1 0 55776 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2613_
timestamp 1698431365
transform -1 0 57456 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2614_
timestamp 1698431365
transform -1 0 58352 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2615_
timestamp 1698431365
transform -1 0 57568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2616_
timestamp 1698431365
transform -1 0 56224 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2617_
timestamp 1698431365
transform -1 0 49840 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2618_
timestamp 1698431365
transform 1 0 43008 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2619_
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2620_
timestamp 1698431365
transform 1 0 39312 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2621_
timestamp 1698431365
transform 1 0 37632 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2622_
timestamp 1698431365
transform -1 0 28560 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2623_
timestamp 1698431365
transform -1 0 55776 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2624_
timestamp 1698431365
transform -1 0 55776 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2625_
timestamp 1698431365
transform -1 0 53648 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2626_
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2627_
timestamp 1698431365
transform -1 0 40096 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2628_
timestamp 1698431365
transform -1 0 37408 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2629_
timestamp 1698431365
transform 1 0 32592 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2630_
timestamp 1698431365
transform 1 0 29344 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2631_
timestamp 1698431365
transform 1 0 35056 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2632_
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2633_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8848 0 -1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2634_
timestamp 1698431365
transform -1 0 27776 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2635_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2636_
timestamp 1698431365
transform 1 0 21392 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2637_
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2638_
timestamp 1698431365
transform 1 0 15232 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2639_
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2640_
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2641_
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2642_
timestamp 1698431365
transform -1 0 24752 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2643_
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2644_
timestamp 1698431365
transform 1 0 15792 0 1 32928
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2645_
timestamp 1698431365
transform 1 0 45136 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2646_
timestamp 1698431365
transform 1 0 40544 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2647_
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2648_
timestamp 1698431365
transform 1 0 38640 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2649_
timestamp 1698431365
transform -1 0 41664 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2650_
timestamp 1698431365
transform 1 0 37408 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2651_
timestamp 1698431365
transform -1 0 47936 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2652_
timestamp 1698431365
transform 1 0 38304 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2653_
timestamp 1698431365
transform -1 0 44688 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2654_
timestamp 1698431365
transform 1 0 44688 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2655_
timestamp 1698431365
transform -1 0 58352 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2656_
timestamp 1698431365
transform -1 0 58352 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2657_
timestamp 1698431365
transform -1 0 58352 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2658_
timestamp 1698431365
transform 1 0 50624 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2659_
timestamp 1698431365
transform 1 0 55104 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2660_
timestamp 1698431365
transform 1 0 55104 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2661_
timestamp 1698431365
transform 1 0 54656 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2662_
timestamp 1698431365
transform 1 0 55104 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2663_
timestamp 1698431365
transform 1 0 36512 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2664_
timestamp 1698431365
transform -1 0 53984 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2665_
timestamp 1698431365
transform -1 0 49840 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2666_
timestamp 1698431365
transform 1 0 43456 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2667_
timestamp 1698431365
transform -1 0 50736 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2668_
timestamp 1698431365
transform 1 0 42336 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2669_
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2670_
timestamp 1698431365
transform -1 0 50176 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2671_
timestamp 1698431365
transform 1 0 46816 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2672_
timestamp 1698431365
transform 1 0 48608 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2673_
timestamp 1698431365
transform 1 0 48608 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2674_
timestamp 1698431365
transform -1 0 55104 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2675_
timestamp 1698431365
transform 1 0 51184 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2676_
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2677_
timestamp 1698431365
transform 1 0 49056 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2678_
timestamp 1698431365
transform 1 0 41104 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2679_
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2680_
timestamp 1698431365
transform 1 0 41216 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2681_
timestamp 1698431365
transform 1 0 37632 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2682_
timestamp 1698431365
transform 1 0 35056 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2683_
timestamp 1698431365
transform 1 0 33376 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2684_
timestamp 1698431365
transform 1 0 26432 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2685_
timestamp 1698431365
transform 1 0 26992 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2686_
timestamp 1698431365
transform 1 0 27664 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2687_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2688_
timestamp 1698431365
transform 1 0 29456 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2689_
timestamp 1698431365
transform 1 0 30464 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2690_
timestamp 1698431365
transform 1 0 15792 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2691_
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2692_
timestamp 1698431365
transform 1 0 15008 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2693_
timestamp 1698431365
transform 1 0 14112 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2694_
timestamp 1698431365
transform 1 0 19712 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2695_
timestamp 1698431365
transform 1 0 19264 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2696_
timestamp 1698431365
transform 1 0 30800 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2697_
timestamp 1698431365
transform 1 0 31024 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2698_
timestamp 1698431365
transform 1 0 27888 0 -1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2699_
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2700_
timestamp 1698431365
transform 1 0 23744 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2701_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2702_
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2703_
timestamp 1698431365
transform 1 0 19376 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2704_
timestamp 1698431365
transform 1 0 4144 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2705_
timestamp 1698431365
transform 1 0 4480 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2706_
timestamp 1698431365
transform 1 0 8400 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2707_
timestamp 1698431365
transform 1 0 9968 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2708_
timestamp 1698431365
transform 1 0 15232 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2709_
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2710_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2711_
timestamp 1698431365
transform -1 0 16912 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2712_
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2713_
timestamp 1698431365
transform 1 0 21504 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2714_
timestamp 1698431365
transform -1 0 31024 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_
timestamp 1698431365
transform 1 0 45472 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2716_
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1698431365
transform 1 0 38416 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__A3 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A3
timestamp 1698431365
transform 1 0 34496 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A1
timestamp 1698431365
transform -1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A2
timestamp 1698431365
transform -1 0 33264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A2
timestamp 1698431365
transform -1 0 22624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A2
timestamp 1698431365
transform -1 0 38640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A2
timestamp 1698431365
transform 1 0 22848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A3
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A1
timestamp 1698431365
transform 1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1698431365
transform 1 0 17472 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__I
timestamp 1698431365
transform 1 0 29120 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A2
timestamp 1698431365
transform 1 0 12320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1698431365
transform 1 0 33712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A2
timestamp 1698431365
transform -1 0 32592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A2
timestamp 1698431365
transform 1 0 13664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A2
timestamp 1698431365
transform -1 0 13776 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__A2
timestamp 1698431365
transform -1 0 33264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A1
timestamp 1698431365
transform 1 0 31920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A2
timestamp 1698431365
transform 1 0 12880 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__A2
timestamp 1698431365
transform -1 0 32592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__I
timestamp 1698431365
transform -1 0 31472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A1
timestamp 1698431365
transform 1 0 14560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A2
timestamp 1698431365
transform 1 0 13552 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__I
timestamp 1698431365
transform 1 0 11760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__I
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1698431365
transform 1 0 27664 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__I
timestamp 1698431365
transform -1 0 26208 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__I
timestamp 1698431365
transform 1 0 30464 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1698431365
transform 1 0 27440 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__I
timestamp 1698431365
transform 1 0 27776 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__I
timestamp 1698431365
transform 1 0 9632 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__I
timestamp 1698431365
transform 1 0 10752 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A2
timestamp 1698431365
transform -1 0 14000 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1698431365
transform 1 0 32256 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A2
timestamp 1698431365
transform 1 0 33600 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform 1 0 15792 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__I
timestamp 1698431365
transform 1 0 15344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__I
timestamp 1698431365
transform 1 0 14224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__A2
timestamp 1698431365
transform 1 0 13328 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__I
timestamp 1698431365
transform 1 0 31584 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__I
timestamp 1698431365
transform 1 0 30912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1698431365
transform -1 0 37408 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A2
timestamp 1698431365
transform 1 0 38640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__A1
timestamp 1698431365
transform 1 0 50400 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__I
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__I
timestamp 1698431365
transform 1 0 41888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__I
timestamp 1698431365
transform 1 0 29792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__I
timestamp 1698431365
transform 1 0 28112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1698431365
transform -1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1698431365
transform -1 0 35392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__C
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__I
timestamp 1698431365
transform -1 0 36064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform 1 0 35392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__I
timestamp 1698431365
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__I
timestamp 1698431365
transform -1 0 23072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__I
timestamp 1698431365
transform -1 0 42000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__B
timestamp 1698431365
transform 1 0 32480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1698431365
transform -1 0 31584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__I
timestamp 1698431365
transform 1 0 34384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__B
timestamp 1698431365
transform -1 0 30240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform 1 0 32032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1698431365
transform -1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__B
timestamp 1698431365
transform 1 0 32256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1698431365
transform -1 0 32144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__I
timestamp 1698431365
transform -1 0 39088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1698431365
transform 1 0 46816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__C
timestamp 1698431365
transform 1 0 46368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__B
timestamp 1698431365
transform 1 0 45808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A1
timestamp 1698431365
transform 1 0 44912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I
timestamp 1698431365
transform 1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__B
timestamp 1698431365
transform 1 0 45472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1698431365
transform 1 0 44912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__B
timestamp 1698431365
transform 1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1698431365
transform 1 0 43904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A1
timestamp 1698431365
transform 1 0 30800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1698431365
transform 1 0 47824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__C
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__B
timestamp 1698431365
transform 1 0 46592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1698431365
transform 1 0 46256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__B
timestamp 1698431365
transform -1 0 47376 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A1
timestamp 1698431365
transform 1 0 45248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__I
timestamp 1698431365
transform -1 0 22736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__I
timestamp 1698431365
transform 1 0 21840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__B
timestamp 1698431365
transform 1 0 46144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1698431365
transform 1 0 45360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__B
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__I
timestamp 1698431365
transform 1 0 49728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I
timestamp 1698431365
transform 1 0 49728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A1
timestamp 1698431365
transform 1 0 41664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1698431365
transform 1 0 23632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__B
timestamp 1698431365
transform 1 0 24080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__A1
timestamp 1698431365
transform 1 0 23184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__I
timestamp 1698431365
transform 1 0 49952 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__I
timestamp 1698431365
transform -1 0 25536 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__B
timestamp 1698431365
transform -1 0 23184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__B
timestamp 1698431365
transform 1 0 20944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__I
timestamp 1698431365
transform 1 0 8512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__B
timestamp 1698431365
transform 1 0 18256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__I
timestamp 1698431365
transform 1 0 22288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A1
timestamp 1698431365
transform 1 0 18368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__B
timestamp 1698431365
transform 1 0 20720 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__B
timestamp 1698431365
transform 1 0 4480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1698431365
transform 1 0 3248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A1
timestamp 1698431365
transform 1 0 3024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1698431365
transform 1 0 3136 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__B
timestamp 1698431365
transform 1 0 4592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__I
timestamp 1698431365
transform 1 0 7728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__B
timestamp 1698431365
transform 1 0 4592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__B
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__I
timestamp 1698431365
transform 1 0 21392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1698431365
transform 1 0 8176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__B
timestamp 1698431365
transform 1 0 7504 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1698431365
transform 1 0 20720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__I
timestamp 1698431365
transform 1 0 41776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__B
timestamp 1698431365
transform 1 0 20832 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__B
timestamp 1698431365
transform 1 0 6832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1698431365
transform -1 0 10416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__I
timestamp 1698431365
transform 1 0 8512 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1698431365
transform 1 0 14000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__I
timestamp 1698431365
transform -1 0 48608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1698431365
transform 1 0 12208 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform -1 0 13776 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1698431365
transform 1 0 15568 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__I
timestamp 1698431365
transform 1 0 25088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__I
timestamp 1698431365
transform -1 0 38752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__B
timestamp 1698431365
transform -1 0 18592 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A2
timestamp 1698431365
transform 1 0 53536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1698431365
transform 1 0 52976 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1698431365
transform 1 0 55104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1698431365
transform 1 0 53088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__I
timestamp 1698431365
transform -1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__A1
timestamp 1698431365
transform -1 0 50736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__I
timestamp 1698431365
transform 1 0 48832 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A1
timestamp 1698431365
transform 1 0 49616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A1
timestamp 1698431365
transform 1 0 50624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1698431365
transform -1 0 50736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1698431365
transform 1 0 48944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__I
timestamp 1698431365
transform 1 0 57568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A2
timestamp 1698431365
transform 1 0 58128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A2
timestamp 1698431365
transform 1 0 58128 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__I
timestamp 1698431365
transform 1 0 44800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A2
timestamp 1698431365
transform 1 0 45248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1698431365
transform -1 0 48272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1698431365
transform 1 0 57792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__I
timestamp 1698431365
transform -1 0 41552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__I
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__I
timestamp 1698431365
transform 1 0 37856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A2
timestamp 1698431365
transform -1 0 44016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A3
timestamp 1698431365
transform -1 0 45920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A1
timestamp 1698431365
transform 1 0 44352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__B
timestamp 1698431365
transform 1 0 42672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__I
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B
timestamp 1698431365
transform 1 0 44912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__B
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1698431365
transform 1 0 45472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A1
timestamp 1698431365
transform 1 0 47712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__B
timestamp 1698431365
transform -1 0 45360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform 1 0 44464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__B
timestamp 1698431365
transform 1 0 35616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__I
timestamp 1698431365
transform -1 0 38528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1698431365
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__B
timestamp 1698431365
transform 1 0 30464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__I
timestamp 1698431365
transform -1 0 27664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__B
timestamp 1698431365
transform 1 0 28448 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A1
timestamp 1698431365
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__B
timestamp 1698431365
transform 1 0 28560 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A2
timestamp 1698431365
transform 1 0 31248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__B
timestamp 1698431365
transform -1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A2
timestamp 1698431365
transform 1 0 30800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1698431365
transform 1 0 31472 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1698431365
transform 1 0 35504 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__C
timestamp 1698431365
transform 1 0 32816 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__I
timestamp 1698431365
transform -1 0 50736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A2
timestamp 1698431365
transform 1 0 52640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1698431365
transform 1 0 50624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__B
timestamp 1698431365
transform 1 0 51968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__I
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__I
timestamp 1698431365
transform -1 0 51184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__I
timestamp 1698431365
transform -1 0 38192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__I
timestamp 1698431365
transform 1 0 37520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__B
timestamp 1698431365
transform -1 0 51296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__C
timestamp 1698431365
transform 1 0 52752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__B
timestamp 1698431365
transform 1 0 51184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__C
timestamp 1698431365
transform -1 0 52752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__B
timestamp 1698431365
transform 1 0 52080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__I
timestamp 1698431365
transform 1 0 43344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__I
timestamp 1698431365
transform 1 0 49504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A1
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__I
timestamp 1698431365
transform 1 0 42784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A1
timestamp 1698431365
transform 1 0 42560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A2
timestamp 1698431365
transform 1 0 43680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__C
timestamp 1698431365
transform 1 0 43232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__A1
timestamp 1698431365
transform 1 0 38416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__I
timestamp 1698431365
transform 1 0 51408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__A1
timestamp 1698431365
transform 1 0 39984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A2
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__B
timestamp 1698431365
transform 1 0 42112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A1
timestamp 1698431365
transform -1 0 37968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A2
timestamp 1698431365
transform 1 0 39200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A1
timestamp 1698431365
transform -1 0 37856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__A2
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__B
timestamp 1698431365
transform 1 0 28336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__A2
timestamp 1698431365
transform -1 0 27664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__A2
timestamp 1698431365
transform 1 0 52416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1698431365
transform 1 0 50400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__B
timestamp 1698431365
transform -1 0 51408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__I
timestamp 1698431365
transform 1 0 42560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__I
timestamp 1698431365
transform 1 0 38976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__I
timestamp 1698431365
transform -1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1698431365
transform -1 0 33376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A1
timestamp 1698431365
transform -1 0 33824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A2
timestamp 1698431365
transform -1 0 33600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__C
timestamp 1698431365
transform -1 0 34048 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__A1
timestamp 1698431365
transform 1 0 35728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__A1
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__A2
timestamp 1698431365
transform 1 0 35056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__B
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A1
timestamp 1698431365
transform 1 0 33040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A2
timestamp 1698431365
transform -1 0 33600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1698431365
transform 1 0 36064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__I
timestamp 1698431365
transform -1 0 39424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A2
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__B
timestamp 1698431365
transform -1 0 11648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A2
timestamp 1698431365
transform 1 0 8400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A2
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A1
timestamp 1698431365
transform -1 0 25984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__B
timestamp 1698431365
transform -1 0 27664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__I
timestamp 1698431365
transform 1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2210__I
timestamp 1698431365
transform 1 0 24528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__I
timestamp 1698431365
transform 1 0 22176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A2
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1698431365
transform -1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1698431365
transform -1 0 20272 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__A1
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A2
timestamp 1698431365
transform -1 0 22176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__C
timestamp 1698431365
transform 1 0 22176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A1
timestamp 1698431365
transform 1 0 24304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A1
timestamp 1698431365
transform -1 0 24304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__A2
timestamp 1698431365
transform -1 0 23408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__B
timestamp 1698431365
transform 1 0 25200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A1
timestamp 1698431365
transform 1 0 22624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__A2
timestamp 1698431365
transform 1 0 22400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__A1
timestamp 1698431365
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A2
timestamp 1698431365
transform 1 0 21056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__B
timestamp 1698431365
transform 1 0 21280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__A2
timestamp 1698431365
transform 1 0 19824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__B
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A1
timestamp 1698431365
transform 1 0 33488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A2
timestamp 1698431365
transform -1 0 34160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A2
timestamp 1698431365
transform -1 0 37968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A1
timestamp 1698431365
transform 1 0 42112 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__B
timestamp 1698431365
transform 1 0 45920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1698431365
transform 1 0 41664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1698431365
transform 1 0 42224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2285__A2
timestamp 1698431365
transform 1 0 39536 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2288__I
timestamp 1698431365
transform -1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__B
timestamp 1698431365
transform 1 0 40992 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1698431365
transform 1 0 45696 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__B
timestamp 1698431365
transform 1 0 41888 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A1
timestamp 1698431365
transform 1 0 43792 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__B
timestamp 1698431365
transform 1 0 44912 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1698431365
transform 1 0 56000 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A2
timestamp 1698431365
transform 1 0 56000 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__C
timestamp 1698431365
transform 1 0 55552 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__C
timestamp 1698431365
transform -1 0 53984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__A1
timestamp 1698431365
transform 1 0 51520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__B
timestamp 1698431365
transform 1 0 51632 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1698431365
transform 1 0 52080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A2
timestamp 1698431365
transform 1 0 47824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A2
timestamp 1698431365
transform 1 0 47488 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A2
timestamp 1698431365
transform 1 0 45808 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A2
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A2
timestamp 1698431365
transform 1 0 44128 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__C2
timestamp 1698431365
transform 1 0 45472 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A2
timestamp 1698431365
transform 1 0 51072 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1698431365
transform -1 0 51296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__I
timestamp 1698431365
transform 1 0 32032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__I
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__B
timestamp 1698431365
transform -1 0 43232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__I
timestamp 1698431365
transform 1 0 23632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A1
timestamp 1698431365
transform 1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1698431365
transform 1 0 39760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__A1
timestamp 1698431365
transform 1 0 37744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__I
timestamp 1698431365
transform -1 0 33936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__A2
timestamp 1698431365
transform -1 0 27776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__A1
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__I
timestamp 1698431365
transform 1 0 35952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1698431365
transform -1 0 27664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__I
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A1
timestamp 1698431365
transform 1 0 30128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__I
timestamp 1698431365
transform 1 0 19600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A1
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A1
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1698431365
transform 1 0 19264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A1
timestamp 1698431365
transform -1 0 18368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A1
timestamp 1698431365
transform -1 0 19152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__B
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A1
timestamp 1698431365
transform -1 0 27888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A2
timestamp 1698431365
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A1
timestamp 1698431365
transform 1 0 32032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__C
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A1
timestamp 1698431365
transform 1 0 31920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A1
timestamp 1698431365
transform 1 0 29232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__A1
timestamp 1698431365
transform 1 0 26880 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A1
timestamp 1698431365
transform -1 0 25536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1698431365
transform -1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A1
timestamp 1698431365
transform 1 0 21168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A1
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A2
timestamp 1698431365
transform 1 0 29344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A1
timestamp 1698431365
transform 1 0 15792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2490__I
timestamp 1698431365
transform 1 0 19600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A1
timestamp 1698431365
transform 1 0 15792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A1
timestamp 1698431365
transform 1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__A1
timestamp 1698431365
transform 1 0 17808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__A1
timestamp 1698431365
transform 1 0 18480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__I
timestamp 1698431365
transform -1 0 35840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A1
timestamp 1698431365
transform 1 0 18592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__C
timestamp 1698431365
transform -1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__A1
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__C
timestamp 1698431365
transform 1 0 18592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1698431365
transform -1 0 15680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__C
timestamp 1698431365
transform -1 0 16240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__B
timestamp 1698431365
transform -1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A1
timestamp 1698431365
transform -1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__B
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__C
timestamp 1698431365
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1698431365
transform 1 0 42448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__B
timestamp 1698431365
transform -1 0 37744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A1
timestamp 1698431365
transform -1 0 36848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1698431365
transform -1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2524__A1
timestamp 1698431365
transform 1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__C
timestamp 1698431365
transform 1 0 37744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__CLK
timestamp 1698431365
transform 1 0 42000 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__D
timestamp 1698431365
transform 1 0 41552 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2527__CLK
timestamp 1698431365
transform 1 0 30688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__CLK
timestamp 1698431365
transform 1 0 31808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__CLK
timestamp 1698431365
transform 1 0 31584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__CLK
timestamp 1698431365
transform 1 0 50288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__CLK
timestamp 1698431365
transform -1 0 44016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__CLK
timestamp 1698431365
transform 1 0 41216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__CLK
timestamp 1698431365
transform 1 0 51184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__CLK
timestamp 1698431365
transform -1 0 50400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__CLK
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__CLK
timestamp 1698431365
transform 1 0 44912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__CLK
timestamp 1698431365
transform 1 0 43456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__CLK
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__CLK
timestamp 1698431365
transform 1 0 22512 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__CLK
timestamp 1698431365
transform 1 0 19040 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__CLK
timestamp 1698431365
transform -1 0 21616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__CLK
timestamp 1698431365
transform 1 0 25872 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__CLK
timestamp 1698431365
transform 1 0 16128 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__CLK
timestamp 1698431365
transform 1 0 23408 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__CLK
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__CLK
timestamp 1698431365
transform 1 0 5488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__CLK
timestamp 1698431365
transform 1 0 5040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__CLK
timestamp 1698431365
transform 1 0 5376 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__CLK
timestamp 1698431365
transform -1 0 5152 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2556__CLK
timestamp 1698431365
transform 1 0 4816 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__CLK
timestamp 1698431365
transform 1 0 5824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__CLK
timestamp 1698431365
transform -1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__CLK
timestamp 1698431365
transform 1 0 21952 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__CLK
timestamp 1698431365
transform 1 0 21392 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__CLK
timestamp 1698431365
transform 1 0 7840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__CLK
timestamp 1698431365
transform 1 0 8400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__CLK
timestamp 1698431365
transform 1 0 9520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__CLK
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__CLK
timestamp 1698431365
transform 1 0 10192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__CLK
timestamp 1698431365
transform -1 0 9856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__CLK
timestamp 1698431365
transform 1 0 9744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__CLK
timestamp 1698431365
transform 1 0 11312 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__CLK
timestamp 1698431365
transform -1 0 12544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__CLK
timestamp 1698431365
transform -1 0 20944 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__CLK
timestamp 1698431365
transform 1 0 56224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__CLK
timestamp 1698431365
transform 1 0 54880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__CLK
timestamp 1698431365
transform 1 0 53312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__CLK
timestamp 1698431365
transform 1 0 52416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__CLK
timestamp 1698431365
transform 1 0 53536 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__CLK
timestamp 1698431365
transform 1 0 48720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__CLK
timestamp 1698431365
transform 1 0 50848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__CLK
timestamp 1698431365
transform 1 0 54656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__CLK
timestamp 1698431365
transform 1 0 53312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__CLK
timestamp 1698431365
transform 1 0 54656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__CLK
timestamp 1698431365
transform 1 0 55552 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__CLK
timestamp 1698431365
transform 1 0 58128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__CLK
timestamp 1698431365
transform 1 0 58128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__CLK
timestamp 1698431365
transform 1 0 58128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__CLK
timestamp 1698431365
transform 1 0 58128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__CLK
timestamp 1698431365
transform 1 0 58128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__CLK
timestamp 1698431365
transform 1 0 54880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__CLK
timestamp 1698431365
transform -1 0 56784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__CLK
timestamp 1698431365
transform 1 0 56000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__CLK
timestamp 1698431365
transform 1 0 51408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__CLK
timestamp 1698431365
transform 1 0 50288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__CLK
timestamp 1698431365
transform 1 0 42896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__CLK
timestamp 1698431365
transform 1 0 44352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__CLK
timestamp 1698431365
transform 1 0 45584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__CLK
timestamp 1698431365
transform 1 0 42112 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__CLK
timestamp 1698431365
transform -1 0 42560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__CLK
timestamp 1698431365
transform 1 0 49952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__CLK
timestamp 1698431365
transform 1 0 49728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__CLK
timestamp 1698431365
transform 1 0 44800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__CLK
timestamp 1698431365
transform 1 0 34384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__CLK
timestamp 1698431365
transform 1 0 25088 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__CLK
timestamp 1698431365
transform 1 0 34944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__CLK
timestamp 1698431365
transform 1 0 23184 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__CLK
timestamp 1698431365
transform 1 0 27664 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__CLK
timestamp 1698431365
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__CLK
timestamp 1698431365
transform -1 0 25536 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__CLK
timestamp 1698431365
transform 1 0 56000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__CLK
timestamp 1698431365
transform 1 0 57456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__CLK
timestamp 1698431365
transform 1 0 58128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__CLK
timestamp 1698431365
transform 1 0 57792 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__CLK
timestamp 1698431365
transform 1 0 56672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__CLK
timestamp 1698431365
transform 1 0 50064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__CLK
timestamp 1698431365
transform 1 0 42784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__CLK
timestamp 1698431365
transform 1 0 41440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__CLK
timestamp 1698431365
transform 1 0 43008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__CLK
timestamp 1698431365
transform 1 0 56000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__CLK
timestamp 1698431365
transform 1 0 56000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__CLK
timestamp 1698431365
transform 1 0 53872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__CLK
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__CLK
timestamp 1698431365
transform 1 0 40320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__CLK
timestamp 1698431365
transform 1 0 37632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__CLK
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__CLK
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__CLK
timestamp 1698431365
transform 1 0 38304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__CLK
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__CLK
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__CLK
timestamp 1698431365
transform 1 0 28336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__CLK
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__CLK
timestamp 1698431365
transform -1 0 21616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__CLK
timestamp 1698431365
transform 1 0 18368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__CLK
timestamp 1698431365
transform 1 0 17696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__CLK
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__CLK
timestamp 1698431365
transform -1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__CLK
timestamp 1698431365
transform 1 0 43792 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__CLK
timestamp 1698431365
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__CLK
timestamp 1698431365
transform 1 0 42112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__CLK
timestamp 1698431365
transform 1 0 42784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__CLK
timestamp 1698431365
transform 1 0 48160 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__CLK
timestamp 1698431365
transform 1 0 41776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__CLK
timestamp 1698431365
transform 1 0 45360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__CLK
timestamp 1698431365
transform 1 0 44912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__CLK
timestamp 1698431365
transform 1 0 54880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__CLK
timestamp 1698431365
transform 1 0 54880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2657__CLK
timestamp 1698431365
transform 1 0 53984 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2658__CLK
timestamp 1698431365
transform 1 0 53872 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__CLK
timestamp 1698431365
transform 1 0 54880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__CLK
timestamp 1698431365
transform 1 0 54880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__CLK
timestamp 1698431365
transform 1 0 58128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__CLK
timestamp 1698431365
transform 1 0 54992 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__CLK
timestamp 1698431365
transform -1 0 41216 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__D
timestamp 1698431365
transform -1 0 40208 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__CLK
timestamp 1698431365
transform 1 0 54208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__CLK
timestamp 1698431365
transform 1 0 49840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__CLK
timestamp 1698431365
transform 1 0 43232 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__CLK
timestamp 1698431365
transform -1 0 51856 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__CLK
timestamp 1698431365
transform 1 0 45808 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__CLK
timestamp 1698431365
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__CLK
timestamp 1698431365
transform 1 0 50400 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__CLK
timestamp 1698431365
transform 1 0 50400 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__CLK
timestamp 1698431365
transform 1 0 52080 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__CLK
timestamp 1698431365
transform 1 0 52752 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__CLK
timestamp 1698431365
transform -1 0 55552 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__CLK
timestamp 1698431365
transform 1 0 54656 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__CLK
timestamp 1698431365
transform 1 0 54208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2677__CLK
timestamp 1698431365
transform -1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__CLK
timestamp 1698431365
transform -1 0 45584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__CLK
timestamp 1698431365
transform -1 0 41664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__CLK
timestamp 1698431365
transform 1 0 41440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__CLK
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__CLK
timestamp 1698431365
transform 1 0 33152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__CLK
timestamp 1698431365
transform 1 0 29904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__CLK
timestamp 1698431365
transform 1 0 30464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__CLK
timestamp 1698431365
transform 1 0 30912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__CLK
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__CLK
timestamp 1698431365
transform 1 0 33936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__CLK
timestamp 1698431365
transform 1 0 19712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__CLK
timestamp 1698431365
transform 1 0 14784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__CLK
timestamp 1698431365
transform -1 0 17808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__CLK
timestamp 1698431365
transform -1 0 19712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__CLK
timestamp 1698431365
transform 1 0 18032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__CLK
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__CLK
timestamp 1698431365
transform 1 0 30240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__CLK
timestamp 1698431365
transform 1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__CLK
timestamp 1698431365
transform 1 0 29680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__CLK
timestamp 1698431365
transform 1 0 27216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__CLK
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__CLK
timestamp 1698431365
transform 1 0 24640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__CLK
timestamp 1698431365
transform 1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__CLK
timestamp 1698431365
transform 1 0 6944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__CLK
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__CLK
timestamp 1698431365
transform 1 0 13440 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__CLK
timestamp 1698431365
transform 1 0 15008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__CLK
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__CLK
timestamp 1698431365
transform 1 0 16576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__CLK
timestamp 1698431365
transform 1 0 23968 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__CLK
timestamp 1698431365
transform -1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__CLK
timestamp 1698431365
transform 1 0 27552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__CLK
timestamp 1698431365
transform 1 0 45248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__CLK
timestamp 1698431365
transform 1 0 38416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__CLK
timestamp 1698431365
transform 1 0 40320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__CLK
timestamp 1698431365
transform 1 0 41888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 28224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 38752 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 39984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 53872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 12432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 20944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 14448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 25648 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 52752 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 39984 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 52528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 58352 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 57680 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 57456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 58128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 58352 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 57680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 57904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 57680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 58352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 57456 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 1792 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 1792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1698431365
transform -1 0 30352 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1698431365
transform 1 0 39424 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1698431365
transform 1 0 43008 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698431365
transform 1 0 29568 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698431365
transform 1 0 12544 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698431365
transform 1 0 38976 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698431365
transform 1 0 53200 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698431365
transform 1 0 40208 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698431365
transform 1 0 54096 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698431365
transform -1 0 12432 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698431365
transform 1 0 18032 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698431365
transform 1 0 11536 0 -1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698431365
transform 1 0 21952 0 -1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698431365
transform 1 0 41216 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698431365
transform 1 0 52976 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698431365
transform 1 0 41104 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698431365
transform 1 0 52752 0 1 58016
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_178 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_181 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_197
timestamp 1698431365
transform 1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_378
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_381
timestamp 1698431365
transform 1 0 44016 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_397 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_405
timestamp 1698431365
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_241
timestamp 1698431365
transform 1 0 28336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_245
timestamp 1698431365
transform 1 0 28784 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_290
timestamp 1698431365
transform 1 0 33824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_292
timestamp 1698431365
transform 1 0 34048 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_322
timestamp 1698431365
transform 1 0 37408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_326
timestamp 1698431365
transform 1 0 37856 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_331
timestamp 1698431365
transform 1 0 38416 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_347
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_410
timestamp 1698431365
transform 1 0 47264 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_418
timestamp 1698431365
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_426
timestamp 1698431365
transform 1 0 49056 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_434
timestamp 1698431365
transform 1 0 49952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_467
timestamp 1698431365
transform 1 0 53648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_471
timestamp 1698431365
transform 1 0 54096 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_487
timestamp 1698431365
transform 1 0 55888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_496
timestamp 1698431365
transform 1 0 56896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_498
timestamp 1698431365
transform 1 0 57120 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_139
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_155
timestamp 1698431365
transform 1 0 18704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_163
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_165
timestamp 1698431365
transform 1 0 19824 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_170
timestamp 1698431365
transform 1 0 20384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_189
timestamp 1698431365
transform 1 0 22512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_197
timestamp 1698431365
transform 1 0 23408 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_213
timestamp 1698431365
transform 1 0 25200 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_217
timestamp 1698431365
transform 1 0 25648 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_255
timestamp 1698431365
transform 1 0 29904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_259
timestamp 1698431365
transform 1 0 30352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_268
timestamp 1698431365
transform 1 0 31360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_272
timestamp 1698431365
transform 1 0 31808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_276
timestamp 1698431365
transform 1 0 32256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_278
timestamp 1698431365
transform 1 0 32480 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_308
timestamp 1698431365
transform 1 0 35840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_346
timestamp 1698431365
transform 1 0 40096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_354
timestamp 1698431365
transform 1 0 40992 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_370
timestamp 1698431365
transform 1 0 42784 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_378
timestamp 1698431365
transform 1 0 43680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_380
timestamp 1698431365
transform 1 0 43904 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_383
timestamp 1698431365
transform 1 0 44240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_391
timestamp 1698431365
transform 1 0 45136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_393
timestamp 1698431365
transform 1 0 45360 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_404
timestamp 1698431365
transform 1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_435
timestamp 1698431365
transform 1 0 50064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_439
timestamp 1698431365
transform 1 0 50512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_443
timestamp 1698431365
transform 1 0 50960 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_448
timestamp 1698431365
transform 1 0 51520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1698431365
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698431365
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_146
timestamp 1698431365
transform 1 0 17696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_162
timestamp 1698431365
transform 1 0 19488 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_178
timestamp 1698431365
transform 1 0 21280 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_187
timestamp 1698431365
transform 1 0 22288 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_205
timestamp 1698431365
transform 1 0 24304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_228
timestamp 1698431365
transform 1 0 26880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_232
timestamp 1698431365
transform 1 0 27328 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_262
timestamp 1698431365
transform 1 0 30688 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_271
timestamp 1698431365
transform 1 0 31696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_286
timestamp 1698431365
transform 1 0 33376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_292
timestamp 1698431365
transform 1 0 34048 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_300
timestamp 1698431365
transform 1 0 34944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_302
timestamp 1698431365
transform 1 0 35168 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_307
timestamp 1698431365
transform 1 0 35728 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_339
timestamp 1698431365
transform 1 0 39312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_387
timestamp 1698431365
transform 1 0 44688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_397
timestamp 1698431365
transform 1 0 45808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_414
timestamp 1698431365
transform 1 0 47712 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_418
timestamp 1698431365
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_165
timestamp 1698431365
transform 1 0 19824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_193
timestamp 1698431365
transform 1 0 22960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_195
timestamp 1698431365
transform 1 0 23184 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_216
timestamp 1698431365
transform 1 0 25536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_236
timestamp 1698431365
transform 1 0 27776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_240
timestamp 1698431365
transform 1 0 28224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_255
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_274
timestamp 1698431365
transform 1 0 32032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_278
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_312
timestamp 1698431365
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698431365
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_337
timestamp 1698431365
transform 1 0 39088 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_341
timestamp 1698431365
transform 1 0 39536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_363
timestamp 1698431365
transform 1 0 42000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_367
timestamp 1698431365
transform 1 0 42448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_369
timestamp 1698431365
transform 1 0 42672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_378
timestamp 1698431365
transform 1 0 43680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_382
timestamp 1698431365
transform 1 0 44128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_395
timestamp 1698431365
transform 1 0 45584 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_399
timestamp 1698431365
transform 1 0 46032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_401
timestamp 1698431365
transform 1 0 46256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_404
timestamp 1698431365
transform 1 0 46592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_408
timestamp 1698431365
transform 1 0 47040 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_416
timestamp 1698431365
transform 1 0 47936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_426
timestamp 1698431365
transform 1 0 49056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_448
timestamp 1698431365
transform 1 0 51520 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_452
timestamp 1698431365
transform 1 0 51968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_454
timestamp 1698431365
transform 1 0 52192 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_486
timestamp 1698431365
transform 1 0 55776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_490
timestamp 1698431365
transform 1 0 56224 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_506
timestamp 1698431365
transform 1 0 58016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_508
timestamp 1698431365
transform 1 0 58240 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_170
timestamp 1698431365
transform 1 0 20384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_180
timestamp 1698431365
transform 1 0 21504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_188
timestamp 1698431365
transform 1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_233
timestamp 1698431365
transform 1 0 27440 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_263
timestamp 1698431365
transform 1 0 30800 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_267
timestamp 1698431365
transform 1 0 31248 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_270
timestamp 1698431365
transform 1 0 31584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_274
timestamp 1698431365
transform 1 0 32032 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_278
timestamp 1698431365
transform 1 0 32480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_298
timestamp 1698431365
transform 1 0 34720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_318
timestamp 1698431365
transform 1 0 36960 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_338
timestamp 1698431365
transform 1 0 39200 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_360
timestamp 1698431365
transform 1 0 41664 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_384
timestamp 1698431365
transform 1 0 44352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_388
timestamp 1698431365
transform 1 0 44800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_396
timestamp 1698431365
transform 1 0 45696 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_399
timestamp 1698431365
transform 1 0 46032 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_415
timestamp 1698431365
transform 1 0 47824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_419
timestamp 1698431365
transform 1 0 48272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_450
timestamp 1698431365
transform 1 0 51744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_454
timestamp 1698431365
transform 1 0 52192 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_459
timestamp 1698431365
transform 1 0 52752 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_475
timestamp 1698431365
transform 1 0 54544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_483
timestamp 1698431365
transform 1 0 55440 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_487
timestamp 1698431365
transform 1 0 55888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_489
timestamp 1698431365
transform 1 0 56112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_233
timestamp 1698431365
transform 1 0 27440 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_259
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_276
timestamp 1698431365
transform 1 0 32256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_280
timestamp 1698431365
transform 1 0 32704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_284
timestamp 1698431365
transform 1 0 33152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_286
timestamp 1698431365
transform 1 0 33376 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_293
timestamp 1698431365
transform 1 0 34160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_297
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_333
timestamp 1698431365
transform 1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_335
timestamp 1698431365
transform 1 0 38864 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_344
timestamp 1698431365
transform 1 0 39872 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_376
timestamp 1698431365
transform 1 0 43456 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1698431365
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_407
timestamp 1698431365
transform 1 0 46928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_450
timestamp 1698431365
transform 1 0 51744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698431365
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_104
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_120
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_124
timestamp 1698431365
transform 1 0 15232 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_126
timestamp 1698431365
transform 1 0 15456 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_131
timestamp 1698431365
transform 1 0 16016 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_162
timestamp 1698431365
transform 1 0 19488 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_178
timestamp 1698431365
transform 1 0 21280 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_182
timestamp 1698431365
transform 1 0 21728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_228
timestamp 1698431365
transform 1 0 26880 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_232
timestamp 1698431365
transform 1 0 27328 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_235
timestamp 1698431365
transform 1 0 27664 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_251
timestamp 1698431365
transform 1 0 29456 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_259
timestamp 1698431365
transform 1 0 30352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_263
timestamp 1698431365
transform 1 0 30800 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_270
timestamp 1698431365
transform 1 0 31584 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_291
timestamp 1698431365
transform 1 0 33936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_307
timestamp 1698431365
transform 1 0 35728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_315
timestamp 1698431365
transform 1 0 36624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_317
timestamp 1698431365
transform 1 0 36848 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_326
timestamp 1698431365
transform 1 0 37856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_334
timestamp 1698431365
transform 1 0 38752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_336
timestamp 1698431365
transform 1 0 38976 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698431365
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_360
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_381
timestamp 1698431365
transform 1 0 44016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_414
timestamp 1698431365
transform 1 0 47712 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_418
timestamp 1698431365
transform 1 0 48160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_430
timestamp 1698431365
transform 1 0 49504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_440
timestamp 1698431365
transform 1 0 50624 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_444
timestamp 1698431365
transform 1 0 51072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_447
timestamp 1698431365
transform 1 0 51408 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_479
timestamp 1698431365
transform 1 0 54992 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_487
timestamp 1698431365
transform 1 0 55888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_489
timestamp 1698431365
transform 1 0 56112 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_144
timestamp 1698431365
transform 1 0 17472 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_165
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_169
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_184
timestamp 1698431365
transform 1 0 21952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_188
timestamp 1698431365
transform 1 0 22400 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_192
timestamp 1698431365
transform 1 0 22848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_194
timestamp 1698431365
transform 1 0 23072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_251
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_253
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_274
timestamp 1698431365
transform 1 0 32032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_297
timestamp 1698431365
transform 1 0 34608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_301
timestamp 1698431365
transform 1 0 35056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_321
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_360
timestamp 1698431365
transform 1 0 41664 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_419
timestamp 1698431365
transform 1 0 48272 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_435
timestamp 1698431365
transform 1 0 50064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_437
timestamp 1698431365
transform 1 0 50288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_445
timestamp 1698431365
transform 1 0 51184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_486
timestamp 1698431365
transform 1 0 55776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_490
timestamp 1698431365
transform 1 0 56224 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_506
timestamp 1698431365
transform 1 0 58016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_508
timestamp 1698431365
transform 1 0 58240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_104
timestamp 1698431365
transform 1 0 12992 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_124
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_126
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_131
timestamp 1698431365
transform 1 0 16016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_174
timestamp 1698431365
transform 1 0 20832 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_178
timestamp 1698431365
transform 1 0 21280 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_216
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_262
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_269
timestamp 1698431365
transform 1 0 31472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_273
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_356
timestamp 1698431365
transform 1 0 41216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_358
timestamp 1698431365
transform 1 0 41440 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_367
timestamp 1698431365
transform 1 0 42448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_369
timestamp 1698431365
transform 1 0 42672 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_401
timestamp 1698431365
transform 1 0 46256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_411
timestamp 1698431365
transform 1 0 47376 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_419
timestamp 1698431365
transform 1 0 48272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_438
timestamp 1698431365
transform 1 0 50400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_442
timestamp 1698431365
transform 1 0 50848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_444
timestamp 1698431365
transform 1 0 51072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_450
timestamp 1698431365
transform 1 0 51744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_454
timestamp 1698431365
transform 1 0 52192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_458
timestamp 1698431365
transform 1 0 52640 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_500
timestamp 1698431365
transform 1 0 57344 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_504
timestamp 1698431365
transform 1 0 57792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_506
timestamp 1698431365
transform 1 0 58016 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_144
timestamp 1698431365
transform 1 0 17472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_148
timestamp 1698431365
transform 1 0 17920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_152
timestamp 1698431365
transform 1 0 18368 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_165
timestamp 1698431365
transform 1 0 19824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_169
timestamp 1698431365
transform 1 0 20272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_183
timestamp 1698431365
transform 1 0 21840 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_199
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_259
timestamp 1698431365
transform 1 0 30352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_261
timestamp 1698431365
transform 1 0 30576 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_264
timestamp 1698431365
transform 1 0 30912 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_268
timestamp 1698431365
transform 1 0 31360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_280
timestamp 1698431365
transform 1 0 32704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_284
timestamp 1698431365
transform 1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_288
timestamp 1698431365
transform 1 0 33600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_292
timestamp 1698431365
transform 1 0 34048 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_300
timestamp 1698431365
transform 1 0 34944 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_303
timestamp 1698431365
transform 1 0 35280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_328
timestamp 1698431365
transform 1 0 38080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_338
timestamp 1698431365
transform 1 0 39200 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_370
timestamp 1698431365
transform 1 0 42784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_374
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_403
timestamp 1698431365
transform 1 0 46480 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_433
timestamp 1698431365
transform 1 0 49840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_437
timestamp 1698431365
transform 1 0 50288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_441
timestamp 1698431365
transform 1 0 50736 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_486
timestamp 1698431365
transform 1 0 55776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_490
timestamp 1698431365
transform 1 0 56224 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_502
timestamp 1698431365
transform 1 0 57568 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_171
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_175
timestamp 1698431365
transform 1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_179
timestamp 1698431365
transform 1 0 21392 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_197
timestamp 1698431365
transform 1 0 23408 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_201
timestamp 1698431365
transform 1 0 23856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_205
timestamp 1698431365
transform 1 0 24304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_228
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_235
timestamp 1698431365
transform 1 0 27664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_239
timestamp 1698431365
transform 1 0 28112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_243
timestamp 1698431365
transform 1 0 28560 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_251
timestamp 1698431365
transform 1 0 29456 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_292
timestamp 1698431365
transform 1 0 34048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_332
timestamp 1698431365
transform 1 0 38528 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_358
timestamp 1698431365
transform 1 0 41440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_362
timestamp 1698431365
transform 1 0 41888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_366
timestamp 1698431365
transform 1 0 42336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_370
timestamp 1698431365
transform 1 0 42784 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_378
timestamp 1698431365
transform 1 0 43680 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_382
timestamp 1698431365
transform 1 0 44128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_384
timestamp 1698431365
transform 1 0 44352 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_389
timestamp 1698431365
transform 1 0 44912 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_405
timestamp 1698431365
transform 1 0 46704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_417
timestamp 1698431365
transform 1 0 48048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1698431365
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_430
timestamp 1698431365
transform 1 0 49504 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_456
timestamp 1698431365
transform 1 0 52416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_460
timestamp 1698431365
transform 1 0 52864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_462
timestamp 1698431365
transform 1 0 53088 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_489
timestamp 1698431365
transform 1 0 56112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698431365
transform 1 0 17360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_183
timestamp 1698431365
transform 1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_211
timestamp 1698431365
transform 1 0 24976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_215
timestamp 1698431365
transform 1 0 25424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_249
timestamp 1698431365
transform 1 0 29232 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_293
timestamp 1698431365
transform 1 0 34160 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_310
timestamp 1698431365
transform 1 0 36064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_333
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_368
timestamp 1698431365
transform 1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_372
timestamp 1698431365
transform 1 0 43008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_374
timestamp 1698431365
transform 1 0 43232 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_399
timestamp 1698431365
transform 1 0 46032 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_407
timestamp 1698431365
transform 1 0 46928 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_420
timestamp 1698431365
transform 1 0 48384 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_436
timestamp 1698431365
transform 1 0 50176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_440
timestamp 1698431365
transform 1 0 50624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_442
timestamp 1698431365
transform 1 0 50848 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_445
timestamp 1698431365
transform 1 0 51184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_449
timestamp 1698431365
transform 1 0 51632 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_453
timestamp 1698431365
transform 1 0 52080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_463
timestamp 1698431365
transform 1 0 53200 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_495
timestamp 1698431365
transform 1 0 56784 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_503
timestamp 1698431365
transform 1 0 57680 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_507
timestamp 1698431365
transform 1 0 58128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698431365
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698431365
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_184
timestamp 1698431365
transform 1 0 21952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_203
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_228
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_258
timestamp 1698431365
transform 1 0 30240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_262
timestamp 1698431365
transform 1 0 30688 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_270
timestamp 1698431365
transform 1 0 31584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_288
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_305
timestamp 1698431365
transform 1 0 35504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_309
timestamp 1698431365
transform 1 0 35952 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_317
timestamp 1698431365
transform 1 0 36848 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_321
timestamp 1698431365
transform 1 0 37296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_325
timestamp 1698431365
transform 1 0 37744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_329
timestamp 1698431365
transform 1 0 38192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_333
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_372
timestamp 1698431365
transform 1 0 43008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_376
timestamp 1698431365
transform 1 0 43456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_385
timestamp 1698431365
transform 1 0 44464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_393
timestamp 1698431365
transform 1 0 45360 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_417
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_430
timestamp 1698431365
transform 1 0 49504 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_434
timestamp 1698431365
transform 1 0 49952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_444
timestamp 1698431365
transform 1 0 51072 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_452
timestamp 1698431365
transform 1 0 51968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_456
timestamp 1698431365
transform 1 0 52416 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_496
timestamp 1698431365
transform 1 0 56896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_504
timestamp 1698431365
transform 1 0 57792 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_149
timestamp 1698431365
transform 1 0 18032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_158
timestamp 1698431365
transform 1 0 19040 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_183
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_186
timestamp 1698431365
transform 1 0 22176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_192
timestamp 1698431365
transform 1 0 22848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_194
timestamp 1698431365
transform 1 0 23072 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_232
timestamp 1698431365
transform 1 0 27328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_279
timestamp 1698431365
transform 1 0 32592 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_287
timestamp 1698431365
transform 1 0 33488 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_290
timestamp 1698431365
transform 1 0 33824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_292
timestamp 1698431365
transform 1 0 34048 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_346
timestamp 1698431365
transform 1 0 40096 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_350
timestamp 1698431365
transform 1 0 40544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_352
timestamp 1698431365
transform 1 0 40768 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_375
timestamp 1698431365
transform 1 0 43344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_377
timestamp 1698431365
transform 1 0 43568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_380
timestamp 1698431365
transform 1 0 43904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_392
timestamp 1698431365
transform 1 0 45248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_400
timestamp 1698431365
transform 1 0 46144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_402
timestamp 1698431365
transform 1 0 46368 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_419
timestamp 1698431365
transform 1 0 48272 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_502
timestamp 1698431365
transform 1 0 57568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_506
timestamp 1698431365
transform 1 0 58016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_508
timestamp 1698431365
transform 1 0 58240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_190
timestamp 1698431365
transform 1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_253
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_257
timestamp 1698431365
transform 1 0 30128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_265
timestamp 1698431365
transform 1 0 31024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_267
timestamp 1698431365
transform 1 0 31248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_288
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_296
timestamp 1698431365
transform 1 0 34496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_348
timestamp 1698431365
transform 1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_397
timestamp 1698431365
transform 1 0 45808 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_401
timestamp 1698431365
transform 1 0 46256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_415
timestamp 1698431365
transform 1 0 47824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698431365
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_431
timestamp 1698431365
transform 1 0 49616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_433
timestamp 1698431365
transform 1 0 49840 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_442
timestamp 1698431365
transform 1 0 50848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_460
timestamp 1698431365
transform 1 0 52864 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_476
timestamp 1698431365
transform 1 0 54656 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_484
timestamp 1698431365
transform 1 0 55552 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_488
timestamp 1698431365
transform 1 0 56000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_500
timestamp 1698431365
transform 1 0 57344 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_504
timestamp 1698431365
transform 1 0 57792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_506
timestamp 1698431365
transform 1 0 58016 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_127
timestamp 1698431365
transform 1 0 15568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_158
timestamp 1698431365
transform 1 0 19040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_162
timestamp 1698431365
transform 1 0 19488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_166
timestamp 1698431365
transform 1 0 19936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_198
timestamp 1698431365
transform 1 0 23520 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_202
timestamp 1698431365
transform 1 0 23968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_204
timestamp 1698431365
transform 1 0 24192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_211
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_215
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_256
timestamp 1698431365
transform 1 0 30016 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_272
timestamp 1698431365
transform 1 0 31808 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_281
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_285
timestamp 1698431365
transform 1 0 33264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_287
timestamp 1698431365
transform 1 0 33488 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_300
timestamp 1698431365
transform 1 0 34944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_308
timestamp 1698431365
transform 1 0 35840 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_327
timestamp 1698431365
transform 1 0 37968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_331
timestamp 1698431365
transform 1 0 38416 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_347
timestamp 1698431365
transform 1 0 40208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_355
timestamp 1698431365
transform 1 0 41104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_357
timestamp 1698431365
transform 1 0 41328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_360
timestamp 1698431365
transform 1 0 41664 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_376
timestamp 1698431365
transform 1 0 43456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_391
timestamp 1698431365
transform 1 0 45136 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_398
timestamp 1698431365
transform 1 0 45920 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_473
timestamp 1698431365
transform 1 0 54320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_477
timestamp 1698431365
transform 1 0 54768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_479
timestamp 1698431365
transform 1 0 54992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698431365
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698431365
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698431365
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_160
timestamp 1698431365
transform 1 0 19264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_193
timestamp 1698431365
transform 1 0 22960 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_232
timestamp 1698431365
transform 1 0 27328 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_286
timestamp 1698431365
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_356
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_392
timestamp 1698431365
transform 1 0 45248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_408
timestamp 1698431365
transform 1 0 47040 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_430
timestamp 1698431365
transform 1 0 49504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_438
timestamp 1698431365
transform 1 0 50400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_442
timestamp 1698431365
transform 1 0 50848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_444
timestamp 1698431365
transform 1 0 51072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_455
timestamp 1698431365
transform 1 0 52304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_459
timestamp 1698431365
transform 1 0 52752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_472
timestamp 1698431365
transform 1 0 54208 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_488
timestamp 1698431365
transform 1 0 56000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_500
timestamp 1698431365
transform 1 0 57344 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_503
timestamp 1698431365
transform 1 0 57680 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_166
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_189
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_196
timestamp 1698431365
transform 1 0 23296 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_228
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_255
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_259
timestamp 1698431365
transform 1 0 30352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_276
timestamp 1698431365
transform 1 0 32256 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_292
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_296
timestamp 1698431365
transform 1 0 34496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_298
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_323
timestamp 1698431365
transform 1 0 37520 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_353
timestamp 1698431365
transform 1 0 40880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_355
timestamp 1698431365
transform 1 0 41104 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_391
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_399
timestamp 1698431365
transform 1 0 46032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_403
timestamp 1698431365
transform 1 0 46480 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_414
timestamp 1698431365
transform 1 0 47712 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_430
timestamp 1698431365
transform 1 0 49504 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_434
timestamp 1698431365
transform 1 0 49952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_436
timestamp 1698431365
transform 1 0 50176 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_453
timestamp 1698431365
transform 1 0 52080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_469
timestamp 1698431365
transform 1 0 53872 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_471
timestamp 1698431365
transform 1 0 54096 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_501
timestamp 1698431365
transform 1 0 57456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_155
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_159
timestamp 1698431365
transform 1 0 19152 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_175
timestamp 1698431365
transform 1 0 20944 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_179
timestamp 1698431365
transform 1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_189
timestamp 1698431365
transform 1 0 22512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_249
timestamp 1698431365
transform 1 0 29232 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_265
timestamp 1698431365
transform 1 0 31024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_267
timestamp 1698431365
transform 1 0 31248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_270
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_300
timestamp 1698431365
transform 1 0 34944 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_330
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_334
timestamp 1698431365
transform 1 0 38752 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_338
timestamp 1698431365
transform 1 0 39200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_348
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_354
timestamp 1698431365
transform 1 0 40992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_371
timestamp 1698431365
transform 1 0 42896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_375
timestamp 1698431365
transform 1 0 43344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_387
timestamp 1698431365
transform 1 0 44688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_418
timestamp 1698431365
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_430
timestamp 1698431365
transform 1 0 49504 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_434
timestamp 1698431365
transform 1 0 49952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_436
timestamp 1698431365
transform 1 0 50176 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_450
timestamp 1698431365
transform 1 0 51744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_452
timestamp 1698431365
transform 1 0 51968 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_477
timestamp 1698431365
transform 1 0 54768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_483
timestamp 1698431365
transform 1 0 55440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_487
timestamp 1698431365
transform 1 0 55888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_489
timestamp 1698431365
transform 1 0 56112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698431365
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_113
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_143
timestamp 1698431365
transform 1 0 17360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_147
timestamp 1698431365
transform 1 0 17808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_149
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_158
timestamp 1698431365
transform 1 0 19040 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_193
timestamp 1698431365
transform 1 0 22960 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_197
timestamp 1698431365
transform 1 0 23408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_207
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_215
timestamp 1698431365
transform 1 0 25424 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_219
timestamp 1698431365
transform 1 0 25872 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_221
timestamp 1698431365
transform 1 0 26096 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_253
timestamp 1698431365
transform 1 0 29680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_262
timestamp 1698431365
transform 1 0 30688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_266
timestamp 1698431365
transform 1 0 31136 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_282
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_286
timestamp 1698431365
transform 1 0 33376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_302
timestamp 1698431365
transform 1 0 35168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_306
timestamp 1698431365
transform 1 0 35616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_341
timestamp 1698431365
transform 1 0 39536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_345
timestamp 1698431365
transform 1 0 39984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_353
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_357
timestamp 1698431365
transform 1 0 41328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_367
timestamp 1698431365
transform 1 0 42448 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_391
timestamp 1698431365
transform 1 0 45136 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_402
timestamp 1698431365
transform 1 0 46368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_406
timestamp 1698431365
transform 1 0 46816 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_436
timestamp 1698431365
transform 1 0 50176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_454
timestamp 1698431365
transform 1 0 52192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_461
timestamp 1698431365
transform 1 0 52976 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_493
timestamp 1698431365
transform 1 0 56560 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_148
timestamp 1698431365
transform 1 0 17920 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_159
timestamp 1698431365
transform 1 0 19152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_189
timestamp 1698431365
transform 1 0 22512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_222
timestamp 1698431365
transform 1 0 26208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_322
timestamp 1698431365
transform 1 0 37408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_324
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_327
timestamp 1698431365
transform 1 0 37968 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_389
timestamp 1698431365
transform 1 0 44912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_397
timestamp 1698431365
transform 1 0 45808 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_430
timestamp 1698431365
transform 1 0 49504 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_434
timestamp 1698431365
transform 1 0 49952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_438
timestamp 1698431365
transform 1 0 50400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_442
timestamp 1698431365
transform 1 0 50848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_446
timestamp 1698431365
transform 1 0 51296 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_478
timestamp 1698431365
transform 1 0 54880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_500
timestamp 1698431365
transform 1 0 57344 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_504
timestamp 1698431365
transform 1 0 57792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_506
timestamp 1698431365
transform 1 0 58016 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698431365
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_119
timestamp 1698431365
transform 1 0 14672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_159
timestamp 1698431365
transform 1 0 19152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_163
timestamp 1698431365
transform 1 0 19600 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_189
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_227
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_235
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_259
timestamp 1698431365
transform 1 0 30352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_289
timestamp 1698431365
transform 1 0 33712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_293
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698431365
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_349
timestamp 1698431365
transform 1 0 40432 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_357
timestamp 1698431365
transform 1 0 41328 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_360
timestamp 1698431365
transform 1 0 41664 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_376
timestamp 1698431365
transform 1 0 43456 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_403
timestamp 1698431365
transform 1 0 46480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_407
timestamp 1698431365
transform 1 0 46928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_411
timestamp 1698431365
transform 1 0 47376 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_443
timestamp 1698431365
transform 1 0 50960 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_473
timestamp 1698431365
transform 1 0 54320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_477
timestamp 1698431365
transform 1 0 54768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_479
timestamp 1698431365
transform 1 0 54992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_168
timestamp 1698431365
transform 1 0 20160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_176
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_249
timestamp 1698431365
transform 1 0 29232 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_265
timestamp 1698431365
transform 1 0 31024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698431365
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_286
timestamp 1698431365
transform 1 0 33376 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_321
timestamp 1698431365
transform 1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_323
timestamp 1698431365
transform 1 0 37520 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_326
timestamp 1698431365
transform 1 0 37856 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_340
timestamp 1698431365
transform 1 0 39424 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_354
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_363
timestamp 1698431365
transform 1 0 42000 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_379
timestamp 1698431365
transform 1 0 43792 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_387
timestamp 1698431365
transform 1 0 44688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_391
timestamp 1698431365
transform 1 0 45136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_395
timestamp 1698431365
transform 1 0 45584 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_399
timestamp 1698431365
transform 1 0 46032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_401
timestamp 1698431365
transform 1 0 46256 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_404
timestamp 1698431365
transform 1 0 46592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_413
timestamp 1698431365
transform 1 0 47600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_434
timestamp 1698431365
transform 1 0 49952 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_450
timestamp 1698431365
transform 1 0 51744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_452
timestamp 1698431365
transform 1 0 51968 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_482
timestamp 1698431365
transform 1 0 55328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_500
timestamp 1698431365
transform 1 0 57344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_193
timestamp 1698431365
transform 1 0 22960 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_197
timestamp 1698431365
transform 1 0 23408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_199
timestamp 1698431365
transform 1 0 23632 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_279
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_283
timestamp 1698431365
transform 1 0 33040 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_353
timestamp 1698431365
transform 1 0 40880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_391
timestamp 1698431365
transform 1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_403
timestamp 1698431365
transform 1 0 46480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_443
timestamp 1698431365
transform 1 0 50960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_447
timestamp 1698431365
transform 1 0 51408 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_473
timestamp 1698431365
transform 1 0 54320 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_482
timestamp 1698431365
transform 1 0 55328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_490
timestamp 1698431365
transform 1 0 56224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_507
timestamp 1698431365
transform 1 0 58128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1698431365
transform 1 0 13440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_162
timestamp 1698431365
transform 1 0 19488 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_165
timestamp 1698431365
transform 1 0 19824 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_181
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_195
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_216
timestamp 1698431365
transform 1 0 25536 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_232
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_265
timestamp 1698431365
transform 1 0 31024 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_294
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_326
timestamp 1698431365
transform 1 0 37856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_336
timestamp 1698431365
transform 1 0 38976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_340
timestamp 1698431365
transform 1 0 39424 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_356
timestamp 1698431365
transform 1 0 41216 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_370
timestamp 1698431365
transform 1 0 42784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_374
timestamp 1698431365
transform 1 0 43232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_384
timestamp 1698431365
transform 1 0 44352 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_438
timestamp 1698431365
transform 1 0 50400 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_468
timestamp 1698431365
transform 1 0 53760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_474
timestamp 1698431365
transform 1 0 54432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_478
timestamp 1698431365
transform 1 0 54880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_497
timestamp 1698431365
transform 1 0 57008 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_505
timestamp 1698431365
transform 1 0 57904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_135
timestamp 1698431365
transform 1 0 16464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_138
timestamp 1698431365
transform 1 0 16800 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_154
timestamp 1698431365
transform 1 0 18592 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_230
timestamp 1698431365
transform 1 0 27104 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_251
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_272
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_276
timestamp 1698431365
transform 1 0 32256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_284
timestamp 1698431365
transform 1 0 33152 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_292
timestamp 1698431365
transform 1 0 34048 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_300
timestamp 1698431365
transform 1 0 34944 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_304
timestamp 1698431365
transform 1 0 35392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_333
timestamp 1698431365
transform 1 0 38640 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_391
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_407
timestamp 1698431365
transform 1 0 46928 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_439
timestamp 1698431365
transform 1 0 50512 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_475
timestamp 1698431365
transform 1 0 54544 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_508
timestamp 1698431365
transform 1 0 58240 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_34
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_58
timestamp 1698431365
transform 1 0 7840 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_62
timestamp 1698431365
transform 1 0 8288 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_65
timestamp 1698431365
transform 1 0 8624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_106
timestamp 1698431365
transform 1 0 13216 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_110
timestamp 1698431365
transform 1 0 13664 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_121
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_125
timestamp 1698431365
transform 1 0 15344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_129
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_152
timestamp 1698431365
transform 1 0 18368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_156
timestamp 1698431365
transform 1 0 18816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_160
timestamp 1698431365
transform 1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_162
timestamp 1698431365
transform 1 0 19488 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_200
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_222
timestamp 1698431365
transform 1 0 26208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_226
timestamp 1698431365
transform 1 0 26656 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_237
timestamp 1698431365
transform 1 0 27888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_241
timestamp 1698431365
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_253
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_257
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_265
timestamp 1698431365
transform 1 0 31024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698431365
transform 1 0 32144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_296
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_300
timestamp 1698431365
transform 1 0 34944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_331
timestamp 1698431365
transform 1 0 38416 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_340
timestamp 1698431365
transform 1 0 39424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_348
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_358
timestamp 1698431365
transform 1 0 41440 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_379
timestamp 1698431365
transform 1 0 43792 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_383
timestamp 1698431365
transform 1 0 44240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_386
timestamp 1698431365
transform 1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_390
timestamp 1698431365
transform 1 0 45024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_394
timestamp 1698431365
transform 1 0 45472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_398
timestamp 1698431365
transform 1 0 45920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_402
timestamp 1698431365
transform 1 0 46368 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_426
timestamp 1698431365
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_462
timestamp 1698431365
transform 1 0 53088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_466
timestamp 1698431365
transform 1 0 53536 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_482
timestamp 1698431365
transform 1 0 55328 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_506
timestamp 1698431365
transform 1 0 58016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_53
timestamp 1698431365
transform 1 0 7280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_94
timestamp 1698431365
transform 1 0 11872 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_100
timestamp 1698431365
transform 1 0 12544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_121
timestamp 1698431365
transform 1 0 14896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_186
timestamp 1698431365
transform 1 0 22176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_190
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_194
timestamp 1698431365
transform 1 0 23072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_210
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_214
timestamp 1698431365
transform 1 0 25312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_256
timestamp 1698431365
transform 1 0 30016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_260
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_262
timestamp 1698431365
transform 1 0 30688 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_269
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_287
timestamp 1698431365
transform 1 0 33488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_295
timestamp 1698431365
transform 1 0 34384 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_302
timestamp 1698431365
transform 1 0 35168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_354
timestamp 1698431365
transform 1 0 40992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_356
timestamp 1698431365
transform 1 0 41216 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_365
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_369
timestamp 1698431365
transform 1 0 42672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_373
timestamp 1698431365
transform 1 0 43120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_375
timestamp 1698431365
transform 1 0 43344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_435
timestamp 1698431365
transform 1 0 50064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_439
timestamp 1698431365
transform 1 0 50512 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_470
timestamp 1698431365
transform 1 0 53984 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_486
timestamp 1698431365
transform 1 0 55776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_490
timestamp 1698431365
transform 1 0 56224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_496
timestamp 1698431365
transform 1 0 56896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_500
timestamp 1698431365
transform 1 0 57344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_26
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_30
timestamp 1698431365
transform 1 0 4704 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_88
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_132
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_161
timestamp 1698431365
transform 1 0 19376 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_177
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_185
timestamp 1698431365
transform 1 0 22064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_217
timestamp 1698431365
transform 1 0 25648 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_238
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_254
timestamp 1698431365
transform 1 0 29792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_261
timestamp 1698431365
transform 1 0 30576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1698431365
transform 1 0 31024 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698431365
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698431365
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_286
timestamp 1698431365
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_288
timestamp 1698431365
transform 1 0 33600 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_293
timestamp 1698431365
transform 1 0 34160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_297
timestamp 1698431365
transform 1 0 34608 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_313
timestamp 1698431365
transform 1 0 36400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_317
timestamp 1698431365
transform 1 0 36848 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_325
timestamp 1698431365
transform 1 0 37744 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_333
timestamp 1698431365
transform 1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_335
timestamp 1698431365
transform 1 0 38864 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_364
timestamp 1698431365
transform 1 0 42112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_395
timestamp 1698431365
transform 1 0 45584 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_403
timestamp 1698431365
transform 1 0 46480 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_407
timestamp 1698431365
transform 1 0 46928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_415
timestamp 1698431365
transform 1 0 47824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_454
timestamp 1698431365
transform 1 0 52192 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_460
timestamp 1698431365
transform 1 0 52864 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_476
timestamp 1698431365
transform 1 0 54656 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_484
timestamp 1698431365
transform 1 0 55552 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_488
timestamp 1698431365
transform 1 0 56000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_500
timestamp 1698431365
transform 1 0 57344 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_504
timestamp 1698431365
transform 1 0 57792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_506
timestamp 1698431365
transform 1 0 58016 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_88
timestamp 1698431365
transform 1 0 11200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_126
timestamp 1698431365
transform 1 0 15456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_130
timestamp 1698431365
transform 1 0 15904 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_146
timestamp 1698431365
transform 1 0 17696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_150
timestamp 1698431365
transform 1 0 18144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_152
timestamp 1698431365
transform 1 0 18368 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_155
timestamp 1698431365
transform 1 0 18704 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_193
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_201
timestamp 1698431365
transform 1 0 23856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_210
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_212
timestamp 1698431365
transform 1 0 25088 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_228
timestamp 1698431365
transform 1 0 26880 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_232
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_234
timestamp 1698431365
transform 1 0 27552 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_249
timestamp 1698431365
transform 1 0 29232 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_252
timestamp 1698431365
transform 1 0 29568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_256
timestamp 1698431365
transform 1 0 30016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_260
timestamp 1698431365
transform 1 0 30464 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_292
timestamp 1698431365
transform 1 0 34048 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_308
timestamp 1698431365
transform 1 0 35840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_331
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_335
timestamp 1698431365
transform 1 0 38864 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_343
timestamp 1698431365
transform 1 0 39760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_373
timestamp 1698431365
transform 1 0 43120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_377
timestamp 1698431365
transform 1 0 43568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_427
timestamp 1698431365
transform 1 0 49168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_443
timestamp 1698431365
transform 1 0 50960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_470
timestamp 1698431365
transform 1 0 53984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_478
timestamp 1698431365
transform 1 0 54880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_67
timestamp 1698431365
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_102
timestamp 1698431365
transform 1 0 12768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_114
timestamp 1698431365
transform 1 0 14112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_116
timestamp 1698431365
transform 1 0 14336 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_127
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_131
timestamp 1698431365
transform 1 0 16016 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_152
timestamp 1698431365
transform 1 0 18368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_156
timestamp 1698431365
transform 1 0 18816 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_160
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_190
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_194
timestamp 1698431365
transform 1 0 23072 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_238
timestamp 1698431365
transform 1 0 28000 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_242
timestamp 1698431365
transform 1 0 28448 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_249
timestamp 1698431365
transform 1 0 29232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_257
timestamp 1698431365
transform 1 0 30128 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_261
timestamp 1698431365
transform 1 0 30576 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_272
timestamp 1698431365
transform 1 0 31808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_294
timestamp 1698431365
transform 1 0 34272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_303
timestamp 1698431365
transform 1 0 35280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_305
timestamp 1698431365
transform 1 0 35504 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_308
timestamp 1698431365
transform 1 0 35840 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_324
timestamp 1698431365
transform 1 0 37632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_342
timestamp 1698431365
transform 1 0 39648 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_382
timestamp 1698431365
transform 1 0 44128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_386
timestamp 1698431365
transform 1 0 44576 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_418
timestamp 1698431365
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_438
timestamp 1698431365
transform 1 0 50400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_442
timestamp 1698431365
transform 1 0 50848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_444
timestamp 1698431365
transform 1 0 51072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_474
timestamp 1698431365
transform 1 0 54432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_478
timestamp 1698431365
transform 1 0 54880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_485
timestamp 1698431365
transform 1 0 55664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_489
timestamp 1698431365
transform 1 0 56112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_49
timestamp 1698431365
transform 1 0 6832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_78
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_127
timestamp 1698431365
transform 1 0 15568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_131
timestamp 1698431365
transform 1 0 16016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_135
timestamp 1698431365
transform 1 0 16464 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_153
timestamp 1698431365
transform 1 0 18480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_161
timestamp 1698431365
transform 1 0 19376 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_165
timestamp 1698431365
transform 1 0 19824 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_257
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_294
timestamp 1698431365
transform 1 0 34272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_360
timestamp 1698431365
transform 1 0 41664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_364
timestamp 1698431365
transform 1 0 42112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_368
timestamp 1698431365
transform 1 0 42560 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_379
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_391
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_423
timestamp 1698431365
transform 1 0 48720 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_427
timestamp 1698431365
transform 1 0 49168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_437
timestamp 1698431365
transform 1 0 50288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_441
timestamp 1698431365
transform 1 0 50736 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_449
timestamp 1698431365
transform 1 0 51632 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_453
timestamp 1698431365
transform 1 0 52080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_468
timestamp 1698431365
transform 1 0 53760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_470
timestamp 1698431365
transform 1 0 53984 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_497
timestamp 1698431365
transform 1 0 57008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_505
timestamp 1698431365
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_18
timestamp 1698431365
transform 1 0 3360 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_22
timestamp 1698431365
transform 1 0 3808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_24
timestamp 1698431365
transform 1 0 4032 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_54
timestamp 1698431365
transform 1 0 7392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_91
timestamp 1698431365
transform 1 0 11536 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_95
timestamp 1698431365
transform 1 0 11984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_173
timestamp 1698431365
transform 1 0 20720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_190
timestamp 1698431365
transform 1 0 22624 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_197
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_218
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_226
timestamp 1698431365
transform 1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_247
timestamp 1698431365
transform 1 0 29008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_251
timestamp 1698431365
transform 1 0 29456 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_255
timestamp 1698431365
transform 1 0 29904 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_259
timestamp 1698431365
transform 1 0 30352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_271
timestamp 1698431365
transform 1 0 31696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_275
timestamp 1698431365
transform 1 0 32144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_300
timestamp 1698431365
transform 1 0 34944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_312
timestamp 1698431365
transform 1 0 36288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_323
timestamp 1698431365
transform 1 0 37520 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_339
timestamp 1698431365
transform 1 0 39312 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_343
timestamp 1698431365
transform 1 0 39760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_415
timestamp 1698431365
transform 1 0 47824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_438
timestamp 1698431365
transform 1 0 50400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_450
timestamp 1698431365
transform 1 0 51744 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_458
timestamp 1698431365
transform 1 0 52640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_460
timestamp 1698431365
transform 1 0 52864 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_467
timestamp 1698431365
transform 1 0 53648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_471
timestamp 1698431365
transform 1 0 54096 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_487
timestamp 1698431365
transform 1 0 55888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_489
timestamp 1698431365
transform 1 0 56112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_499
timestamp 1698431365
transform 1 0 57232 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_505
timestamp 1698431365
transform 1 0 57904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_49
timestamp 1698431365
transform 1 0 6832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_64
timestamp 1698431365
transform 1 0 8512 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_98
timestamp 1698431365
transform 1 0 12320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_102
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_121
timestamp 1698431365
transform 1 0 14896 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_129
timestamp 1698431365
transform 1 0 15792 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_145
timestamp 1698431365
transform 1 0 17584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_149
timestamp 1698431365
transform 1 0 18032 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_165
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_189
timestamp 1698431365
transform 1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_201
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_213
timestamp 1698431365
transform 1 0 25200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_215
timestamp 1698431365
transform 1 0 25424 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_262
timestamp 1698431365
transform 1 0 30688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_264
timestamp 1698431365
transform 1 0 30912 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_346
timestamp 1698431365
transform 1 0 40096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_350
timestamp 1698431365
transform 1 0 40544 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_382
timestamp 1698431365
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_395
timestamp 1698431365
transform 1 0 45584 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_399
timestamp 1698431365
transform 1 0 46032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_440
timestamp 1698431365
transform 1 0 50624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_444
timestamp 1698431365
transform 1 0 51072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_452
timestamp 1698431365
transform 1 0 51968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_463
timestamp 1698431365
transform 1 0 53200 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_471
timestamp 1698431365
transform 1 0 54096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_473
timestamp 1698431365
transform 1 0 54320 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_34
timestamp 1698431365
transform 1 0 5152 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_50
timestamp 1698431365
transform 1 0 6944 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_99
timestamp 1698431365
transform 1 0 12432 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_107
timestamp 1698431365
transform 1 0 13328 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698431365
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_174
timestamp 1698431365
transform 1 0 20832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_176
timestamp 1698431365
transform 1 0 21056 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_199
timestamp 1698431365
transform 1 0 23632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_216
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_232
timestamp 1698431365
transform 1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_234
timestamp 1698431365
transform 1 0 27552 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_268
timestamp 1698431365
transform 1 0 31360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_294
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_298
timestamp 1698431365
transform 1 0 34720 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_330
timestamp 1698431365
transform 1 0 38304 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_360
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_393
timestamp 1698431365
transform 1 0 45360 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_397
timestamp 1698431365
transform 1 0 45808 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_413
timestamp 1698431365
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_424
timestamp 1698431365
transform 1 0 48832 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_427
timestamp 1698431365
transform 1 0 49168 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_431
timestamp 1698431365
transform 1 0 49616 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_438
timestamp 1698431365
transform 1 0 50400 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_470
timestamp 1698431365
transform 1 0 53984 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_484
timestamp 1698431365
transform 1 0 55552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_488
timestamp 1698431365
transform 1 0 56000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_500
timestamp 1698431365
transform 1 0 57344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_502
timestamp 1698431365
transform 1 0 57568 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_45
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_47
timestamp 1698431365
transform 1 0 6608 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_117
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_121
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_163
timestamp 1698431365
transform 1 0 19600 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_167
timestamp 1698431365
transform 1 0 20048 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_197
timestamp 1698431365
transform 1 0 23408 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_199
timestamp 1698431365
transform 1 0 23632 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_229
timestamp 1698431365
transform 1 0 26992 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_233
timestamp 1698431365
transform 1 0 27440 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_255
timestamp 1698431365
transform 1 0 29904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_259
timestamp 1698431365
transform 1 0 30352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_287
timestamp 1698431365
transform 1 0 33488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_331
timestamp 1698431365
transform 1 0 38416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_362
timestamp 1698431365
transform 1 0 41888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_366
timestamp 1698431365
transform 1 0 42336 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_374
timestamp 1698431365
transform 1 0 43232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_376
timestamp 1698431365
transform 1 0 43456 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_421
timestamp 1698431365
transform 1 0 48496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_425
timestamp 1698431365
transform 1 0 48944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_443
timestamp 1698431365
transform 1 0 50960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_473
timestamp 1698431365
transform 1 0 54320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_477
timestamp 1698431365
transform 1 0 54768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_479
timestamp 1698431365
transform 1 0 54992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_50
timestamp 1698431365
transform 1 0 6944 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_58
timestamp 1698431365
transform 1 0 7840 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_62
timestamp 1698431365
transform 1 0 8288 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_86
timestamp 1698431365
transform 1 0 10976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_127
timestamp 1698431365
transform 1 0 15568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_129
timestamp 1698431365
transform 1 0 15792 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_174
timestamp 1698431365
transform 1 0 20832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_178
timestamp 1698431365
transform 1 0 21280 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_194
timestamp 1698431365
transform 1 0 23072 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_228
timestamp 1698431365
transform 1 0 26880 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_236
timestamp 1698431365
transform 1 0 27776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_240
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_242
timestamp 1698431365
transform 1 0 28448 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_245
timestamp 1698431365
transform 1 0 28784 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_261
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_265
timestamp 1698431365
transform 1 0 31024 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_344
timestamp 1698431365
transform 1 0 39872 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_372
timestamp 1698431365
transform 1 0 43008 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_387
timestamp 1698431365
transform 1 0 44688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_391
timestamp 1698431365
transform 1 0 45136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_399
timestamp 1698431365
transform 1 0 46032 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_413
timestamp 1698431365
transform 1 0 47600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_417
timestamp 1698431365
transform 1 0 48048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_432
timestamp 1698431365
transform 1 0 49728 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_444
timestamp 1698431365
transform 1 0 51072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_446
timestamp 1698431365
transform 1 0 51296 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_449
timestamp 1698431365
transform 1 0 51632 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_455
timestamp 1698431365
transform 1 0 52304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_465
timestamp 1698431365
transform 1 0 53424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_472
timestamp 1698431365
transform 1 0 54208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_482
timestamp 1698431365
transform 1 0 55328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_500
timestamp 1698431365
transform 1 0 57344 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_504
timestamp 1698431365
transform 1 0 57792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_506
timestamp 1698431365
transform 1 0 58016 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_69
timestamp 1698431365
transform 1 0 9072 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_77
timestamp 1698431365
transform 1 0 9968 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_81
timestamp 1698431365
transform 1 0 10416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_83
timestamp 1698431365
transform 1 0 10640 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_109
timestamp 1698431365
transform 1 0 13552 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_127
timestamp 1698431365
transform 1 0 15568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_173
timestamp 1698431365
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_206
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_210
timestamp 1698431365
transform 1 0 24864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_220
timestamp 1698431365
transform 1 0 25984 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_228
timestamp 1698431365
transform 1 0 26880 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_232
timestamp 1698431365
transform 1 0 27328 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_253
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_261
timestamp 1698431365
transform 1 0 30576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_309
timestamp 1698431365
transform 1 0 35952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_367
timestamp 1698431365
transform 1 0 42448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_375
timestamp 1698431365
transform 1 0 43344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_403
timestamp 1698431365
transform 1 0 46480 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_411
timestamp 1698431365
transform 1 0 47376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_415
timestamp 1698431365
transform 1 0 47824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_417
timestamp 1698431365
transform 1 0 48048 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_486
timestamp 1698431365
transform 1 0 55776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_490
timestamp 1698431365
transform 1 0 56224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_494
timestamp 1698431365
transform 1 0 56672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_505
timestamp 1698431365
transform 1 0 57904 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_34
timestamp 1698431365
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_50
timestamp 1698431365
transform 1 0 6944 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_54
timestamp 1698431365
transform 1 0 7392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_61
timestamp 1698431365
transform 1 0 8176 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_91
timestamp 1698431365
transform 1 0 11536 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_107
timestamp 1698431365
transform 1 0 13328 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_134
timestamp 1698431365
transform 1 0 16352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_176
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_180
timestamp 1698431365
transform 1 0 21504 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_204
timestamp 1698431365
transform 1 0 24192 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_251
timestamp 1698431365
transform 1 0 29456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_253
timestamp 1698431365
transform 1 0 29680 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_278
timestamp 1698431365
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_368
timestamp 1698431365
transform 1 0 42560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_376
timestamp 1698431365
transform 1 0 43456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_387
timestamp 1698431365
transform 1 0 44688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_391
timestamp 1698431365
transform 1 0 45136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_393
timestamp 1698431365
transform 1 0 45360 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_412
timestamp 1698431365
transform 1 0 47488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_454
timestamp 1698431365
transform 1 0 52192 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_470
timestamp 1698431365
transform 1 0 53984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_474
timestamp 1698431365
transform 1 0 54432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_481
timestamp 1698431365
transform 1 0 55216 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_489
timestamp 1698431365
transform 1 0 56112 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_501
timestamp 1698431365
transform 1 0 57456 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_6
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_22
timestamp 1698431365
transform 1 0 3808 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_30
timestamp 1698431365
transform 1 0 4704 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_49
timestamp 1698431365
transform 1 0 6832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_63
timestamp 1698431365
transform 1 0 8400 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_71
timestamp 1698431365
transform 1 0 9296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_73
timestamp 1698431365
transform 1 0 9520 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_89
timestamp 1698431365
transform 1 0 11312 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_97
timestamp 1698431365
transform 1 0 12208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_149
timestamp 1698431365
transform 1 0 18032 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_157
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_169
timestamp 1698431365
transform 1 0 20272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_206
timestamp 1698431365
transform 1 0 24416 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_222
timestamp 1698431365
transform 1 0 26208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_230
timestamp 1698431365
transform 1 0 27104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_232
timestamp 1698431365
transform 1 0 27328 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_330
timestamp 1698431365
transform 1 0 38304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_334
timestamp 1698431365
transform 1 0 38752 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_340
timestamp 1698431365
transform 1 0 39424 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_348
timestamp 1698431365
transform 1 0 40320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_354
timestamp 1698431365
transform 1 0 40992 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_370
timestamp 1698431365
transform 1 0 42784 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_374
timestamp 1698431365
transform 1 0 43232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_392
timestamp 1698431365
transform 1 0 45248 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_396
timestamp 1698431365
transform 1 0 45696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_427
timestamp 1698431365
transform 1 0 49168 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_432
timestamp 1698431365
transform 1 0 49728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_436
timestamp 1698431365
transform 1 0 50176 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_452
timestamp 1698431365
transform 1 0 51968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_454
timestamp 1698431365
transform 1 0 52192 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_467
timestamp 1698431365
transform 1 0 53648 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_488
timestamp 1698431365
transform 1 0 56000 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_499
timestamp 1698431365
transform 1 0 57232 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_507
timestamp 1698431365
transform 1 0 58128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_10
timestamp 1698431365
transform 1 0 2464 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_42
timestamp 1698431365
transform 1 0 6048 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_58
timestamp 1698431365
transform 1 0 7840 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_82
timestamp 1698431365
transform 1 0 10528 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_86
timestamp 1698431365
transform 1 0 10976 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_88
timestamp 1698431365
transform 1 0 11200 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_104
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_106
timestamp 1698431365
transform 1 0 13216 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_115
timestamp 1698431365
transform 1 0 14224 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_134
timestamp 1698431365
transform 1 0 16352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_146
timestamp 1698431365
transform 1 0 17696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_148
timestamp 1698431365
transform 1 0 17920 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_189
timestamp 1698431365
transform 1 0 22512 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_198
timestamp 1698431365
transform 1 0 23520 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_234
timestamp 1698431365
transform 1 0 27552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_238
timestamp 1698431365
transform 1 0 28000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_240
timestamp 1698431365
transform 1 0 28224 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_243
timestamp 1698431365
transform 1 0 28560 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_272
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_274
timestamp 1698431365
transform 1 0 32032 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_284
timestamp 1698431365
transform 1 0 33152 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_339
timestamp 1698431365
transform 1 0 39312 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_347
timestamp 1698431365
transform 1 0 40208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_397
timestamp 1698431365
transform 1 0 45808 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_413
timestamp 1698431365
transform 1 0 47600 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_417
timestamp 1698431365
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_430
timestamp 1698431365
transform 1 0 49504 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_434
timestamp 1698431365
transform 1 0 49952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_442
timestamp 1698431365
transform 1 0 50848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_446
timestamp 1698431365
transform 1 0 51296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_448
timestamp 1698431365
transform 1 0 51520 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_455
timestamp 1698431365
transform 1 0 52304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_467
timestamp 1698431365
transform 1 0 53648 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_475
timestamp 1698431365
transform 1 0 54544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_477
timestamp 1698431365
transform 1 0 54768 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_506
timestamp 1698431365
transform 1 0 58016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_61
timestamp 1698431365
transform 1 0 8176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_63
timestamp 1698431365
transform 1 0 8400 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_77
timestamp 1698431365
transform 1 0 9968 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_81
timestamp 1698431365
transform 1 0 10416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_83
timestamp 1698431365
transform 1 0 10640 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_112
timestamp 1698431365
transform 1 0 13888 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_120
timestamp 1698431365
transform 1 0 14784 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_124
timestamp 1698431365
transform 1 0 15232 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_135
timestamp 1698431365
transform 1 0 16464 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698431365
transform 1 0 19824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_183
timestamp 1698431365
transform 1 0 21840 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_187
timestamp 1698431365
transform 1 0 22288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_196
timestamp 1698431365
transform 1 0 23296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_210
timestamp 1698431365
transform 1 0 24864 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_218
timestamp 1698431365
transform 1 0 25760 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_222
timestamp 1698431365
transform 1 0 26208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_224
timestamp 1698431365
transform 1 0 26432 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_259
timestamp 1698431365
transform 1 0 30352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_294
timestamp 1698431365
transform 1 0 34272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_296
timestamp 1698431365
transform 1 0 34496 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_312
timestamp 1698431365
transform 1 0 36288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_328
timestamp 1698431365
transform 1 0 38080 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_344
timestamp 1698431365
transform 1 0 39872 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_358
timestamp 1698431365
transform 1 0 41440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_362
timestamp 1698431365
transform 1 0 41888 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_370
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_374
timestamp 1698431365
transform 1 0 43232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_376
timestamp 1698431365
transform 1 0 43456 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_383
timestamp 1698431365
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_419
timestamp 1698431365
transform 1 0 48272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_423
timestamp 1698431365
transform 1 0 48720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_425
timestamp 1698431365
transform 1 0 48944 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_461
timestamp 1698431365
transform 1 0 52976 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_491
timestamp 1698431365
transform 1 0 56336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_495
timestamp 1698431365
transform 1 0 56784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_503
timestamp 1698431365
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_507
timestamp 1698431365
transform 1 0 58128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_56
timestamp 1698431365
transform 1 0 7616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_91
timestamp 1698431365
transform 1 0 11536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_106
timestamp 1698431365
transform 1 0 13216 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_146
timestamp 1698431365
transform 1 0 17696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_183
timestamp 1698431365
transform 1 0 21840 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_256
timestamp 1698431365
transform 1 0 30016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_260
timestamp 1698431365
transform 1 0 30464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_269
timestamp 1698431365
transform 1 0 31472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698431365
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_330
timestamp 1698431365
transform 1 0 38304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_345
timestamp 1698431365
transform 1 0 39984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_381
timestamp 1698431365
transform 1 0 44016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_385
timestamp 1698431365
transform 1 0 44464 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_407
timestamp 1698431365
transform 1 0 46928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_415
timestamp 1698431365
transform 1 0 47824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_419
timestamp 1698431365
transform 1 0 48272 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_18
timestamp 1698431365
transform 1 0 3360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_20
timestamp 1698431365
transform 1 0 3584 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_26
timestamp 1698431365
transform 1 0 4256 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_30
timestamp 1698431365
transform 1 0 4704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_55
timestamp 1698431365
transform 1 0 7504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_59
timestamp 1698431365
transform 1 0 7952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_78
timestamp 1698431365
transform 1 0 10080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_80
timestamp 1698431365
transform 1 0 10304 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_123
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_196
timestamp 1698431365
transform 1 0 23296 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_200
timestamp 1698431365
transform 1 0 23744 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_209
timestamp 1698431365
transform 1 0 24752 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_217
timestamp 1698431365
transform 1 0 25648 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_252
timestamp 1698431365
transform 1 0 29568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_256
timestamp 1698431365
transform 1 0 30016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_331
timestamp 1698431365
transform 1 0 38416 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_355
timestamp 1698431365
transform 1 0 41104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_357
timestamp 1698431365
transform 1 0 41328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_366
timestamp 1698431365
transform 1 0 42336 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_430
timestamp 1698431365
transform 1 0 49504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_434
timestamp 1698431365
transform 1 0 49952 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_450
timestamp 1698431365
transform 1 0 51744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_454
timestamp 1698431365
transform 1 0 52192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_465
timestamp 1698431365
transform 1 0 53424 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_468
timestamp 1698431365
transform 1 0 53760 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_476
timestamp 1698431365
transform 1 0 54656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_34
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_38
timestamp 1698431365
transform 1 0 5600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_40
timestamp 1698431365
transform 1 0 5824 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_62
timestamp 1698431365
transform 1 0 8288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_84
timestamp 1698431365
transform 1 0 10752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_93
timestamp 1698431365
transform 1 0 11760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_108
timestamp 1698431365
transform 1 0 13440 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_116
timestamp 1698431365
transform 1 0 14336 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_120
timestamp 1698431365
transform 1 0 14784 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_159
timestamp 1698431365
transform 1 0 19152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_187
timestamp 1698431365
transform 1 0 22288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_191
timestamp 1698431365
transform 1 0 22736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_240
timestamp 1698431365
transform 1 0 28224 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_248
timestamp 1698431365
transform 1 0 29120 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_252
timestamp 1698431365
transform 1 0 29568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_286
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_303
timestamp 1698431365
transform 1 0 35280 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_319
timestamp 1698431365
transform 1 0 37072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_321
timestamp 1698431365
transform 1 0 37296 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_328
timestamp 1698431365
transform 1 0 38080 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_332
timestamp 1698431365
transform 1 0 38528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_334
timestamp 1698431365
transform 1 0 38752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_384
timestamp 1698431365
transform 1 0 44352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_390
timestamp 1698431365
transform 1 0 45024 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_394
timestamp 1698431365
transform 1 0 45472 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_396
timestamp 1698431365
transform 1 0 45696 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_405
timestamp 1698431365
transform 1 0 46704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_413
timestamp 1698431365
transform 1 0 47600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_417
timestamp 1698431365
transform 1 0 48048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_419
timestamp 1698431365
transform 1 0 48272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_431
timestamp 1698431365
transform 1 0 49616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_464
timestamp 1698431365
transform 1 0 53312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_474
timestamp 1698431365
transform 1 0 54432 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_496
timestamp 1698431365
transform 1 0 56896 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_500
timestamp 1698431365
transform 1 0 57344 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_6
timestamp 1698431365
transform 1 0 2016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_8
timestamp 1698431365
transform 1 0 2240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_43
timestamp 1698431365
transform 1 0 6160 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_47
timestamp 1698431365
transform 1 0 6608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_51
timestamp 1698431365
transform 1 0 7056 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_83
timestamp 1698431365
transform 1 0 10640 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_87
timestamp 1698431365
transform 1 0 11088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_113
timestamp 1698431365
transform 1 0 14000 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_173
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_183
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_240
timestamp 1698431365
transform 1 0 28224 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_285
timestamp 1698431365
transform 1 0 33264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_293
timestamp 1698431365
transform 1 0 34160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_295
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_304
timestamp 1698431365
transform 1 0 35392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1698431365
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_349
timestamp 1698431365
transform 1 0 40432 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_357
timestamp 1698431365
transform 1 0 41328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_367
timestamp 1698431365
transform 1 0 42448 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_371
timestamp 1698431365
transform 1 0 42896 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_400
timestamp 1698431365
transform 1 0 46144 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_408
timestamp 1698431365
transform 1 0 47040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_414
timestamp 1698431365
transform 1 0 47712 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_422
timestamp 1698431365
transform 1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_430
timestamp 1698431365
transform 1 0 49504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_434
timestamp 1698431365
transform 1 0 49952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_438
timestamp 1698431365
transform 1 0 50400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_448
timestamp 1698431365
transform 1 0 51520 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_452
timestamp 1698431365
transform 1 0 51968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698431365
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_506
timestamp 1698431365
transform 1 0 58016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_508
timestamp 1698431365
transform 1 0 58240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_31
timestamp 1698431365
transform 1 0 4816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_35
timestamp 1698431365
transform 1 0 5264 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_39
timestamp 1698431365
transform 1 0 5712 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_41
timestamp 1698431365
transform 1 0 5936 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_48
timestamp 1698431365
transform 1 0 6720 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_62
timestamp 1698431365
transform 1 0 8288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_88
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_96
timestamp 1698431365
transform 1 0 12096 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_102
timestamp 1698431365
transform 1 0 12768 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_181
timestamp 1698431365
transform 1 0 21616 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_185
timestamp 1698431365
transform 1 0 22064 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698431365
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_224
timestamp 1698431365
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_336
timestamp 1698431365
transform 1 0 38976 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_344
timestamp 1698431365
transform 1 0 39872 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_368
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_372
timestamp 1698431365
transform 1 0 43008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_374
timestamp 1698431365
transform 1 0 43232 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698431365
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_430
timestamp 1698431365
transform 1 0 49504 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_438
timestamp 1698431365
transform 1 0 50400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_454
timestamp 1698431365
transform 1 0 52192 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_470
timestamp 1698431365
transform 1 0 53984 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_478
timestamp 1698431365
transform 1 0 54880 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_482
timestamp 1698431365
transform 1 0 55328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_484
timestamp 1698431365
transform 1 0 55552 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_505
timestamp 1698431365
transform 1 0 57904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_10
timestamp 1698431365
transform 1 0 2464 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_17
timestamp 1698431365
transform 1 0 3248 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_19
timestamp 1698431365
transform 1 0 3472 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_42
timestamp 1698431365
transform 1 0 6048 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_81
timestamp 1698431365
transform 1 0 10416 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_103
timestamp 1698431365
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_185
timestamp 1698431365
transform 1 0 22064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_189
timestamp 1698431365
transform 1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_191
timestamp 1698431365
transform 1 0 22736 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_202
timestamp 1698431365
transform 1 0 23968 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_220
timestamp 1698431365
transform 1 0 25984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_239
timestamp 1698431365
transform 1 0 28112 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_243
timestamp 1698431365
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_252
timestamp 1698431365
transform 1 0 29568 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_268
timestamp 1698431365
transform 1 0 31360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698431365
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_329
timestamp 1698431365
transform 1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_333
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_341
timestamp 1698431365
transform 1 0 39536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_374
timestamp 1698431365
transform 1 0 43232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_378
timestamp 1698431365
transform 1 0 43680 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_389
timestamp 1698431365
transform 1 0 44912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_396
timestamp 1698431365
transform 1 0 45696 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_428
timestamp 1698431365
transform 1 0 49280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_442
timestamp 1698431365
transform 1 0 50848 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_446
timestamp 1698431365
transform 1 0 51296 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_467
timestamp 1698431365
transform 1 0 53648 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_475
timestamp 1698431365
transform 1 0 54544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_10
timestamp 1698431365
transform 1 0 2464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_14
timestamp 1698431365
transform 1 0 2912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_16
timestamp 1698431365
transform 1 0 3136 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_19
timestamp 1698431365
transform 1 0 3472 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_27
timestamp 1698431365
transform 1 0 4368 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_31
timestamp 1698431365
transform 1 0 4816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_33
timestamp 1698431365
transform 1 0 5040 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_63
timestamp 1698431365
transform 1 0 8400 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_77
timestamp 1698431365
transform 1 0 9968 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_81
timestamp 1698431365
transform 1 0 10416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_83
timestamp 1698431365
transform 1 0 10640 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_113
timestamp 1698431365
transform 1 0 14000 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_186
timestamp 1698431365
transform 1 0 22176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_190
timestamp 1698431365
transform 1 0 22624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_194
timestamp 1698431365
transform 1 0 23072 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_196
timestamp 1698431365
transform 1 0 23296 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_202
timestamp 1698431365
transform 1 0 23968 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_261
timestamp 1698431365
transform 1 0 30576 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_284
timestamp 1698431365
transform 1 0 33152 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_310
timestamp 1698431365
transform 1 0 36064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_343
timestamp 1698431365
transform 1 0 39760 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_347
timestamp 1698431365
transform 1 0 40208 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_362
timestamp 1698431365
transform 1 0 41888 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_366
timestamp 1698431365
transform 1 0 42336 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_374
timestamp 1698431365
transform 1 0 43232 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_381
timestamp 1698431365
transform 1 0 44016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_387
timestamp 1698431365
transform 1 0 44688 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_424
timestamp 1698431365
transform 1 0 48832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_454
timestamp 1698431365
transform 1 0 52192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_458
timestamp 1698431365
transform 1 0 52640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_489
timestamp 1698431365
transform 1 0 56112 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_504
timestamp 1698431365
transform 1 0 57792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_506
timestamp 1698431365
transform 1 0 58016 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_10
timestamp 1698431365
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_12
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_25
timestamp 1698431365
transform 1 0 4144 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_53
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_61
timestamp 1698431365
transform 1 0 8176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_71
timestamp 1698431365
transform 1 0 9296 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_87
timestamp 1698431365
transform 1 0 11088 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_95
timestamp 1698431365
transform 1 0 11984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_109
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_116
timestamp 1698431365
transform 1 0 14336 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_124
timestamp 1698431365
transform 1 0 15232 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_183
timestamp 1698431365
transform 1 0 21840 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_187
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_203
timestamp 1698431365
transform 1 0 24080 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_207
timestamp 1698431365
transform 1 0 24528 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_225
timestamp 1698431365
transform 1 0 26544 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_237
timestamp 1698431365
transform 1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_239
timestamp 1698431365
transform 1 0 28112 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_269
timestamp 1698431365
transform 1 0 31472 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_277
timestamp 1698431365
transform 1 0 32368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_281
timestamp 1698431365
transform 1 0 32816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_285
timestamp 1698431365
transform 1 0 33264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_289
timestamp 1698431365
transform 1 0 33712 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_293
timestamp 1698431365
transform 1 0 34160 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_309
timestamp 1698431365
transform 1 0 35952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_335
timestamp 1698431365
transform 1 0 38864 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_355
timestamp 1698431365
transform 1 0 41104 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_398
timestamp 1698431365
transform 1 0 45920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_408
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_424
timestamp 1698431365
transform 1 0 48832 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_428
timestamp 1698431365
transform 1 0 49280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_430
timestamp 1698431365
transform 1 0 49504 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_438
timestamp 1698431365
transform 1 0 50400 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_446
timestamp 1698431365
transform 1 0 51296 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_461
timestamp 1698431365
transform 1 0 52976 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_35
timestamp 1698431365
transform 1 0 5264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_39
timestamp 1698431365
transform 1 0 5712 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_55
timestamp 1698431365
transform 1 0 7504 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_63
timestamp 1698431365
transform 1 0 8400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_67
timestamp 1698431365
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_104
timestamp 1698431365
transform 1 0 12992 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_108
timestamp 1698431365
transform 1 0 13440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_193
timestamp 1698431365
transform 1 0 22960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_197
timestamp 1698431365
transform 1 0 23408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_205
timestamp 1698431365
transform 1 0 24304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_244
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_260
timestamp 1698431365
transform 1 0 30464 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_268
timestamp 1698431365
transform 1 0 31360 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_270
timestamp 1698431365
transform 1 0 31584 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_382
timestamp 1698431365
transform 1 0 44128 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_386
timestamp 1698431365
transform 1 0 44576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_388
timestamp 1698431365
transform 1 0 44800 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_454
timestamp 1698431365
transform 1 0 52192 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_458
timestamp 1698431365
transform 1 0 52640 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_487
timestamp 1698431365
transform 1 0 55888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_502
timestamp 1698431365
transform 1 0 57568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_506
timestamp 1698431365
transform 1 0 58016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_6
timestamp 1698431365
transform 1 0 2016 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_8
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_15
timestamp 1698431365
transform 1 0 3024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_45
timestamp 1698431365
transform 1 0 6384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_49
timestamp 1698431365
transform 1 0 6832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_71
timestamp 1698431365
transform 1 0 9296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_75
timestamp 1698431365
transform 1 0 9744 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_91
timestamp 1698431365
transform 1 0 11536 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_99
timestamp 1698431365
transform 1 0 12432 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_103
timestamp 1698431365
transform 1 0 12880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_113
timestamp 1698431365
transform 1 0 14000 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_121
timestamp 1698431365
transform 1 0 14896 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_142
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_146
timestamp 1698431365
transform 1 0 17696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_148
timestamp 1698431365
transform 1 0 17920 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_197
timestamp 1698431365
transform 1 0 23408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_201
timestamp 1698431365
transform 1 0 23856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_211
timestamp 1698431365
transform 1 0 24976 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_221
timestamp 1698431365
transform 1 0 26096 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_237
timestamp 1698431365
transform 1 0 27888 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_263
timestamp 1698431365
transform 1 0 30800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_285
timestamp 1698431365
transform 1 0 33264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_287
timestamp 1698431365
transform 1 0 33488 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_304
timestamp 1698431365
transform 1 0 35392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_308
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_327
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_343
timestamp 1698431365
transform 1 0 39760 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_347
timestamp 1698431365
transform 1 0 40208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_349
timestamp 1698431365
transform 1 0 40432 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_410
timestamp 1698431365
transform 1 0 47264 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_465
timestamp 1698431365
transform 1 0 53424 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_469
timestamp 1698431365
transform 1 0 53872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_485
timestamp 1698431365
transform 1 0 55664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_487
timestamp 1698431365
transform 1 0 55888 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_498
timestamp 1698431365
transform 1 0 57120 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_504
timestamp 1698431365
transform 1 0 57792 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_506
timestamp 1698431365
transform 1 0 58016 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_10
timestamp 1698431365
transform 1 0 2464 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_14
timestamp 1698431365
transform 1 0 2912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_17
timestamp 1698431365
transform 1 0 3248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_25
timestamp 1698431365
transform 1 0 4144 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_29
timestamp 1698431365
transform 1 0 4592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_35
timestamp 1698431365
transform 1 0 5264 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_39
timestamp 1698431365
transform 1 0 5712 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_69
timestamp 1698431365
transform 1 0 9072 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_80
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_96
timestamp 1698431365
transform 1 0 12096 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_98
timestamp 1698431365
transform 1 0 12320 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_101
timestamp 1698431365
transform 1 0 12656 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_109
timestamp 1698431365
transform 1 0 13552 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_113
timestamp 1698431365
transform 1 0 14000 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_131
timestamp 1698431365
transform 1 0 16016 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_139
timestamp 1698431365
transform 1 0 16912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_156
timestamp 1698431365
transform 1 0 18816 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_172
timestamp 1698431365
transform 1 0 20608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_174
timestamp 1698431365
transform 1 0 20832 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_177
timestamp 1698431365
transform 1 0 21168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_179
timestamp 1698431365
transform 1 0 21392 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_201
timestamp 1698431365
transform 1 0 23856 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_230
timestamp 1698431365
transform 1 0 27104 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_238
timestamp 1698431365
transform 1 0 28000 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_246
timestamp 1698431365
transform 1 0 28896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_250
timestamp 1698431365
transform 1 0 29344 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_266
timestamp 1698431365
transform 1 0 31136 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_313
timestamp 1698431365
transform 1 0 36400 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_317
timestamp 1698431365
transform 1 0 36848 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_325
timestamp 1698431365
transform 1 0 37744 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_329
timestamp 1698431365
transform 1 0 38192 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_332
timestamp 1698431365
transform 1 0 38528 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_348
timestamp 1698431365
transform 1 0 40320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_368
timestamp 1698431365
transform 1 0 42560 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_376
timestamp 1698431365
transform 1 0 43456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_378
timestamp 1698431365
transform 1 0 43680 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_381
timestamp 1698431365
transform 1 0 44016 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_413
timestamp 1698431365
transform 1 0 47600 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_417
timestamp 1698431365
transform 1 0 48048 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_428
timestamp 1698431365
transform 1 0 49280 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_432
timestamp 1698431365
transform 1 0 49728 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_462
timestamp 1698431365
transform 1 0 53088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_466
timestamp 1698431365
transform 1 0 53536 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_474
timestamp 1698431365
transform 1 0 54432 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_478
timestamp 1698431365
transform 1 0 54880 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_500
timestamp 1698431365
transform 1 0 57344 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_53
timestamp 1698431365
transform 1 0 7280 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_57
timestamp 1698431365
transform 1 0 7728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_67
timestamp 1698431365
transform 1 0 8848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_111
timestamp 1698431365
transform 1 0 13776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_115
timestamp 1698431365
transform 1 0 14224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_130
timestamp 1698431365
transform 1 0 15904 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_155
timestamp 1698431365
transform 1 0 18704 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_163
timestamp 1698431365
transform 1 0 19600 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_181
timestamp 1698431365
transform 1 0 21616 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_189
timestamp 1698431365
transform 1 0 22512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_195
timestamp 1698431365
transform 1 0 23184 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_227
timestamp 1698431365
transform 1 0 26768 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_262
timestamp 1698431365
transform 1 0 30688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_293
timestamp 1698431365
transform 1 0 34160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_297
timestamp 1698431365
transform 1 0 34608 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1698431365
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_321
timestamp 1698431365
transform 1 0 37296 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_330
timestamp 1698431365
transform 1 0 38304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_332
timestamp 1698431365
transform 1 0 38528 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_362
timestamp 1698431365
transform 1 0 41888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_366
timestamp 1698431365
transform 1 0 42336 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_382
timestamp 1698431365
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_396
timestamp 1698431365
transform 1 0 45696 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_400
timestamp 1698431365
transform 1 0 46144 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_422
timestamp 1698431365
transform 1 0 48608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_432
timestamp 1698431365
transform 1 0 49728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_436
timestamp 1698431365
transform 1 0 50176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_438
timestamp 1698431365
transform 1 0 50400 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_447
timestamp 1698431365
transform 1 0 51408 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_473
timestamp 1698431365
transform 1 0 54320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_477
timestamp 1698431365
transform 1 0 54768 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_6
timestamp 1698431365
transform 1 0 2016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_14
timestamp 1698431365
transform 1 0 2912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_41
timestamp 1698431365
transform 1 0 5936 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_57
timestamp 1698431365
transform 1 0 7728 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_105
timestamp 1698431365
transform 1 0 13104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_133
timestamp 1698431365
transform 1 0 16240 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_137
timestamp 1698431365
transform 1 0 16688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_167
timestamp 1698431365
transform 1 0 20048 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_183
timestamp 1698431365
transform 1 0 21840 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_191
timestamp 1698431365
transform 1 0 22736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_195
timestamp 1698431365
transform 1 0 23184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_216
timestamp 1698431365
transform 1 0 25536 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_236
timestamp 1698431365
transform 1 0 27776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_240
timestamp 1698431365
transform 1 0 28224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_276
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_294
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_296
timestamp 1698431365
transform 1 0 34496 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_305
timestamp 1698431365
transform 1 0 35504 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_358
timestamp 1698431365
transform 1 0 41440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_362
timestamp 1698431365
transform 1 0 41888 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_378
timestamp 1698431365
transform 1 0 43680 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_382
timestamp 1698431365
transform 1 0 44128 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_403
timestamp 1698431365
transform 1 0 46480 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_411
timestamp 1698431365
transform 1 0 47376 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_446
timestamp 1698431365
transform 1 0 51296 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_454
timestamp 1698431365
transform 1 0 52192 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_458
timestamp 1698431365
transform 1 0 52640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_460
timestamp 1698431365
transform 1 0 52864 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_469
timestamp 1698431365
transform 1 0 53872 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_483
timestamp 1698431365
transform 1 0 55440 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_487
timestamp 1698431365
transform 1 0 55888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_489
timestamp 1698431365
transform 1 0 56112 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_43
timestamp 1698431365
transform 1 0 6160 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_75
timestamp 1698431365
transform 1 0 9744 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_98
timestamp 1698431365
transform 1 0 12320 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_120
timestamp 1698431365
transform 1 0 14784 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_124
timestamp 1698431365
transform 1 0 15232 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_139
timestamp 1698431365
transform 1 0 16912 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_163
timestamp 1698431365
transform 1 0 19600 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_185
timestamp 1698431365
transform 1 0 22064 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_212
timestamp 1698431365
transform 1 0 25088 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_255
timestamp 1698431365
transform 1 0 29904 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_287
timestamp 1698431365
transform 1 0 33488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_291
timestamp 1698431365
transform 1 0 33936 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_293
timestamp 1698431365
transform 1 0 34160 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_307
timestamp 1698431365
transform 1 0 35728 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_343
timestamp 1698431365
transform 1 0 39760 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_351
timestamp 1698431365
transform 1 0 40656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_376
timestamp 1698431365
transform 1 0 43456 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_380
timestamp 1698431365
transform 1 0 43904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_382
timestamp 1698431365
transform 1 0 44128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_416
timestamp 1698431365
transform 1 0 47936 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_422
timestamp 1698431365
transform 1 0 48608 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_430
timestamp 1698431365
transform 1 0 49504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_434
timestamp 1698431365
transform 1 0 49952 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_450
timestamp 1698431365
transform 1 0 51744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698431365
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_488
timestamp 1698431365
transform 1 0 56000 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_492
timestamp 1698431365
transform 1 0 56448 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_508
timestamp 1698431365
transform 1 0 58240 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_18
timestamp 1698431365
transform 1 0 3360 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_46
timestamp 1698431365
transform 1 0 6496 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_54
timestamp 1698431365
transform 1 0 7392 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_76
timestamp 1698431365
transform 1 0 9856 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_101
timestamp 1698431365
transform 1 0 12656 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_105
timestamp 1698431365
transform 1 0 13104 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_112
timestamp 1698431365
transform 1 0 13888 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_133
timestamp 1698431365
transform 1 0 16240 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_137
timestamp 1698431365
transform 1 0 16688 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_139
timestamp 1698431365
transform 1 0 16912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_172
timestamp 1698431365
transform 1 0 20608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_174
timestamp 1698431365
transform 1 0 20832 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_177
timestamp 1698431365
transform 1 0 21168 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_228
timestamp 1698431365
transform 1 0 26880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_238
timestamp 1698431365
transform 1 0 28000 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_244
timestamp 1698431365
transform 1 0 28672 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_298
timestamp 1698431365
transform 1 0 34720 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_306
timestamp 1698431365
transform 1 0 35616 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_308
timestamp 1698431365
transform 1 0 35840 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_324
timestamp 1698431365
transform 1 0 37632 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_340
timestamp 1698431365
transform 1 0 39424 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_348
timestamp 1698431365
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_356
timestamp 1698431365
transform 1 0 41216 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_362
timestamp 1698431365
transform 1 0 41888 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_364
timestamp 1698431365
transform 1 0 42112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_370
timestamp 1698431365
transform 1 0 42784 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_372
timestamp 1698431365
transform 1 0 43008 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_381
timestamp 1698431365
transform 1 0 44016 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_413
timestamp 1698431365
transform 1 0 47600 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_417
timestamp 1698431365
transform 1 0 48048 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_419
timestamp 1698431365
transform 1 0 48272 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_438
timestamp 1698431365
transform 1 0 50400 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_440
timestamp 1698431365
transform 1 0 50624 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_470
timestamp 1698431365
transform 1 0 53984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_474
timestamp 1698431365
transform 1 0 54432 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_480
timestamp 1698431365
transform 1 0 55104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_39
timestamp 1698431365
transform 1 0 5712 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_77
timestamp 1698431365
transform 1 0 9968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_81
timestamp 1698431365
transform 1 0 10416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_85
timestamp 1698431365
transform 1 0 10864 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_92
timestamp 1698431365
transform 1 0 11648 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_100
timestamp 1698431365
transform 1 0 12544 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_104
timestamp 1698431365
transform 1 0 12992 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_115
timestamp 1698431365
transform 1 0 14224 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_164
timestamp 1698431365
transform 1 0 19712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_174
timestamp 1698431365
transform 1 0 20832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_185
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_220
timestamp 1698431365
transform 1 0 25984 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_236
timestamp 1698431365
transform 1 0 27776 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_263
timestamp 1698431365
transform 1 0 30800 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_265
timestamp 1698431365
transform 1 0 31024 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_287
timestamp 1698431365
transform 1 0 33488 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_291
timestamp 1698431365
transform 1 0 33936 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_307
timestamp 1698431365
transform 1 0 35728 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_349
timestamp 1698431365
transform 1 0 40432 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_357
timestamp 1698431365
transform 1 0 41328 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_359
timestamp 1698431365
transform 1 0 41552 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_369
timestamp 1698431365
transform 1 0 42672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_375
timestamp 1698431365
transform 1 0 43344 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_383
timestamp 1698431365
transform 1 0 44240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_403
timestamp 1698431365
transform 1 0 46480 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_433
timestamp 1698431365
transform 1 0 49840 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_435
timestamp 1698431365
transform 1 0 50064 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_446
timestamp 1698431365
transform 1 0 51296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_450
timestamp 1698431365
transform 1 0 51744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_452
timestamp 1698431365
transform 1 0 51968 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_465
timestamp 1698431365
transform 1 0 53424 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_467
timestamp 1698431365
transform 1 0 53648 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_10
timestamp 1698431365
transform 1 0 2464 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_34
timestamp 1698431365
transform 1 0 5152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_38
timestamp 1698431365
transform 1 0 5600 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_54
timestamp 1698431365
transform 1 0 7392 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_82
timestamp 1698431365
transform 1 0 10528 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_108
timestamp 1698431365
transform 1 0 13440 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_122
timestamp 1698431365
transform 1 0 15008 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_138
timestamp 1698431365
transform 1 0 16800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_183
timestamp 1698431365
transform 1 0 21840 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_191
timestamp 1698431365
transform 1 0 22736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_195
timestamp 1698431365
transform 1 0 23184 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_202
timestamp 1698431365
transform 1 0 23968 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_228
timestamp 1698431365
transform 1 0 26880 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_236
timestamp 1698431365
transform 1 0 27776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_258
timestamp 1698431365
transform 1 0 30240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_262
timestamp 1698431365
transform 1 0 30688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_294
timestamp 1698431365
transform 1 0 34272 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_306
timestamp 1698431365
transform 1 0 35616 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_314
timestamp 1698431365
transform 1 0 36512 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_341
timestamp 1698431365
transform 1 0 39536 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_366
timestamp 1698431365
transform 1 0 42336 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_398
timestamp 1698431365
transform 1 0 45920 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_406
timestamp 1698431365
transform 1 0 46816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_408
timestamp 1698431365
transform 1 0 47040 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_413
timestamp 1698431365
transform 1 0 47600 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_417
timestamp 1698431365
transform 1 0 48048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_419
timestamp 1698431365
transform 1 0 48272 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_430
timestamp 1698431365
transform 1 0 49504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_432
timestamp 1698431365
transform 1 0 49728 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_435
timestamp 1698431365
transform 1 0 50064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_437
timestamp 1698431365
transform 1 0 50288 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_445
timestamp 1698431365
transform 1 0 51184 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_459
timestamp 1698431365
transform 1 0 52752 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_475
timestamp 1698431365
transform 1 0 54544 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_483
timestamp 1698431365
transform 1 0 55440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_487
timestamp 1698431365
transform 1 0 55888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_489
timestamp 1698431365
transform 1 0 56112 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_42
timestamp 1698431365
transform 1 0 6048 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_58
timestamp 1698431365
transform 1 0 7840 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_81
timestamp 1698431365
transform 1 0 10416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_83
timestamp 1698431365
transform 1 0 10640 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_94
timestamp 1698431365
transform 1 0 11872 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_102
timestamp 1698431365
transform 1 0 12768 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_104
timestamp 1698431365
transform 1 0 12992 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_109
timestamp 1698431365
transform 1 0 13552 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_118
timestamp 1698431365
transform 1 0 14560 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_150
timestamp 1698431365
transform 1 0 18144 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_158
timestamp 1698431365
transform 1 0 19040 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_166
timestamp 1698431365
transform 1 0 19936 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698431365
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_209
timestamp 1698431365
transform 1 0 24752 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_211
timestamp 1698431365
transform 1 0 24976 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_243
timestamp 1698431365
transform 1 0 28560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_267
timestamp 1698431365
transform 1 0 31248 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_271
timestamp 1698431365
transform 1 0 31696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_273
timestamp 1698431365
transform 1 0 31920 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_289
timestamp 1698431365
transform 1 0 33712 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_293
timestamp 1698431365
transform 1 0 34160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_295
timestamp 1698431365
transform 1 0 34384 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_325
timestamp 1698431365
transform 1 0 37744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_329
timestamp 1698431365
transform 1 0 38192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_368
timestamp 1698431365
transform 1 0 42560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_372
timestamp 1698431365
transform 1 0 43008 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_380
timestamp 1698431365
transform 1 0 43904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_395
timestamp 1698431365
transform 1 0 45584 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_399
timestamp 1698431365
transform 1 0 46032 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_403
timestamp 1698431365
transform 1 0 46480 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_413
timestamp 1698431365
transform 1 0 47600 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_417
timestamp 1698431365
transform 1 0 48048 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_449
timestamp 1698431365
transform 1 0 51632 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_453
timestamp 1698431365
transform 1 0 52080 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_473
timestamp 1698431365
transform 1 0 54320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_477
timestamp 1698431365
transform 1 0 54768 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_10
timestamp 1698431365
transform 1 0 2464 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_14
timestamp 1698431365
transform 1 0 2912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_44
timestamp 1698431365
transform 1 0 6272 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_60
timestamp 1698431365
transform 1 0 8064 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1698431365
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_88
timestamp 1698431365
transform 1 0 11200 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_96
timestamp 1698431365
transform 1 0 12096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_100
timestamp 1698431365
transform 1 0 12544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_102
timestamp 1698431365
transform 1 0 12768 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_110
timestamp 1698431365
transform 1 0 13664 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_126
timestamp 1698431365
transform 1 0 15456 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_134
timestamp 1698431365
transform 1 0 16352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_138
timestamp 1698431365
transform 1 0 16800 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_228
timestamp 1698431365
transform 1 0 26880 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_236
timestamp 1698431365
transform 1 0 27776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_240
timestamp 1698431365
transform 1 0 28224 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_260
timestamp 1698431365
transform 1 0 30464 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_279
timestamp 1698431365
transform 1 0 32592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_298
timestamp 1698431365
transform 1 0 34720 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_306
timestamp 1698431365
transform 1 0 35616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_335
timestamp 1698431365
transform 1 0 38864 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_343
timestamp 1698431365
transform 1 0 39760 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_347
timestamp 1698431365
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_363
timestamp 1698431365
transform 1 0 42000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_367
timestamp 1698431365
transform 1 0 42448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_371
timestamp 1698431365
transform 1 0 42896 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_373
timestamp 1698431365
transform 1 0 43120 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_405
timestamp 1698431365
transform 1 0 46704 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_426
timestamp 1698431365
transform 1 0 49056 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_442
timestamp 1698431365
transform 1 0 50848 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_446
timestamp 1698431365
transform 1 0 51296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_448
timestamp 1698431365
transform 1 0 51520 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_465
timestamp 1698431365
transform 1 0 53424 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_473
timestamp 1698431365
transform 1 0 54320 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_477
timestamp 1698431365
transform 1 0 54768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1698431365
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_500
timestamp 1698431365
transform 1 0 57344 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_18
timestamp 1698431365
transform 1 0 3360 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_26
timestamp 1698431365
transform 1 0 4256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_28
timestamp 1698431365
transform 1 0 4480 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_31
timestamp 1698431365
transform 1 0 4816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_45
timestamp 1698431365
transform 1 0 6384 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_49
timestamp 1698431365
transform 1 0 6832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_51
timestamp 1698431365
transform 1 0 7056 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_69
timestamp 1698431365
transform 1 0 9072 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_73
timestamp 1698431365
transform 1 0 9520 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_82
timestamp 1698431365
transform 1 0 10528 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_86
timestamp 1698431365
transform 1 0 10976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_88
timestamp 1698431365
transform 1 0 11200 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_95
timestamp 1698431365
transform 1 0 11984 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_104
timestamp 1698431365
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_137
timestamp 1698431365
transform 1 0 16688 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_145
timestamp 1698431365
transform 1 0 17584 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_149
timestamp 1698431365
transform 1 0 18032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_151
timestamp 1698431365
transform 1 0 18256 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_164
timestamp 1698431365
transform 1 0 19712 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_166
timestamp 1698431365
transform 1 0 19936 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_181
timestamp 1698431365
transform 1 0 21616 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_185
timestamp 1698431365
transform 1 0 22064 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_210
timestamp 1698431365
transform 1 0 24864 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_242
timestamp 1698431365
transform 1 0 28448 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1698431365
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_255
timestamp 1698431365
transform 1 0 29904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_259
timestamp 1698431365
transform 1 0 30352 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_292
timestamp 1698431365
transform 1 0 34048 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_300
timestamp 1698431365
transform 1 0 34944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_302
timestamp 1698431365
transform 1 0 35168 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1698431365
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_321
timestamp 1698431365
transform 1 0 37296 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_329
timestamp 1698431365
transform 1 0 38192 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_333
timestamp 1698431365
transform 1 0 38640 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_342
timestamp 1698431365
transform 1 0 39648 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_358
timestamp 1698431365
transform 1 0 41440 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_366
timestamp 1698431365
transform 1 0 42336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_370
timestamp 1698431365
transform 1 0 42784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_380
timestamp 1698431365
transform 1 0 43904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_447
timestamp 1698431365
transform 1 0 51408 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698431365
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_465
timestamp 1698431365
transform 1 0 53424 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_469
timestamp 1698431365
transform 1 0 53872 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_476
timestamp 1698431365
transform 1 0 54656 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_484
timestamp 1698431365
transform 1 0 55552 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_493
timestamp 1698431365
transform 1 0 56560 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_18
timestamp 1698431365
transform 1 0 3360 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_26
timestamp 1698431365
transform 1 0 4256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_30
timestamp 1698431365
transform 1 0 4704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_32
timestamp 1698431365
transform 1 0 4928 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_76
timestamp 1698431365
transform 1 0 9856 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_107
timestamp 1698431365
transform 1 0 13328 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_111
timestamp 1698431365
transform 1 0 13776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_115
timestamp 1698431365
transform 1 0 14224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_117
timestamp 1698431365
transform 1 0 14448 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_123
timestamp 1698431365
transform 1 0 15120 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698431365
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_216
timestamp 1698431365
transform 1 0 25536 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_248
timestamp 1698431365
transform 1 0 29120 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_264
timestamp 1698431365
transform 1 0 30912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_284
timestamp 1698431365
transform 1 0 33152 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_297
timestamp 1698431365
transform 1 0 34608 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_318
timestamp 1698431365
transform 1 0 36960 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_356
timestamp 1698431365
transform 1 0 41216 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_364
timestamp 1698431365
transform 1 0 42112 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_395
timestamp 1698431365
transform 1 0 45584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_399
timestamp 1698431365
transform 1 0 46032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_410
timestamp 1698431365
transform 1 0 47264 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_414
timestamp 1698431365
transform 1 0 47712 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1698431365
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_438
timestamp 1698431365
transform 1 0 50400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_477
timestamp 1698431365
transform 1 0 54768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_481
timestamp 1698431365
transform 1 0 55216 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_496
timestamp 1698431365
transform 1 0 56896 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_498
timestamp 1698431365
transform 1 0 57120 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_10
timestamp 1698431365
transform 1 0 2464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_12
timestamp 1698431365
transform 1 0 2688 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_30
timestamp 1698431365
transform 1 0 4704 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_45
timestamp 1698431365
transform 1 0 6384 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_49
timestamp 1698431365
transform 1 0 6832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_71
timestamp 1698431365
transform 1 0 9296 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_85
timestamp 1698431365
transform 1 0 10864 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_139
timestamp 1698431365
transform 1 0 16912 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_143
timestamp 1698431365
transform 1 0 17360 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698431365
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_185
timestamp 1698431365
transform 1 0 22064 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_211
timestamp 1698431365
transform 1 0 24976 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_261
timestamp 1698431365
transform 1 0 30576 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_277
timestamp 1698431365
transform 1 0 32368 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_281
timestamp 1698431365
transform 1 0 32816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_285
timestamp 1698431365
transform 1 0 33264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_287
timestamp 1698431365
transform 1 0 33488 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_337
timestamp 1698431365
transform 1 0 39088 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_351
timestamp 1698431365
transform 1 0 40656 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_362
timestamp 1698431365
transform 1 0 41888 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_378
timestamp 1698431365
transform 1 0 43680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_382
timestamp 1698431365
transform 1 0 44128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1698431365
transform 1 0 44352 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_419
timestamp 1698431365
transform 1 0 48272 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_435
timestamp 1698431365
transform 1 0 50064 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_443
timestamp 1698431365
transform 1 0 50960 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_463
timestamp 1698431365
transform 1 0 53200 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_467
timestamp 1698431365
transform 1 0 53648 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_39
timestamp 1698431365
transform 1 0 5712 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_55
timestamp 1698431365
transform 1 0 7504 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_63
timestamp 1698431365
transform 1 0 8400 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_67
timestamp 1698431365
transform 1 0 8848 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_69
timestamp 1698431365
transform 1 0 9072 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_80
timestamp 1698431365
transform 1 0 10304 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_84
timestamp 1698431365
transform 1 0 10752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_91
timestamp 1698431365
transform 1 0 11536 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_107
timestamp 1698431365
transform 1 0 13328 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_111
timestamp 1698431365
transform 1 0 13776 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_139
timestamp 1698431365
transform 1 0 16912 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_150
timestamp 1698431365
transform 1 0 18144 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_153
timestamp 1698431365
transform 1 0 18480 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_185
timestamp 1698431365
transform 1 0 22064 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_201
timestamp 1698431365
transform 1 0 23856 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698431365
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_220
timestamp 1698431365
transform 1 0 25984 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_224
timestamp 1698431365
transform 1 0 26432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_253
timestamp 1698431365
transform 1 0 29680 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_257
timestamp 1698431365
transform 1 0 30128 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_271
timestamp 1698431365
transform 1 0 31696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_275
timestamp 1698431365
transform 1 0 32144 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_279
timestamp 1698431365
transform 1 0 32592 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_314
timestamp 1698431365
transform 1 0 36512 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_330
timestamp 1698431365
transform 1 0 38304 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_338
timestamp 1698431365
transform 1 0 39200 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_347
timestamp 1698431365
transform 1 0 40208 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1698431365
transform 1 0 40432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_369
timestamp 1698431365
transform 1 0 42672 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_385
timestamp 1698431365
transform 1 0 44464 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_393
timestamp 1698431365
transform 1 0 45360 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_410
timestamp 1698431365
transform 1 0 47264 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_418
timestamp 1698431365
transform 1 0 48160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_438
timestamp 1698431365
transform 1 0 50400 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_440
timestamp 1698431365
transform 1 0 50624 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_453
timestamp 1698431365
transform 1 0 52080 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_469
timestamp 1698431365
transform 1 0 53872 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_473
timestamp 1698431365
transform 1 0 54320 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_482
timestamp 1698431365
transform 1 0 55328 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_500
timestamp 1698431365
transform 1 0 57344 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_10
timestamp 1698431365
transform 1 0 2464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_12
timestamp 1698431365
transform 1 0 2688 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_69
timestamp 1698431365
transform 1 0 9072 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_90
timestamp 1698431365
transform 1 0 11424 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_92
timestamp 1698431365
transform 1 0 11648 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_95
timestamp 1698431365
transform 1 0 11984 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_99
timestamp 1698431365
transform 1 0 12432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_103
timestamp 1698431365
transform 1 0 12880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_111
timestamp 1698431365
transform 1 0 13776 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_115
timestamp 1698431365
transform 1 0 14224 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_120
timestamp 1698431365
transform 1 0 14784 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_154
timestamp 1698431365
transform 1 0 18592 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_170
timestamp 1698431365
transform 1 0 20384 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1698431365
transform 1 0 20832 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_193
timestamp 1698431365
transform 1 0 22960 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_203
timestamp 1698431365
transform 1 0 24080 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_219
timestamp 1698431365
transform 1 0 25872 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_227
timestamp 1698431365
transform 1 0 26768 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_231
timestamp 1698431365
transform 1 0 27216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_233
timestamp 1698431365
transform 1 0 27440 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_242
timestamp 1698431365
transform 1 0 28448 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1698431365
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_272
timestamp 1698431365
transform 1 0 31808 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_292
timestamp 1698431365
transform 1 0 34048 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_294
timestamp 1698431365
transform 1 0 34272 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_305
timestamp 1698431365
transform 1 0 35504 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_313
timestamp 1698431365
transform 1 0 36400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_321
timestamp 1698431365
transform 1 0 37296 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_375
timestamp 1698431365
transform 1 0 43344 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_416
timestamp 1698431365
transform 1 0 47936 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_424
timestamp 1698431365
transform 1 0 48832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_432
timestamp 1698431365
transform 1 0 49728 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_439
timestamp 1698431365
transform 1 0 50512 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_466
timestamp 1698431365
transform 1 0 53536 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_474
timestamp 1698431365
transform 1 0 54432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_505
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_26
timestamp 1698431365
transform 1 0 4256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_28
timestamp 1698431365
transform 1 0 4480 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_31
timestamp 1698431365
transform 1 0 4816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_33
timestamp 1698431365
transform 1 0 5040 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_52
timestamp 1698431365
transform 1 0 7168 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_68
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_74
timestamp 1698431365
transform 1 0 9632 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_77
timestamp 1698431365
transform 1 0 9968 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_86
timestamp 1698431365
transform 1 0 10976 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_93
timestamp 1698431365
transform 1 0 11760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_116
timestamp 1698431365
transform 1 0 14336 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_133
timestamp 1698431365
transform 1 0 16240 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_137
timestamp 1698431365
transform 1 0 16688 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_139
timestamp 1698431365
transform 1 0 16912 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_152
timestamp 1698431365
transform 1 0 18368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_177
timestamp 1698431365
transform 1 0 21168 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_185
timestamp 1698431365
transform 1 0 22064 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_209
timestamp 1698431365
transform 1 0 24752 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_216
timestamp 1698431365
transform 1 0 25536 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_232
timestamp 1698431365
transform 1 0 27328 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_244
timestamp 1698431365
transform 1 0 28672 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_260
timestamp 1698431365
transform 1 0 30464 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_264
timestamp 1698431365
transform 1 0 30912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_266
timestamp 1698431365
transform 1 0 31136 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_269
timestamp 1698431365
transform 1 0 31472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_344
timestamp 1698431365
transform 1 0 39872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_348
timestamp 1698431365
transform 1 0 40320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_384
timestamp 1698431365
transform 1 0 44352 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_392
timestamp 1698431365
transform 1 0 45248 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_397
timestamp 1698431365
transform 1 0 45808 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_419
timestamp 1698431365
transform 1 0 48272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_426
timestamp 1698431365
transform 1 0 49056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_430
timestamp 1698431365
transform 1 0 49504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_432
timestamp 1698431365
transform 1 0 49728 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_439
timestamp 1698431365
transform 1 0 50512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_470
timestamp 1698431365
transform 1 0 53984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_474
timestamp 1698431365
transform 1 0 54432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_488
timestamp 1698431365
transform 1 0 56000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_492
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_18
timestamp 1698431365
transform 1 0 3360 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_45
timestamp 1698431365
transform 1 0 6384 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_87
timestamp 1698431365
transform 1 0 11088 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_91
timestamp 1698431365
transform 1 0 11536 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_93
timestamp 1698431365
transform 1 0 11760 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_102
timestamp 1698431365
transform 1 0 12768 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_104
timestamp 1698431365
transform 1 0 12992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_125
timestamp 1698431365
transform 1 0 15344 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_129
timestamp 1698431365
transform 1 0 15792 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_131
timestamp 1698431365
transform 1 0 16016 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_171
timestamp 1698431365
transform 1 0 20496 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_233
timestamp 1698431365
transform 1 0 27440 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_237
timestamp 1698431365
transform 1 0 27888 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_249
timestamp 1698431365
transform 1 0 29232 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_265
timestamp 1698431365
transform 1 0 31024 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_298
timestamp 1698431365
transform 1 0 34720 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_302
timestamp 1698431365
transform 1 0 35168 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_306
timestamp 1698431365
transform 1 0 35616 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_329
timestamp 1698431365
transform 1 0 38192 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_361
timestamp 1698431365
transform 1 0 41776 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_379
timestamp 1698431365
transform 1 0 43792 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_383
timestamp 1698431365
transform 1 0 44240 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_403
timestamp 1698431365
transform 1 0 46480 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_436
timestamp 1698431365
transform 1 0 50176 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_440
timestamp 1698431365
transform 1 0 50624 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_448
timestamp 1698431365
transform 1 0 51520 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_452
timestamp 1698431365
transform 1 0 51968 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_454
timestamp 1698431365
transform 1 0 52192 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_473
timestamp 1698431365
transform 1 0 54320 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_477
timestamp 1698431365
transform 1 0 54768 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_479
timestamp 1698431365
transform 1 0 54992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_486
timestamp 1698431365
transform 1 0 55776 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_502
timestamp 1698431365
transform 1 0 57568 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_506
timestamp 1698431365
transform 1 0 58016 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_508
timestamp 1698431365
transform 1 0 58240 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_51
timestamp 1698431365
transform 1 0 7056 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_55
timestamp 1698431365
transform 1 0 7504 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_57
timestamp 1698431365
transform 1 0 7728 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_66
timestamp 1698431365
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_85
timestamp 1698431365
transform 1 0 10864 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_101
timestamp 1698431365
transform 1 0 12656 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_105
timestamp 1698431365
transform 1 0 13104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_114
timestamp 1698431365
transform 1 0 14112 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_130
timestamp 1698431365
transform 1 0 15904 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_138
timestamp 1698431365
transform 1 0 16800 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_158
timestamp 1698431365
transform 1 0 19040 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_160
timestamp 1698431365
transform 1 0 19264 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_174
timestamp 1698431365
transform 1 0 20832 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_182
timestamp 1698431365
transform 1 0 21728 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_186
timestamp 1698431365
transform 1 0 22176 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_188
timestamp 1698431365
transform 1 0 22400 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_243
timestamp 1698431365
transform 1 0 28560 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_247
timestamp 1698431365
transform 1 0 29008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_272
timestamp 1698431365
transform 1 0 31808 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_279
timestamp 1698431365
transform 1 0 32592 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_286
timestamp 1698431365
transform 1 0 33376 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_302
timestamp 1698431365
transform 1 0 35168 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_306
timestamp 1698431365
transform 1 0 35616 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_308
timestamp 1698431365
transform 1 0 35840 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_338
timestamp 1698431365
transform 1 0 39200 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_346
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_360
timestamp 1698431365
transform 1 0 41664 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_393
timestamp 1698431365
transform 1 0 45360 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_409
timestamp 1698431365
transform 1 0 47152 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_417
timestamp 1698431365
transform 1 0 48048 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_419
timestamp 1698431365
transform 1 0 48272 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_438
timestamp 1698431365
transform 1 0 50400 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_442
timestamp 1698431365
transform 1 0 50848 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_454
timestamp 1698431365
transform 1 0 52192 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_456
timestamp 1698431365
transform 1 0 52416 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_459
timestamp 1698431365
transform 1 0 52752 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_475
timestamp 1698431365
transform 1 0 54544 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_483
timestamp 1698431365
transform 1 0 55440 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_487
timestamp 1698431365
transform 1 0 55888 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_489
timestamp 1698431365
transform 1 0 56112 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_508
timestamp 1698431365
transform 1 0 58240 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_10
timestamp 1698431365
transform 1 0 2464 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_18
timestamp 1698431365
transform 1 0 3360 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_20
timestamp 1698431365
transform 1 0 3584 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_29
timestamp 1698431365
transform 1 0 4592 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_33
timestamp 1698431365
transform 1 0 5040 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_42
timestamp 1698431365
transform 1 0 6048 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_74
timestamp 1698431365
transform 1 0 9632 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_76
timestamp 1698431365
transform 1 0 9856 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_100
timestamp 1698431365
transform 1 0 12544 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_104
timestamp 1698431365
transform 1 0 12992 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_113
timestamp 1698431365
transform 1 0 14000 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_119
timestamp 1698431365
transform 1 0 14672 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_123
timestamp 1698431365
transform 1 0 15120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_127
timestamp 1698431365
transform 1 0 15568 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_139
timestamp 1698431365
transform 1 0 16912 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_171
timestamp 1698431365
transform 1 0 20496 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_209
timestamp 1698431365
transform 1 0 24752 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_218
timestamp 1698431365
transform 1 0 25760 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_222
timestamp 1698431365
transform 1 0 26208 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1698431365
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_251
timestamp 1698431365
transform 1 0 29456 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_264
timestamp 1698431365
transform 1 0 30912 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_296
timestamp 1698431365
transform 1 0 34496 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_304
timestamp 1698431365
transform 1 0 35392 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_314
timestamp 1698431365
transform 1 0 36512 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_325
timestamp 1698431365
transform 1 0 37744 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_329
timestamp 1698431365
transform 1 0 38192 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_359
timestamp 1698431365
transform 1 0 41552 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_363
timestamp 1698431365
transform 1 0 42000 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_376
timestamp 1698431365
transform 1 0 43456 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_384
timestamp 1698431365
transform 1 0 44352 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_416
timestamp 1698431365
transform 1 0 47936 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_420
timestamp 1698431365
transform 1 0 48384 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_436
timestamp 1698431365
transform 1 0 50176 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_444
timestamp 1698431365
transform 1 0 51072 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_448
timestamp 1698431365
transform 1 0 51520 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_450
timestamp 1698431365
transform 1 0 51744 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_457
timestamp 1698431365
transform 1 0 52528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_485
timestamp 1698431365
transform 1 0 55664 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_501
timestamp 1698431365
transform 1 0 57456 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_505
timestamp 1698431365
transform 1 0 57904 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_6
timestamp 1698431365
transform 1 0 2016 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_38
timestamp 1698431365
transform 1 0 5600 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_46
timestamp 1698431365
transform 1 0 6496 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_50
timestamp 1698431365
transform 1 0 6944 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_52
timestamp 1698431365
transform 1 0 7168 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_59
timestamp 1698431365
transform 1 0 7952 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_63
timestamp 1698431365
transform 1 0 8400 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_67
timestamp 1698431365
transform 1 0 8848 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_69
timestamp 1698431365
transform 1 0 9072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_88
timestamp 1698431365
transform 1 0 11200 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_125
timestamp 1698431365
transform 1 0 15344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_139
timestamp 1698431365
transform 1 0 16912 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_151
timestamp 1698431365
transform 1 0 18256 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_183
timestamp 1698431365
transform 1 0 21840 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_199
timestamp 1698431365
transform 1 0 23632 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_207
timestamp 1698431365
transform 1 0 24528 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_209
timestamp 1698431365
transform 1 0 24752 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_234
timestamp 1698431365
transform 1 0 27552 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_238
timestamp 1698431365
transform 1 0 28000 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_254
timestamp 1698431365
transform 1 0 29792 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_262
timestamp 1698431365
transform 1 0 30688 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_266
timestamp 1698431365
transform 1 0 31136 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_274
timestamp 1698431365
transform 1 0 32032 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_278
timestamp 1698431365
transform 1 0 32480 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_298
timestamp 1698431365
transform 1 0 34720 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_302
timestamp 1698431365
transform 1 0 35168 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_323
timestamp 1698431365
transform 1 0 37520 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_331
timestamp 1698431365
transform 1 0 38416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_335
timestamp 1698431365
transform 1 0 38864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_337
timestamp 1698431365
transform 1 0 39088 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_360
timestamp 1698431365
transform 1 0 41664 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_375
timestamp 1698431365
transform 1 0 43344 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_383
timestamp 1698431365
transform 1 0 44240 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_387
timestamp 1698431365
transform 1 0 44688 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_394
timestamp 1698431365
transform 1 0 45472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_398
timestamp 1698431365
transform 1 0 45920 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_414
timestamp 1698431365
transform 1 0 47712 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_436
timestamp 1698431365
transform 1 0 50176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_440
timestamp 1698431365
transform 1 0 50624 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_444
timestamp 1698431365
transform 1 0 51072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_474
timestamp 1698431365
transform 1 0 54432 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_478
timestamp 1698431365
transform 1 0 54880 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_482
timestamp 1698431365
transform 1 0 55328 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_486
timestamp 1698431365
transform 1 0 55776 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_498
timestamp 1698431365
transform 1 0 57120 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_500
timestamp 1698431365
transform 1 0 57344 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_39
timestamp 1698431365
transform 1 0 5712 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_42
timestamp 1698431365
transform 1 0 6048 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_59
timestamp 1698431365
transform 1 0 7952 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_90
timestamp 1698431365
transform 1 0 11424 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_130
timestamp 1698431365
transform 1 0 15904 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_149
timestamp 1698431365
transform 1 0 18032 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_181
timestamp 1698431365
transform 1 0 21616 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_183
timestamp 1698431365
transform 1 0 21840 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_186
timestamp 1698431365
transform 1 0 22176 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_188
timestamp 1698431365
transform 1 0 22400 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_231
timestamp 1698431365
transform 1 0 27216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_243
timestamp 1698431365
transform 1 0 28560 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_252
timestamp 1698431365
transform 1 0 29568 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_256
timestamp 1698431365
transform 1 0 30016 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_286
timestamp 1698431365
transform 1 0 33376 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_290
timestamp 1698431365
transform 1 0 33824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_300
timestamp 1698431365
transform 1 0 34944 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_308
timestamp 1698431365
transform 1 0 35840 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_312
timestamp 1698431365
transform 1 0 36288 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_314
timestamp 1698431365
transform 1 0 36512 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_335
timestamp 1698431365
transform 1 0 38864 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_343
timestamp 1698431365
transform 1 0 39760 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_403
timestamp 1698431365
transform 1 0 46480 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_405
timestamp 1698431365
transform 1 0 46704 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_457
timestamp 1698431365
transform 1 0 52528 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_473
timestamp 1698431365
transform 1 0 54320 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_477
timestamp 1698431365
transform 1 0 54768 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_2
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_10
timestamp 1698431365
transform 1 0 2464 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_63
timestamp 1698431365
transform 1 0 8400 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_67
timestamp 1698431365
transform 1 0 8848 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_69
timestamp 1698431365
transform 1 0 9072 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_80
timestamp 1698431365
transform 1 0 10304 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_82
timestamp 1698431365
transform 1 0 10528 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_109
timestamp 1698431365
transform 1 0 13552 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_113
timestamp 1698431365
transform 1 0 14000 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_117
timestamp 1698431365
transform 1 0 14448 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_133
timestamp 1698431365
transform 1 0 16240 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_137
timestamp 1698431365
transform 1 0 16688 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_139
timestamp 1698431365
transform 1 0 16912 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_152
timestamp 1698431365
transform 1 0 18368 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_154
timestamp 1698431365
transform 1 0 18592 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_223
timestamp 1698431365
transform 1 0 26320 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_227
timestamp 1698431365
transform 1 0 26768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_258
timestamp 1698431365
transform 1 0 30240 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_262
timestamp 1698431365
transform 1 0 30688 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_278
timestamp 1698431365
transform 1 0 32480 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_318
timestamp 1698431365
transform 1 0 36960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_348
timestamp 1698431365
transform 1 0 40320 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_360
timestamp 1698431365
transform 1 0 41664 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_364
timestamp 1698431365
transform 1 0 42112 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_372
timestamp 1698431365
transform 1 0 43008 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_404
timestamp 1698431365
transform 1 0 46592 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_422
timestamp 1698431365
transform 1 0 48608 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_437
timestamp 1698431365
transform 1 0 50288 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_441
timestamp 1698431365
transform 1 0 50736 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_448
timestamp 1698431365
transform 1 0 51520 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_456
timestamp 1698431365
transform 1 0 52416 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_466
timestamp 1698431365
transform 1 0 53536 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_508
timestamp 1698431365
transform 1 0 58240 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698431365
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_52
timestamp 1698431365
transform 1 0 7168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_54
timestamp 1698431365
transform 1 0 7392 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_57
timestamp 1698431365
transform 1 0 7728 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_89
timestamp 1698431365
transform 1 0 11312 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_99
timestamp 1698431365
transform 1 0 12432 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_103
timestamp 1698431365
transform 1 0 12880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_139
timestamp 1698431365
transform 1 0 16912 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_155
timestamp 1698431365
transform 1 0 18704 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_163
timestamp 1698431365
transform 1 0 19600 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_171
timestamp 1698431365
transform 1 0 20496 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_179
timestamp 1698431365
transform 1 0 21392 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_213
timestamp 1698431365
transform 1 0 25200 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_217
timestamp 1698431365
transform 1 0 25648 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_221
timestamp 1698431365
transform 1 0 26096 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_237
timestamp 1698431365
transform 1 0 27888 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_263
timestamp 1698431365
transform 1 0 30800 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_271
timestamp 1698431365
transform 1 0 31696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_275
timestamp 1698431365
transform 1 0 32144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_282
timestamp 1698431365
transform 1 0 32928 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_290
timestamp 1698431365
transform 1 0 33824 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_325
timestamp 1698431365
transform 1 0 37744 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_327
timestamp 1698431365
transform 1 0 37968 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_334
timestamp 1698431365
transform 1 0 38752 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_366
timestamp 1698431365
transform 1 0 42336 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_380
timestamp 1698431365
transform 1 0 43904 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_384
timestamp 1698431365
transform 1 0 44352 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_387
timestamp 1698431365
transform 1 0 44688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_391
timestamp 1698431365
transform 1 0 45136 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_423
timestamp 1698431365
transform 1 0 48720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_429
timestamp 1698431365
transform 1 0 49392 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_445
timestamp 1698431365
transform 1 0 51184 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_453
timestamp 1698431365
transform 1 0 52080 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_507
timestamp 1698431365
transform 1 0 58128 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_34
timestamp 1698431365
transform 1 0 5152 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_42
timestamp 1698431365
transform 1 0 6048 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_46
timestamp 1698431365
transform 1 0 6496 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_55
timestamp 1698431365
transform 1 0 7504 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_67
timestamp 1698431365
transform 1 0 8848 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_69
timestamp 1698431365
transform 1 0 9072 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_87
timestamp 1698431365
transform 1 0 11088 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_95
timestamp 1698431365
transform 1 0 11984 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_99
timestamp 1698431365
transform 1 0 12432 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_101
timestamp 1698431365
transform 1 0 12656 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_115
timestamp 1698431365
transform 1 0 14224 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_125
timestamp 1698431365
transform 1 0 15344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_129
timestamp 1698431365
transform 1 0 15792 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_138
timestamp 1698431365
transform 1 0 16800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_150
timestamp 1698431365
transform 1 0 18144 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_154
timestamp 1698431365
transform 1 0 18592 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_172
timestamp 1698431365
transform 1 0 20608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_176
timestamp 1698431365
transform 1 0 21056 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_208
timestamp 1698431365
transform 1 0 24640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_228
timestamp 1698431365
transform 1 0 26880 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_232
timestamp 1698431365
transform 1 0 27328 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_234
timestamp 1698431365
transform 1 0 27552 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_237
timestamp 1698431365
transform 1 0 27888 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_253
timestamp 1698431365
transform 1 0 29680 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_261
timestamp 1698431365
transform 1 0 30576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_265
timestamp 1698431365
transform 1 0 31024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_269
timestamp 1698431365
transform 1 0 31472 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_277
timestamp 1698431365
transform 1 0 32368 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_279
timestamp 1698431365
transform 1 0 32592 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_314
timestamp 1698431365
transform 1 0 36512 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_328
timestamp 1698431365
transform 1 0 38080 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_342
timestamp 1698431365
transform 1 0 39648 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_384
timestamp 1698431365
transform 1 0 44352 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_412
timestamp 1698431365
transform 1 0 47488 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_451
timestamp 1698431365
transform 1 0 51856 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_463
timestamp 1698431365
transform 1 0 53200 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_503
timestamp 1698431365
transform 1 0 57680 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_507
timestamp 1698431365
transform 1 0 58128 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_2
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_53
timestamp 1698431365
transform 1 0 7280 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_67
timestamp 1698431365
transform 1 0 8848 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_83
timestamp 1698431365
transform 1 0 10640 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_91
timestamp 1698431365
transform 1 0 11536 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_103
timestamp 1698431365
transform 1 0 12880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_111
timestamp 1698431365
transform 1 0 13776 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_150
timestamp 1698431365
transform 1 0 18144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_154
timestamp 1698431365
transform 1 0 18592 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_168
timestamp 1698431365
transform 1 0 20160 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_172
timestamp 1698431365
transform 1 0 20608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_174
timestamp 1698431365
transform 1 0 20832 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_203
timestamp 1698431365
transform 1 0 24080 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_219
timestamp 1698431365
transform 1 0 25872 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_241
timestamp 1698431365
transform 1 0 28336 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_249
timestamp 1698431365
transform 1 0 29232 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_262
timestamp 1698431365
transform 1 0 30688 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_264
timestamp 1698431365
transform 1 0 30912 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_270
timestamp 1698431365
transform 1 0 31584 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_279
timestamp 1698431365
transform 1 0 32592 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_283
timestamp 1698431365
transform 1 0 33040 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_333
timestamp 1698431365
transform 1 0 38640 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_341
timestamp 1698431365
transform 1 0 39536 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_345
timestamp 1698431365
transform 1 0 39984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_378
timestamp 1698431365
transform 1 0 43680 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_416
timestamp 1698431365
transform 1 0 47936 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_432
timestamp 1698431365
transform 1 0 49728 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_436
timestamp 1698431365
transform 1 0 50176 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_452
timestamp 1698431365
transform 1 0 51968 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_454
timestamp 1698431365
transform 1 0 52192 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_457
timestamp 1698431365
transform 1 0 52528 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_459
timestamp 1698431365
transform 1 0 52752 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_476
timestamp 1698431365
transform 1 0 54656 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_34
timestamp 1698431365
transform 1 0 5152 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_50
timestamp 1698431365
transform 1 0 6944 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_58
timestamp 1698431365
transform 1 0 7840 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_66
timestamp 1698431365
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_80
timestamp 1698431365
transform 1 0 10304 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_150
timestamp 1698431365
transform 1 0 18144 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_195
timestamp 1698431365
transform 1 0 23184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_199
timestamp 1698431365
transform 1 0 23632 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_207
timestamp 1698431365
transform 1 0 24528 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_209
timestamp 1698431365
transform 1 0 24752 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_266
timestamp 1698431365
transform 1 0 31136 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_306
timestamp 1698431365
transform 1 0 35616 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_338
timestamp 1698431365
transform 1 0 39200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_342
timestamp 1698431365
transform 1 0 39648 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_352
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_356
timestamp 1698431365
transform 1 0 41216 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_358
timestamp 1698431365
transform 1 0 41440 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_361
timestamp 1698431365
transform 1 0 41776 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_365
timestamp 1698431365
transform 1 0 42224 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_369
timestamp 1698431365
transform 1 0 42672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_377
timestamp 1698431365
transform 1 0 43568 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_381
timestamp 1698431365
transform 1 0 44016 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_397
timestamp 1698431365
transform 1 0 45808 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_401
timestamp 1698431365
transform 1 0 46256 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_410
timestamp 1698431365
transform 1 0 47264 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_418
timestamp 1698431365
transform 1 0 48160 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_422
timestamp 1698431365
transform 1 0 48608 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_426
timestamp 1698431365
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_442
timestamp 1698431365
transform 1 0 50848 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_444
timestamp 1698431365
transform 1 0 51072 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_479
timestamp 1698431365
transform 1 0 54992 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_487
timestamp 1698431365
transform 1 0 55888 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_498
timestamp 1698431365
transform 1 0 57120 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_506
timestamp 1698431365
transform 1 0 58016 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_508
timestamp 1698431365
transform 1 0 58240 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_2
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_66
timestamp 1698431365
transform 1 0 8736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_68
timestamp 1698431365
transform 1 0 8960 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_98
timestamp 1698431365
transform 1 0 12320 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_113
timestamp 1698431365
transform 1 0 14000 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_145
timestamp 1698431365
transform 1 0 17584 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_177
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_181
timestamp 1698431365
transform 1 0 21616 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_189
timestamp 1698431365
transform 1 0 22512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_193
timestamp 1698431365
transform 1 0 22960 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_238
timestamp 1698431365
transform 1 0 28000 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_242
timestamp 1698431365
transform 1 0 28448 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_255
timestamp 1698431365
transform 1 0 29904 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_267
timestamp 1698431365
transform 1 0 31248 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_271
timestamp 1698431365
transform 1 0 31696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_275
timestamp 1698431365
transform 1 0 32144 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_321
timestamp 1698431365
transform 1 0 37296 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_329
timestamp 1698431365
transform 1 0 38192 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_387
timestamp 1698431365
transform 1 0 44688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_391
timestamp 1698431365
transform 1 0 45136 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_395
timestamp 1698431365
transform 1 0 45584 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_403
timestamp 1698431365
transform 1 0 46480 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_407
timestamp 1698431365
transform 1 0 46928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_439
timestamp 1698431365
transform 1 0 50512 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_447
timestamp 1698431365
transform 1 0 51408 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_452
timestamp 1698431365
transform 1 0 51968 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_454
timestamp 1698431365
transform 1 0 52192 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_457
timestamp 1698431365
transform 1 0 52528 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_461
timestamp 1698431365
transform 1 0 52976 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_469
timestamp 1698431365
transform 1 0 53872 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_478
timestamp 1698431365
transform 1 0 54880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_2
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_68
timestamp 1698431365
transform 1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_88
timestamp 1698431365
transform 1 0 11200 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_96
timestamp 1698431365
transform 1 0 12096 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_100
timestamp 1698431365
transform 1 0 12544 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_132
timestamp 1698431365
transform 1 0 16128 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_171
timestamp 1698431365
transform 1 0 20496 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_175
timestamp 1698431365
transform 1 0 20944 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_179
timestamp 1698431365
transform 1 0 21392 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_216
timestamp 1698431365
transform 1 0 25536 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_224
timestamp 1698431365
transform 1 0 26432 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_228
timestamp 1698431365
transform 1 0 26880 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_255
timestamp 1698431365
transform 1 0 29904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_259
timestamp 1698431365
transform 1 0 30352 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_275
timestamp 1698431365
transform 1 0 32144 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_279
timestamp 1698431365
transform 1 0 32592 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_290
timestamp 1698431365
transform 1 0 33824 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_294
timestamp 1698431365
transform 1 0 34272 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_296
timestamp 1698431365
transform 1 0 34496 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_303
timestamp 1698431365
transform 1 0 35280 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_307
timestamp 1698431365
transform 1 0 35728 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_311
timestamp 1698431365
transform 1 0 36176 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_313
timestamp 1698431365
transform 1 0 36400 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_343
timestamp 1698431365
transform 1 0 39760 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_347
timestamp 1698431365
transform 1 0 40208 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_349
timestamp 1698431365
transform 1 0 40432 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_352
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_356
timestamp 1698431365
transform 1 0 41216 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_416
timestamp 1698431365
transform 1 0 47936 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_480
timestamp 1698431365
transform 1 0 55104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_484
timestamp 1698431365
transform 1 0 55552 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_488
timestamp 1698431365
transform 1 0 56000 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_492
timestamp 1698431365
transform 1 0 56448 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_500
timestamp 1698431365
transform 1 0 57344 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_2
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_10
timestamp 1698431365
transform 1 0 2464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_12
timestamp 1698431365
transform 1 0 2688 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_17
timestamp 1698431365
transform 1 0 3248 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_33
timestamp 1698431365
transform 1 0 5040 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_40
timestamp 1698431365
transform 1 0 5824 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_48
timestamp 1698431365
transform 1 0 6720 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_53
timestamp 1698431365
transform 1 0 7280 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_61
timestamp 1698431365
transform 1 0 8176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_65
timestamp 1698431365
transform 1 0 8624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_67
timestamp 1698431365
transform 1 0 8848 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_74
timestamp 1698431365
transform 1 0 9632 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_82
timestamp 1698431365
transform 1 0 10528 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_84
timestamp 1698431365
transform 1 0 10752 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_89
timestamp 1698431365
transform 1 0 11312 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_97
timestamp 1698431365
transform 1 0 12208 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_101
timestamp 1698431365
transform 1 0 12656 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_108
timestamp 1698431365
transform 1 0 13440 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_116
timestamp 1698431365
transform 1 0 14336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_120
timestamp 1698431365
transform 1 0 14784 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_125
timestamp 1698431365
transform 1 0 15344 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_133
timestamp 1698431365
transform 1 0 16240 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_135
timestamp 1698431365
transform 1 0 16464 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_138
timestamp 1698431365
transform 1 0 16800 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_143
timestamp 1698431365
transform 1 0 17360 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_172
timestamp 1698431365
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_176
timestamp 1698431365
transform 1 0 21056 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_206
timestamp 1698431365
transform 1 0 24416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_210
timestamp 1698431365
transform 1 0 24864 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_237
timestamp 1698431365
transform 1 0 27888 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_240
timestamp 1698431365
transform 1 0 28224 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_244
timestamp 1698431365
transform 1 0 28672 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_246
timestamp 1698431365
transform 1 0 28896 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_251
timestamp 1698431365
transform 1 0 29456 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_259
timestamp 1698431365
transform 1 0 30352 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_263
timestamp 1698431365
transform 1 0 30800 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_269
timestamp 1698431365
transform 1 0 31472 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_271
timestamp 1698431365
transform 1 0 31696 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_274
timestamp 1698431365
transform 1 0 32032 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_282
timestamp 1698431365
transform 1 0 32928 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_287
timestamp 1698431365
transform 1 0 33488 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_295
timestamp 1698431365
transform 1 0 34384 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_299
timestamp 1698431365
transform 1 0 34832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_305
timestamp 1698431365
transform 1 0 35504 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_308
timestamp 1698431365
transform 1 0 35840 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_312
timestamp 1698431365
transform 1 0 36288 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_368
timestamp 1698431365
transform 1 0 42560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_402
timestamp 1698431365
transform 1 0 46368 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_406
timestamp 1698431365
transform 1 0 46816 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_436
timestamp 1698431365
transform 1 0 50176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_440
timestamp 1698431365
transform 1 0 50624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_470
timestamp 1698431365
transform 1 0 53984 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_474
timestamp 1698431365
transform 1 0 54432 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_504
timestamp 1698431365
transform 1 0 57792 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_508
timestamp 1698431365
transform 1 0 58240 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform -1 0 58352 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 58352 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform -1 0 58352 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 58352 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform -1 0 58352 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 58352 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 58352 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1698431365
transform -1 0 58352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1698431365
transform -1 0 58352 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform -1 0 58352 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input12
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform -1 0 24192 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform 1 0 24976 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform -1 0 29904 0 -1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform -1 0 39424 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 39648 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 41552 0 1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform -1 0 46368 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 47264 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform -1 0 50064 0 1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 51072 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 51184 0 -1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 54880 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 55216 0 1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 53312 0 -1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform 1 0 17472 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_81 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_110
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_111
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_112
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_113
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_114
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_115
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_116
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_117
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_118
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_119
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_120
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_121
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_122
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_123
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_124
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_125
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_126
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_127
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_128
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_129
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_130
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_131
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_132
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_133
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_134
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_135
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_136
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_137
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_138
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_139
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_140
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_141
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_142
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_143
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_144
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_145
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_146
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_147
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_148
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_149
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 58576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_150
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 58576 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_151
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 58576 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_152
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 58576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_153
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 58576 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_154
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 58576 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_155
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 58576 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_156
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 58576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_157
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 58576 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_158
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 58576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_159
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 58576 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_160
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 58576 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_161
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 58576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer1
timestamp 1698431365
transform 1 0 13664 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer2
timestamp 1698431365
transform 1 0 19152 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer3
timestamp 1698431365
transform -1 0 21840 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer4
timestamp 1698431365
transform -1 0 54880 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer5
timestamp 1698431365
transform 1 0 56448 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer6
timestamp 1698431365
transform -1 0 17248 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer7
timestamp 1698431365
transform 1 0 11424 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer8
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer9
timestamp 1698431365
transform -1 0 41104 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer10
timestamp 1698431365
transform -1 0 12880 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer11
timestamp 1698431365
transform -1 0 6720 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer12
timestamp 1698431365
transform -1 0 21840 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer13
timestamp 1698431365
transform -1 0 16016 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer14
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer15
timestamp 1698431365
transform 1 0 37520 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer16
timestamp 1698431365
transform -1 0 28560 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer17
timestamp 1698431365
transform -1 0 12880 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  rebuffer18
timestamp 1698431365
transform 1 0 18480 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer19 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer20
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_162 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_163
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_164
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_165
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_166
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_167
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_168
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_169
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_170
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_171
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_172
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_173
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_174
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_175
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_176
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_177
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_178
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_179
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_180
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_181
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_182
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_183
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_184
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_185
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_186
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_187
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_188
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_189
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_190
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_191
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_192
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_193
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_194
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_195
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_196
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_197
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_198
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_199
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_200
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_201
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_202
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_203
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_204
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_205
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_206
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_207
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_208
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_209
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_210
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_211
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_212
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_213
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_214
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_215
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_216
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_217
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_218
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_219
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_220
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_221
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_222
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_223
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_224
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_225
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_226
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_227
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_228
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_229
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_230
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_231
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_232
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_233
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_234
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_235
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_236
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_237
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_238
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_239
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_240
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_241
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_242
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_243
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_244
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_245
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_246
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_247
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_248
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_249
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_250
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_251
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_252
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_253
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_254
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_255
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_256
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_257
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_258
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_259
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_260
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_261
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_262
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_263
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_264
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_265
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_266
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_267
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_268
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_269
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_270
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_271
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_272
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_273
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_274
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_275
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_276
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_277
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_278
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_279
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_280
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_281
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_282
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_283
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_284
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_285
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_286
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_287
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_288
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_289
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_290
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_291
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_292
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_293
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_294
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_295
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_296
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_297
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_298
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_299
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_300
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_301
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_302
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_303
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_304
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_305
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_306
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_307
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_308
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_309
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_310
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_311
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_312
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_313
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_314
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_315
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_316
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_317
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_318
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_319
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_320
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_321
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_322
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_323
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_324
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_325
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_326
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_327
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_328
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_329
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_330
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_331
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_332
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_333
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_334
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_335
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_336
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_337
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_338
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_339
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_340
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_341
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_342
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_343
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_344
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_345
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_346
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_347
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_348
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_349
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_350
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_351
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_352
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_353
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_354
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_355
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_356
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_357
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_358
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_359
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_360
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_361
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_362
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_363
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_364
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_365
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_366
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_367
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_368
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_369
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_370
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_371
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_372
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_373
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_374
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_375
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_376
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_377
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_378
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_379
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_380
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_381
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_382
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_383
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_384
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_385
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_386
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_387
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_388
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_389
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_390
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_391
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_392
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_393
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_394
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_395
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_396
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_397
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_398
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_399
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_400
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_401
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_402
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_403
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_404
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_405
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_406
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_407
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_408
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_409
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_410
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_411
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_412
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_413
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_414
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_415
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_416
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_417
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_418
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_419
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_420
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_421
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_422
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_423
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_424
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_425
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_426
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_427
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_428
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_429
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_430
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_431
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_432
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_433
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_434
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_435
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_436
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_437
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_438
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_439
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_440
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_441
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_442
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_443
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_444
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_445
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_446
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_447
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_448
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_449
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_450
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_451
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_452
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_453
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_454
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_455
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_456
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_457
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_458
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_459
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_460
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_461
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_462
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_463
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_464
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_465
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_466
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_467
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_468
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_469
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_470
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_471
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_472
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_473
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_474
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_475
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_476
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_477
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_478
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_479
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_480
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_481
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_482
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_483
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_484
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_485
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_486
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_487
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_488
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_489
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_490
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_491
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_492
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_493
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_494
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_495
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_496
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_497
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_498
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_499
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_500
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_501
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_502
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_503
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_504
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_505
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_506
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_507
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_508
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_509
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_510
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_511
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_512
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_513
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_514
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_515
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_516
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_517
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_518
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_519
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_520
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_521
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_522
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_523
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_524
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_525
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_526
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_527
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_528
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_529
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_530
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_531
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_532
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_533
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_534
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_535
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_536
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_537
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_538
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_539
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_540
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_541
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_542
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_543
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_544
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_545
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_546
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_547
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_548
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_549
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_550
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_551
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_552
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_553
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_554
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_555
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_556
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_557
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_558
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_559
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_560
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_561
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_562
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_563
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_564
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_565
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_566
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_567
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_568
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_569
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_570
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_571
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_572
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_573
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_574
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_575
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_576
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_577
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_578
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_579
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_580
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_581
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_582
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_583
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_584
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_585
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_586
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_587
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_588
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_589
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_590
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_591
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_592
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_593
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_594
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_595
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_596
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_597
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_598
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_599
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_600
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_601
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_602
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_603
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_604
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_605
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_606
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_607
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_608
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_609
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_610
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_611
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_612
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_613
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_614
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_615
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_616
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_617
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_618
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_619
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_620
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_621
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_622
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_623
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_624
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_625
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_626
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_627
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_628
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_629
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_630
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_631
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_632
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_633
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_634
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_635
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_636
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_637
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_638
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_639
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_640
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_641
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_642
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_643
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_644
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_645
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_646
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_647
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_648
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_649
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_650
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_651
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_652
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_653
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_654
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_655
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_656
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_657
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_658
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_659
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_660
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_661
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_662
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_663
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_664
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_665
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_666
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_667
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_668
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_669
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_670
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_671
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_672
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_673
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_674
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_675
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_676
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_677
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_678
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_679
timestamp 1698431365
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_680
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_681
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_682
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_683
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_684
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_685
timestamp 1698431365
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_686
timestamp 1698431365
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_687
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_688
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_689
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_690
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_691
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_692
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_693
timestamp 1698431365
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_694
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_695
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_696
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_697
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_698
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_699
timestamp 1698431365
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_700
timestamp 1698431365
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_701
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_702
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_703
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_704
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_705
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_706
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_707
timestamp 1698431365
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_708
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_709
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_710
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_711
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_712
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_713
timestamp 1698431365
transform 1 0 48384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_714
timestamp 1698431365
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_715
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_716
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_717
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_718
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_719
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_720
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_721
timestamp 1698431365
transform 1 0 52304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_722
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_723
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_724
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_725
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_726
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_727
timestamp 1698431365
transform 1 0 48384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_728
timestamp 1698431365
transform 1 0 56224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_729
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_730
timestamp 1698431365
transform 1 0 8960 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_731
timestamp 1698431365
transform 1 0 12768 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_732
timestamp 1698431365
transform 1 0 16576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_733
timestamp 1698431365
transform 1 0 20384 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_734
timestamp 1698431365
transform 1 0 24192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_735
timestamp 1698431365
transform 1 0 28000 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_736
timestamp 1698431365
transform 1 0 31808 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_737
timestamp 1698431365
transform 1 0 35616 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_738
timestamp 1698431365
transform 1 0 39424 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_739
timestamp 1698431365
transform 1 0 43232 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_740
timestamp 1698431365
transform 1 0 47040 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_741
timestamp 1698431365
transform 1 0 50848 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_742
timestamp 1698431365
transform 1 0 54656 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_29 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3248 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_30
timestamp 1698431365
transform -1 0 5824 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_31
timestamp 1698431365
transform -1 0 7280 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_32
timestamp 1698431365
transform -1 0 9632 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_33
timestamp 1698431365
transform -1 0 11312 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_34
timestamp 1698431365
transform -1 0 13440 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_35
timestamp 1698431365
transform -1 0 15344 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_36
timestamp 1698431365
transform -1 0 17360 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_37
timestamp 1698431365
transform -1 0 29456 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_38
timestamp 1698431365
transform -1 0 31472 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_39
timestamp 1698431365
transform -1 0 33488 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_40
timestamp 1698431365
transform -1 0 35504 0 1 65856
box -86 -86 534 870
<< labels >>
flabel metal3 s 59200 59136 60000 59248 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 59200 66080 60000 66192 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 59200 3584 60000 3696 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 59200 10528 60000 10640 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 59200 17472 60000 17584 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 59200 24416 60000 24528 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 59200 31360 60000 31472 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 59200 38304 60000 38416 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 59200 45248 60000 45360 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 59200 52192 60000 52304 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal3 s 0 58240 800 58352 0 FreeSans 448 0 0 0 io_in_2
port 10 nsew signal input
flabel metal2 s 2688 69200 2800 70000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal tristate
flabel metal2 s 22848 69200 22960 70000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal tristate
flabel metal2 s 24864 69200 24976 70000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal tristate
flabel metal2 s 26880 69200 26992 70000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal tristate
flabel metal2 s 28896 69200 29008 70000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal tristate
flabel metal2 s 30912 69200 31024 70000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal tristate
flabel metal2 s 32928 69200 33040 70000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal tristate
flabel metal2 s 34944 69200 35056 70000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal tristate
flabel metal2 s 36960 69200 37072 70000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal tristate
flabel metal2 s 38976 69200 39088 70000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal tristate
flabel metal2 s 40992 69200 41104 70000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal tristate
flabel metal2 s 4704 69200 4816 70000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal tristate
flabel metal2 s 43008 69200 43120 70000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal tristate
flabel metal2 s 45024 69200 45136 70000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal tristate
flabel metal2 s 47040 69200 47152 70000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal tristate
flabel metal2 s 49056 69200 49168 70000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal tristate
flabel metal2 s 51072 69200 51184 70000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal tristate
flabel metal2 s 53088 69200 53200 70000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal tristate
flabel metal2 s 55104 69200 55216 70000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal tristate
flabel metal2 s 57120 69200 57232 70000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal tristate
flabel metal2 s 6720 69200 6832 70000 0 FreeSans 448 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 8736 69200 8848 70000 0 FreeSans 448 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 10752 69200 10864 70000 0 FreeSans 448 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 12768 69200 12880 70000 0 FreeSans 448 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 14784 69200 14896 70000 0 FreeSans 448 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 16800 69200 16912 70000 0 FreeSans 448 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 18816 69200 18928 70000 0 FreeSans 448 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 20832 69200 20944 70000 0 FreeSans 448 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 rst_n
port 39 nsew signal input
flabel metal4 s 4448 3076 4768 66700 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 35168 3076 35488 66700 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 19808 3076 20128 66700 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 66700 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal3 s 0 11648 800 11760 0 FreeSans 448 0 0 0 wb_clk_i
port 42 nsew signal input
rlabel metal1 29960 66640 29960 66640 0 vdd
rlabel metal1 29960 65856 29960 65856 0 vss
rlabel metal2 47600 64344 47600 64344 0 _0000_
rlabel metal2 29736 10192 29736 10192 0 _0001_
rlabel metal2 29848 7784 29848 7784 0 _0002_
rlabel metal2 31080 5152 31080 5152 0 _0003_
rlabel metal2 31472 4424 31472 4424 0 _0004_
rlabel metal2 47768 5488 47768 5488 0 _0005_
rlabel metal2 45416 8624 45416 8624 0 _0006_
rlabel metal2 45080 4424 45080 4424 0 _0007_
rlabel metal2 43736 6048 43736 6048 0 _0008_
rlabel metal2 47544 22288 47544 22288 0 _0009_
rlabel metal2 47880 19600 47880 19600 0 _0010_
rlabel metal2 45864 18760 45864 18760 0 _0011_
rlabel metal2 45864 22736 45864 22736 0 _0012_
rlabel metal2 41160 40824 41160 40824 0 _0013_
rlabel metal2 41272 36904 41272 36904 0 _0014_
rlabel metal3 21056 43400 21056 43400 0 _0015_
rlabel metal2 23688 49392 23688 49392 0 _0016_
rlabel metal3 18816 48888 18816 48888 0 _0017_
rlabel metal2 18200 53256 18200 53256 0 _0018_
rlabel metal2 21336 53032 21336 53032 0 _0019_
rlabel metal2 22120 57288 22120 57288 0 _0020_
rlabel metal2 22624 60200 22624 60200 0 _0021_
rlabel metal2 17864 56336 17864 56336 0 _0022_
rlabel metal2 20552 59248 20552 59248 0 _0023_
rlabel metal2 2520 36680 2520 36680 0 _0024_
rlabel metal2 2520 40880 2520 40880 0 _0025_
rlabel metal2 2632 44072 2632 44072 0 _0026_
rlabel metal2 2632 47096 2632 47096 0 _0027_
rlabel metal2 2520 50232 2520 50232 0 _0028_
rlabel metal2 2520 54656 2520 54656 0 _0029_
rlabel metal2 2520 57960 2520 57960 0 _0030_
rlabel metal3 5600 59416 5600 59416 0 _0031_
rlabel metal2 6664 63896 6664 63896 0 _0032_
rlabel metal2 21000 61320 21000 61320 0 _0033_
rlabel metal2 19656 63952 19656 63952 0 _0034_
rlabel metal2 5320 37464 5320 37464 0 _0035_
rlabel metal3 7448 41832 7448 41832 0 _0036_
rlabel metal2 7336 44688 7336 44688 0 _0037_
rlabel metal2 12152 46256 12152 46256 0 _0038_
rlabel metal3 8064 48888 8064 48888 0 _0039_
rlabel metal2 5992 53256 5992 53256 0 _0040_
rlabel metal2 7448 57064 7448 57064 0 _0041_
rlabel metal3 10472 60088 10472 60088 0 _0042_
rlabel metal3 11200 63336 11200 63336 0 _0043_
rlabel metal2 14952 63168 14952 63168 0 _0044_
rlabel metal2 17640 64736 17640 64736 0 _0045_
rlabel metal2 54264 39088 54264 39088 0 _0046_
rlabel metal2 53592 47096 53592 47096 0 _0047_
rlabel metal2 57176 45472 57176 45472 0 _0048_
rlabel metal2 53816 42112 53816 42112 0 _0049_
rlabel metal2 50848 45192 50848 45192 0 _0050_
rlabel metal2 50568 41328 50568 41328 0 _0051_
rlabel metal2 51016 39312 51016 39312 0 _0052_
rlabel metal3 48496 31640 48496 31640 0 _0053_
rlabel metal2 49112 29848 49112 29848 0 _0054_
rlabel metal3 52472 26936 52472 26936 0 _0055_
rlabel metal2 50232 25032 50232 25032 0 _0056_
rlabel metal2 51464 23464 51464 23464 0 _0057_
rlabel metal2 54376 21728 54376 21728 0 _0058_
rlabel metal2 56056 20944 56056 20944 0 _0059_
rlabel metal2 57288 24472 57288 24472 0 _0060_
rlabel metal3 56560 26488 56560 26488 0 _0061_
rlabel metal2 56056 30744 56056 30744 0 _0062_
rlabel metal2 56112 31864 56112 31864 0 _0063_
rlabel metal2 56728 35896 56728 35896 0 _0064_
rlabel metal2 55160 36120 55160 36120 0 _0065_
rlabel metal3 52752 33208 52752 33208 0 _0066_
rlabel metal2 49112 32984 49112 32984 0 _0067_
rlabel metal2 49112 25816 49112 25816 0 _0068_
rlabel metal2 43288 25928 43288 25928 0 _0069_
rlabel metal2 41832 28560 41832 28560 0 _0070_
rlabel metal2 43064 31696 43064 31696 0 _0071_
rlabel metal2 39592 32088 39592 32088 0 _0072_
rlabel metal2 44856 35840 44856 35840 0 _0073_
rlabel metal2 47320 34160 47320 34160 0 _0074_
rlabel metal2 46536 37688 46536 37688 0 _0075_
rlabel metal2 45976 40880 45976 40880 0 _0076_
rlabel metal2 33992 44520 33992 44520 0 _0077_
rlabel metal3 32648 45752 32648 45752 0 _0078_
rlabel metal3 28448 50456 28448 50456 0 _0079_
rlabel metal2 26040 53984 26040 53984 0 _0080_
rlabel metal3 33096 56952 33096 56952 0 _0081_
rlabel metal3 25536 63224 25536 63224 0 _0082_
rlabel metal2 29064 63168 29064 63168 0 _0083_
rlabel metal2 35672 65072 35672 65072 0 _0084_
rlabel metal3 23072 64904 23072 64904 0 _0085_
rlabel metal3 53256 11480 53256 11480 0 _0086_
rlabel metal2 56504 17976 56504 17976 0 _0087_
rlabel metal2 57400 16464 57400 16464 0 _0088_
rlabel metal3 55384 14392 55384 14392 0 _0089_
rlabel metal3 54040 13832 54040 13832 0 _0090_
rlabel metal3 48384 11480 48384 11480 0 _0091_
rlabel metal2 43960 11312 43960 11312 0 _0092_
rlabel metal2 42616 15148 42616 15148 0 _0093_
rlabel metal2 40208 11480 40208 11480 0 _0094_
rlabel metal2 38584 22288 38584 22288 0 _0095_
rlabel metal2 27944 33712 27944 33712 0 _0096_
rlabel metal3 53256 9688 53256 9688 0 _0097_
rlabel metal3 53704 6664 53704 6664 0 _0098_
rlabel metal2 52696 4648 52696 4648 0 _0099_
rlabel metal3 41272 4424 41272 4424 0 _0100_
rlabel metal2 38248 4816 38248 4816 0 _0101_
rlabel metal2 36456 5040 36456 5040 0 _0102_
rlabel metal2 33544 5432 33544 5432 0 _0103_
rlabel metal2 30296 12880 30296 12880 0 _0104_
rlabel metal2 36008 12376 36008 12376 0 _0105_
rlabel metal2 35672 15792 35672 15792 0 _0106_
rlabel metal2 7896 25704 7896 25704 0 _0107_
rlabel metal2 26824 11032 26824 11032 0 _0108_
rlabel metal2 26040 4648 26040 4648 0 _0109_
rlabel metal2 22344 4648 22344 4648 0 _0110_
rlabel metal2 19096 4648 19096 4648 0 _0111_
rlabel metal2 17416 6328 17416 6328 0 _0112_
rlabel metal2 15736 9464 15736 9464 0 _0113_
rlabel metal2 15736 11032 15736 11032 0 _0114_
rlabel metal2 14728 13888 14728 13888 0 _0115_
rlabel metal2 23800 11144 23800 11144 0 _0116_
rlabel metal2 24472 14616 24472 14616 0 _0117_
rlabel metal2 18648 32984 18648 32984 0 _0118_
rlabel metal2 46648 43876 46648 43876 0 _0119_
rlabel metal2 41496 43932 41496 43932 0 _0120_
rlabel metal2 45528 45640 45528 45640 0 _0121_
rlabel metal2 39592 46200 39592 46200 0 _0122_
rlabel metal2 40712 50904 40712 50904 0 _0123_
rlabel metal2 39592 54936 39592 54936 0 _0124_
rlabel metal3 46144 58520 46144 58520 0 _0125_
rlabel metal2 39256 58800 39256 58800 0 _0126_
rlabel metal2 43624 64512 43624 64512 0 _0127_
rlabel metal2 46144 62216 46144 62216 0 _0128_
rlabel metal2 57400 63448 57400 63448 0 _0129_
rlabel metal2 56840 59640 56840 59640 0 _0130_
rlabel metal2 57064 61880 57064 61880 0 _0131_
rlabel metal3 52528 54712 52528 54712 0 _0132_
rlabel metal2 55944 48664 55944 48664 0 _0133_
rlabel metal2 56056 51296 56056 51296 0 _0134_
rlabel metal2 55384 55412 55384 55412 0 _0135_
rlabel metal2 56000 53816 56000 53816 0 _0136_
rlabel metal2 51240 52640 51240 52640 0 _0137_
rlabel metal2 53032 48552 53032 48552 0 _0138_
rlabel metal2 48888 49336 48888 49336 0 _0139_
rlabel metal2 44968 50960 44968 50960 0 _0140_
rlabel metal2 48888 51800 48888 51800 0 _0141_
rlabel metal2 43288 52528 43288 52528 0 _0142_
rlabel metal2 45640 55608 45640 55608 0 _0143_
rlabel metal2 48888 56504 48888 56504 0 _0144_
rlabel metal2 48104 59640 48104 59640 0 _0145_
rlabel metal2 49392 62216 49392 62216 0 _0146_
rlabel metal2 50232 65128 50232 65128 0 _0147_
rlabel metal2 51800 65128 51800 65128 0 _0148_
rlabel metal2 52136 58856 52136 58856 0 _0149_
rlabel metal2 51632 56168 51632 56168 0 _0150_
rlabel metal2 50456 36120 50456 36120 0 _0151_
rlabel metal2 41496 22008 41496 22008 0 _0152_
rlabel metal3 41832 19880 41832 19880 0 _0153_
rlabel metal2 42224 17752 42224 17752 0 _0154_
rlabel metal2 38528 17752 38528 17752 0 _0155_
rlabel metal2 36008 18480 36008 18480 0 _0156_
rlabel metal2 34440 22008 34440 22008 0 _0157_
rlabel metal2 27384 15456 27384 15456 0 _0158_
rlabel metal2 28000 16744 28000 16744 0 _0159_
rlabel metal2 28616 20160 28616 20160 0 _0160_
rlabel metal2 26040 18592 26040 18592 0 _0161_
rlabel metal2 30408 17024 30408 17024 0 _0162_
rlabel metal2 31360 20216 31360 20216 0 _0163_
rlabel metal2 16744 16576 16744 16576 0 _0164_
rlabel metal2 14728 17192 14728 17192 0 _0165_
rlabel metal3 17248 20664 17248 20664 0 _0166_
rlabel metal2 15064 18760 15064 18760 0 _0167_
rlabel metal2 20664 17024 20664 17024 0 _0168_
rlabel metal2 20272 20104 20272 20104 0 _0169_
rlabel metal2 31752 27440 31752 27440 0 _0170_
rlabel metal2 31920 28728 31920 28728 0 _0171_
rlabel metal2 29176 30576 29176 30576 0 _0172_
rlabel metal2 26488 29680 26488 29680 0 _0173_
rlabel metal2 25032 30968 25032 30968 0 _0174_
rlabel metal2 21728 30296 21728 30296 0 _0175_
rlabel metal4 22120 31976 22120 31976 0 _0176_
rlabel metal2 20328 28280 20328 28280 0 _0177_
rlabel metal2 5096 29120 5096 29120 0 _0178_
rlabel metal2 13384 28224 13384 28224 0 _0179_
rlabel metal2 13944 25480 13944 25480 0 _0180_
rlabel metal3 12656 24584 12656 24584 0 _0181_
rlabel metal2 16128 30296 16128 30296 0 _0182_
rlabel metal2 17752 24976 17752 24976 0 _0183_
rlabel metal3 17696 28392 17696 28392 0 _0184_
rlabel metal2 15960 24416 15960 24416 0 _0185_
rlabel metal2 20552 24864 20552 24864 0 _0186_
rlabel metal2 22512 21672 22512 21672 0 _0187_
rlabel metal2 30072 23464 30072 23464 0 _0188_
rlabel metal3 43960 26376 43960 26376 0 _0189_
rlabel metal2 36120 25032 36120 25032 0 _0190_
rlabel metal2 37240 29848 37240 29848 0 _0191_
rlabel metal2 39480 28112 39480 28112 0 _0192_
rlabel metal2 8624 56280 8624 56280 0 _0193_
rlabel metal2 47656 46760 47656 46760 0 _0194_
rlabel metal2 10248 56840 10248 56840 0 _0195_
rlabel metal2 10472 56560 10472 56560 0 _0196_
rlabel metal2 11816 58352 11816 58352 0 _0197_
rlabel metal2 12376 58968 12376 58968 0 _0198_
rlabel metal2 11144 60704 11144 60704 0 _0199_
rlabel metal2 12824 60872 12824 60872 0 _0200_
rlabel metal2 13160 61544 13160 61544 0 _0201_
rlabel metal2 12712 63728 12712 63728 0 _0202_
rlabel metal3 12544 64456 12544 64456 0 _0203_
rlabel metal2 12936 63392 12936 63392 0 _0204_
rlabel metal2 13832 62832 13832 62832 0 _0205_
rlabel metal3 16408 63112 16408 63112 0 _0206_
rlabel metal2 14840 62720 14840 62720 0 _0207_
rlabel metal2 16744 63280 16744 63280 0 _0208_
rlabel metal3 41160 32648 41160 32648 0 _0209_
rlabel metal2 28840 49896 28840 49896 0 _0210_
rlabel metal2 17528 63336 17528 63336 0 _0211_
rlabel metal2 55048 45976 55048 45976 0 _0212_
rlabel metal3 52528 11368 52528 11368 0 _0213_
rlabel metal2 53928 46648 53928 46648 0 _0214_
rlabel metal2 51240 46536 51240 46536 0 _0215_
rlabel metal2 56840 45192 56840 45192 0 _0216_
rlabel metal3 54936 44520 54936 44520 0 _0217_
rlabel metal2 53984 44408 53984 44408 0 _0218_
rlabel metal3 54264 43736 54264 43736 0 _0219_
rlabel metal2 50680 46088 50680 46088 0 _0220_
rlabel metal2 51240 45136 51240 45136 0 _0221_
rlabel metal2 50736 40936 50736 40936 0 _0222_
rlabel metal3 48440 48104 48440 48104 0 _0223_
rlabel metal2 49672 48160 49672 48160 0 _0224_
rlabel metal2 51688 42728 51688 42728 0 _0225_
rlabel metal2 50344 42168 50344 42168 0 _0226_
rlabel metal2 51352 40040 51352 40040 0 _0227_
rlabel metal2 39144 33992 39144 33992 0 _0228_
rlabel metal2 50344 35112 50344 35112 0 _0229_
rlabel metal2 53256 35168 53256 35168 0 _0230_
rlabel metal2 53200 29624 53200 29624 0 _0231_
rlabel metal2 50232 30352 50232 30352 0 _0232_
rlabel metal2 49896 31416 49896 31416 0 _0233_
rlabel metal2 55160 29736 55160 29736 0 _0234_
rlabel metal2 50120 31808 50120 31808 0 _0235_
rlabel metal2 51240 29680 51240 29680 0 _0236_
rlabel metal2 52192 32648 52192 32648 0 _0237_
rlabel metal3 53536 24696 53536 24696 0 _0238_
rlabel metal2 53256 29008 53256 29008 0 _0239_
rlabel metal2 53256 25312 53256 25312 0 _0240_
rlabel metal2 53816 24696 53816 24696 0 _0241_
rlabel metal2 53032 26908 53032 26908 0 _0242_
rlabel metal2 52360 26684 52360 26684 0 _0243_
rlabel metal2 53032 25536 53032 25536 0 _0244_
rlabel metal2 52584 25200 52584 25200 0 _0245_
rlabel metal3 53200 23800 53200 23800 0 _0246_
rlabel metal3 53872 23912 53872 23912 0 _0247_
rlabel metal2 54936 22792 54936 22792 0 _0248_
rlabel metal2 56784 25480 56784 25480 0 _0249_
rlabel metal3 55832 22232 55832 22232 0 _0250_
rlabel metal2 57176 21840 57176 21840 0 _0251_
rlabel metal3 57288 23240 57288 23240 0 _0252_
rlabel metal2 56952 21896 56952 21896 0 _0253_
rlabel metal2 56504 21840 56504 21840 0 _0254_
rlabel metal2 56952 24024 56952 24024 0 _0255_
rlabel metal2 56448 24696 56448 24696 0 _0256_
rlabel metal3 57456 27608 57456 27608 0 _0257_
rlabel metal2 57344 26264 57344 26264 0 _0258_
rlabel metal2 56728 30296 56728 30296 0 _0259_
rlabel metal2 55048 33432 55048 33432 0 _0260_
rlabel metal2 57288 32256 57288 32256 0 _0261_
rlabel metal3 56000 30968 56000 30968 0 _0262_
rlabel metal2 55832 34720 55832 34720 0 _0263_
rlabel metal2 57064 33824 57064 33824 0 _0264_
rlabel metal2 56728 34440 56728 34440 0 _0265_
rlabel metal3 57512 35672 57512 35672 0 _0266_
rlabel metal2 56616 35280 56616 35280 0 _0267_
rlabel metal2 55440 34888 55440 34888 0 _0268_
rlabel metal2 54712 35000 54712 35000 0 _0269_
rlabel metal2 53872 32312 53872 32312 0 _0270_
rlabel metal2 51800 32816 51800 32816 0 _0271_
rlabel metal2 46536 31416 46536 31416 0 _0272_
rlabel metal3 48216 32536 48216 32536 0 _0273_
rlabel metal3 50064 32536 50064 32536 0 _0274_
rlabel metal2 57624 40320 57624 40320 0 _0275_
rlabel metal3 56336 40488 56336 40488 0 _0276_
rlabel metal2 57064 40096 57064 40096 0 _0277_
rlabel metal2 55720 40880 55720 40880 0 _0278_
rlabel metal2 55384 41440 55384 41440 0 _0279_
rlabel metal2 51464 12544 51464 12544 0 _0280_
rlabel metal2 24248 12488 24248 12488 0 _0281_
rlabel metal3 46984 25480 46984 25480 0 _0282_
rlabel metal2 50120 46480 50120 46480 0 _0283_
rlabel metal2 57512 41104 57512 41104 0 _0284_
rlabel metal2 56952 40320 56952 40320 0 _0285_
rlabel metal3 24752 14392 24752 14392 0 _0286_
rlabel metal2 24360 14112 24360 14112 0 _0287_
rlabel metal2 43064 9968 43064 9968 0 _0288_
rlabel metal2 26096 10808 26096 10808 0 _0289_
rlabel metal3 44464 25704 44464 25704 0 _0290_
rlabel metal3 44744 26936 44744 26936 0 _0291_
rlabel metal2 44128 26824 44128 26824 0 _0292_
rlabel metal2 44016 31976 44016 31976 0 _0293_
rlabel metal2 43456 28728 43456 28728 0 _0294_
rlabel metal2 43904 33320 43904 33320 0 _0295_
rlabel metal2 43736 33768 43736 33768 0 _0296_
rlabel metal3 44520 18368 44520 18368 0 _0297_
rlabel metal3 43848 32424 43848 32424 0 _0298_
rlabel metal2 44296 34608 44296 34608 0 _0299_
rlabel metal2 41664 33320 41664 33320 0 _0300_
rlabel metal2 44072 35224 44072 35224 0 _0301_
rlabel metal3 45192 34104 45192 34104 0 _0302_
rlabel metal2 44968 35728 44968 35728 0 _0303_
rlabel metal2 46816 33992 46816 33992 0 _0304_
rlabel metal2 45864 39144 45864 39144 0 _0305_
rlabel metal2 46424 37408 46424 37408 0 _0306_
rlabel metal2 43848 40264 43848 40264 0 _0307_
rlabel metal3 44688 39480 44688 39480 0 _0308_
rlabel metal2 45304 40320 45304 40320 0 _0309_
rlabel metal2 44744 40096 44744 40096 0 _0310_
rlabel metal2 44688 41384 44688 41384 0 _0311_
rlabel metal3 39144 44072 39144 44072 0 _0312_
rlabel metal2 33656 44240 33656 44240 0 _0313_
rlabel metal2 34552 44296 34552 44296 0 _0314_
rlabel metal2 32536 47264 32536 47264 0 _0315_
rlabel metal2 31752 44800 31752 44800 0 _0316_
rlabel metal2 32480 43736 32480 43736 0 _0317_
rlabel metal2 31192 46480 31192 46480 0 _0318_
rlabel metal2 31584 46536 31584 46536 0 _0319_
rlabel metal2 29512 46592 29512 46592 0 _0320_
rlabel metal2 29008 46648 29008 46648 0 _0321_
rlabel metal2 29288 47936 29288 47936 0 _0322_
rlabel metal2 28504 50204 28504 50204 0 _0323_
rlabel metal2 29568 50008 29568 50008 0 _0324_
rlabel metal3 30184 50792 30184 50792 0 _0325_
rlabel metal3 29288 49784 29288 49784 0 _0326_
rlabel metal2 30128 50008 30128 50008 0 _0327_
rlabel metal2 29400 54824 29400 54824 0 _0328_
rlabel metal3 26796 54600 26796 54600 0 _0329_
rlabel metal2 28224 47880 28224 47880 0 _0330_
rlabel metal2 27272 54376 27272 54376 0 _0331_
rlabel metal2 29736 54152 29736 54152 0 _0332_
rlabel metal2 29512 54992 29512 54992 0 _0333_
rlabel metal2 30184 57232 30184 57232 0 _0334_
rlabel metal2 31864 57512 31864 57512 0 _0335_
rlabel metal2 29960 57568 29960 57568 0 _0336_
rlabel metal2 30856 57512 30856 57512 0 _0337_
rlabel metal2 27272 62608 27272 62608 0 _0338_
rlabel metal2 27048 63336 27048 63336 0 _0339_
rlabel metal3 26936 63112 26936 63112 0 _0340_
rlabel metal2 27832 63448 27832 63448 0 _0341_
rlabel metal2 27440 64008 27440 64008 0 _0342_
rlabel metal3 29960 64680 29960 64680 0 _0343_
rlabel metal2 29512 62944 29512 62944 0 _0344_
rlabel metal2 29400 62832 29400 62832 0 _0345_
rlabel metal2 33096 63896 33096 63896 0 _0346_
rlabel metal2 32424 63504 32424 63504 0 _0347_
rlabel metal2 34664 64176 34664 64176 0 _0348_
rlabel metal2 35168 64008 35168 64008 0 _0349_
rlabel metal2 32200 63784 32200 63784 0 _0350_
rlabel metal2 32088 63560 32088 63560 0 _0351_
rlabel metal3 29288 63784 29288 63784 0 _0352_
rlabel metal2 22120 14056 22120 14056 0 _0353_
rlabel metal2 51912 11760 51912 11760 0 _0354_
rlabel metal2 20328 10808 20328 10808 0 _0355_
rlabel metal2 51688 16464 51688 16464 0 _0356_
rlabel metal2 47768 15736 47768 15736 0 _0357_
rlabel metal2 49336 16520 49336 16520 0 _0358_
rlabel metal2 50960 11368 50960 11368 0 _0359_
rlabel metal2 51464 11256 51464 11256 0 _0360_
rlabel metal2 51296 12152 51296 12152 0 _0361_
rlabel metal2 51744 14392 51744 14392 0 _0362_
rlabel metal2 51520 17864 51520 17864 0 _0363_
rlabel metal3 52976 18200 52976 18200 0 _0364_
rlabel metal2 24584 12936 24584 12936 0 _0365_
rlabel metal2 20216 12656 20216 12656 0 _0366_
rlabel metal3 51912 18424 51912 18424 0 _0367_
rlabel metal3 53872 18312 53872 18312 0 _0368_
rlabel metal2 52136 17472 52136 17472 0 _0369_
rlabel metal3 53480 17864 53480 17864 0 _0370_
rlabel metal2 52024 16912 52024 16912 0 _0371_
rlabel metal2 53480 17304 53480 17304 0 _0372_
rlabel metal3 46480 15848 46480 15848 0 _0373_
rlabel metal2 52696 15232 52696 15232 0 _0374_
rlabel metal2 51240 14896 51240 14896 0 _0375_
rlabel metal2 52640 14728 52640 14728 0 _0376_
rlabel metal3 52360 14280 52360 14280 0 _0377_
rlabel metal2 53872 14616 53872 14616 0 _0378_
rlabel metal2 50960 13720 50960 13720 0 _0379_
rlabel metal3 49168 14504 49168 14504 0 _0380_
rlabel metal2 50008 9016 50008 9016 0 _0381_
rlabel metal2 50848 13944 50848 13944 0 _0382_
rlabel metal3 52304 13720 52304 13720 0 _0383_
rlabel metal2 51184 7560 51184 7560 0 _0384_
rlabel metal2 47656 14504 47656 14504 0 _0385_
rlabel metal2 47544 13664 47544 13664 0 _0386_
rlabel metal2 48216 13216 48216 13216 0 _0387_
rlabel metal2 47768 12320 47768 12320 0 _0388_
rlabel metal2 45080 15624 45080 15624 0 _0389_
rlabel metal2 45192 15148 45192 15148 0 _0390_
rlabel metal2 44968 13384 44968 13384 0 _0391_
rlabel metal2 43064 14448 43064 14448 0 _0392_
rlabel metal2 44632 13160 44632 13160 0 _0393_
rlabel metal3 45192 12264 45192 12264 0 _0394_
rlabel metal2 42560 13720 42560 13720 0 _0395_
rlabel metal2 22456 12600 22456 12600 0 _0396_
rlabel metal2 41496 14840 41496 14840 0 _0397_
rlabel metal3 40264 14392 40264 14392 0 _0398_
rlabel metal2 41272 12152 41272 12152 0 _0399_
rlabel metal2 41496 14056 41496 14056 0 _0400_
rlabel metal2 39704 15148 39704 15148 0 _0401_
rlabel metal2 38976 15512 38976 15512 0 _0402_
rlabel metal2 51016 12040 51016 12040 0 _0403_
rlabel metal2 39256 12040 39256 12040 0 _0404_
rlabel metal2 39592 12264 39592 12264 0 _0405_
rlabel metal2 38136 23184 38136 23184 0 _0406_
rlabel metal2 38360 22288 38360 22288 0 _0407_
rlabel metal2 38136 21728 38136 21728 0 _0408_
rlabel metal2 28392 33488 28392 33488 0 _0409_
rlabel metal2 51800 10192 51800 10192 0 _0410_
rlabel metal2 49336 7952 49336 7952 0 _0411_
rlabel metal3 38472 9688 38472 9688 0 _0412_
rlabel metal2 39592 9408 39592 9408 0 _0413_
rlabel metal2 50792 8232 50792 8232 0 _0414_
rlabel metal2 51296 9800 51296 9800 0 _0415_
rlabel metal3 50848 8344 50848 8344 0 _0416_
rlabel metal2 50680 7504 50680 7504 0 _0417_
rlabel metal2 50344 8176 50344 8176 0 _0418_
rlabel metal2 50904 7448 50904 7448 0 _0419_
rlabel metal3 52024 7336 52024 7336 0 _0420_
rlabel metal3 49784 6720 49784 6720 0 _0421_
rlabel metal2 50456 6664 50456 6664 0 _0422_
rlabel metal2 50344 7056 50344 7056 0 _0423_
rlabel metal2 51184 5208 51184 5208 0 _0424_
rlabel via2 39368 7336 39368 7336 0 _0425_
rlabel metal3 39536 9128 39536 9128 0 _0426_
rlabel metal3 40768 7672 40768 7672 0 _0427_
rlabel metal3 39928 6888 39928 6888 0 _0428_
rlabel metal3 39984 7448 39984 7448 0 _0429_
rlabel metal2 40936 7336 40936 7336 0 _0430_
rlabel metal2 40712 5488 40712 5488 0 _0431_
rlabel metal2 37744 7448 37744 7448 0 _0432_
rlabel metal2 38808 6944 38808 6944 0 _0433_
rlabel metal2 38920 7056 38920 7056 0 _0434_
rlabel metal2 38136 5432 38136 5432 0 _0435_
rlabel metal2 35448 8456 35448 8456 0 _0436_
rlabel metal2 35000 7616 35000 7616 0 _0437_
rlabel metal2 36064 7448 36064 7448 0 _0438_
rlabel metal3 25256 6440 25256 6440 0 _0439_
rlabel metal2 35504 5992 35504 5992 0 _0440_
rlabel metal3 32760 15176 32760 15176 0 _0441_
rlabel metal2 33488 9128 33488 9128 0 _0442_
rlabel metal2 33712 7448 33712 7448 0 _0443_
rlabel metal2 32872 9464 32872 9464 0 _0444_
rlabel metal2 33488 7448 33488 7448 0 _0445_
rlabel metal2 33880 6272 33880 6272 0 _0446_
rlabel metal2 31640 11872 31640 11872 0 _0447_
rlabel metal3 32648 13048 32648 13048 0 _0448_
rlabel metal3 34888 13048 34888 13048 0 _0449_
rlabel metal2 32312 11760 32312 11760 0 _0450_
rlabel metal2 32648 11648 32648 11648 0 _0451_
rlabel metal2 34776 13664 34776 13664 0 _0452_
rlabel metal2 35000 14056 35000 14056 0 _0453_
rlabel metal2 34944 12264 34944 12264 0 _0454_
rlabel metal3 34888 12376 34888 12376 0 _0455_
rlabel metal2 41776 46536 41776 46536 0 _0456_
rlabel metal3 8036 25480 8036 25480 0 _0457_
rlabel metal2 34328 15512 34328 15512 0 _0458_
rlabel metal2 35336 15540 35336 15540 0 _0459_
rlabel metal2 46200 46200 46200 46200 0 _0460_
rlabel metal2 8232 25816 8232 25816 0 _0461_
rlabel metal2 27048 11424 27048 11424 0 _0462_
rlabel metal2 24808 8036 24808 8036 0 _0463_
rlabel metal2 19880 10024 19880 10024 0 _0464_
rlabel metal3 26040 8456 26040 8456 0 _0465_
rlabel metal2 26376 7728 26376 7728 0 _0466_
rlabel metal2 26600 10472 26600 10472 0 _0467_
rlabel metal3 23072 6664 23072 6664 0 _0468_
rlabel metal2 26768 7560 26768 7560 0 _0469_
rlabel metal2 23800 6832 23800 6832 0 _0470_
rlabel metal2 26824 7896 26824 7896 0 _0471_
rlabel metal2 25928 5992 25928 5992 0 _0472_
rlabel metal2 23576 5936 23576 5936 0 _0473_
rlabel metal2 21336 7168 21336 7168 0 _0474_
rlabel metal2 24192 5880 24192 5880 0 _0475_
rlabel metal2 23576 6104 23576 6104 0 _0476_
rlabel metal2 23240 5992 23240 5992 0 _0477_
rlabel metal2 21560 11032 21560 11032 0 _0478_
rlabel metal2 20776 6384 20776 6384 0 _0479_
rlabel metal2 21448 7056 21448 7056 0 _0480_
rlabel metal2 20664 6720 20664 6720 0 _0481_
rlabel metal2 20440 8008 20440 8008 0 _0482_
rlabel metal2 20216 5992 20216 5992 0 _0483_
rlabel metal2 19096 6776 19096 6776 0 _0484_
rlabel metal2 19152 5656 19152 5656 0 _0485_
rlabel metal2 19712 6888 19712 6888 0 _0486_
rlabel metal2 17584 5880 17584 5880 0 _0487_
rlabel metal2 18144 10024 18144 10024 0 _0488_
rlabel metal3 18648 12712 18648 12712 0 _0489_
rlabel metal2 18872 9184 18872 9184 0 _0490_
rlabel metal2 15848 9352 15848 9352 0 _0491_
rlabel metal2 21336 11368 21336 11368 0 _0492_
rlabel metal2 18984 13048 18984 13048 0 _0493_
rlabel metal2 19432 11480 19432 11480 0 _0494_
rlabel metal2 18312 13440 18312 13440 0 _0495_
rlabel metal2 19824 13160 19824 13160 0 _0496_
rlabel metal2 15848 10920 15848 10920 0 _0497_
rlabel metal2 20552 13440 20552 13440 0 _0498_
rlabel metal2 19208 13720 19208 13720 0 _0499_
rlabel metal2 21280 13160 21280 13160 0 _0500_
rlabel metal2 21448 13384 21448 13384 0 _0501_
rlabel metal3 20328 13720 20328 13720 0 _0502_
rlabel metal3 23016 13720 23016 13720 0 _0503_
rlabel metal2 24360 12936 24360 12936 0 _0504_
rlabel metal2 23016 12768 23016 12768 0 _0505_
rlabel metal2 24136 12880 24136 12880 0 _0506_
rlabel metal3 22120 16184 22120 16184 0 _0507_
rlabel metal2 23688 15512 23688 15512 0 _0508_
rlabel metal2 24248 15680 24248 15680 0 _0509_
rlabel metal2 19096 32872 19096 32872 0 _0510_
rlabel metal2 46536 44408 46536 44408 0 _0511_
rlabel metal2 46872 44408 46872 44408 0 _0512_
rlabel metal2 44184 42896 44184 42896 0 _0513_
rlabel metal2 34888 41496 34888 41496 0 _0514_
rlabel metal2 39368 42392 39368 42392 0 _0515_
rlabel metal2 43960 43932 43960 43932 0 _0516_
rlabel metal3 41888 42616 41888 42616 0 _0517_
rlabel metal2 43904 41720 43904 41720 0 _0518_
rlabel metal2 44520 44296 44520 44296 0 _0519_
rlabel metal2 45976 46928 45976 46928 0 _0520_
rlabel metal3 44100 46648 44100 46648 0 _0521_
rlabel metal3 45584 46648 45584 46648 0 _0522_
rlabel metal2 45080 46200 45080 46200 0 _0523_
rlabel metal2 42560 49000 42560 49000 0 _0524_
rlabel metal2 42392 48552 42392 48552 0 _0525_
rlabel metal2 42504 47712 42504 47712 0 _0526_
rlabel metal3 42784 49672 42784 49672 0 _0527_
rlabel metal2 41328 46760 41328 46760 0 _0528_
rlabel metal2 41944 49448 41944 49448 0 _0529_
rlabel metal2 41272 49672 41272 49672 0 _0530_
rlabel metal3 41608 50008 41608 50008 0 _0531_
rlabel metal3 41888 49784 41888 49784 0 _0532_
rlabel metal3 41440 50792 41440 50792 0 _0533_
rlabel metal2 41384 50092 41384 50092 0 _0534_
rlabel metal2 41272 51184 41272 51184 0 _0535_
rlabel metal2 41272 54152 41272 54152 0 _0536_
rlabel metal2 39984 53480 39984 53480 0 _0537_
rlabel metal3 40152 54600 40152 54600 0 _0538_
rlabel metal2 40656 45304 40656 45304 0 _0539_
rlabel metal2 40040 54152 40040 54152 0 _0540_
rlabel metal2 49448 49896 49448 49896 0 _0541_
rlabel metal2 42504 54768 42504 54768 0 _0542_
rlabel metal2 42728 57008 42728 57008 0 _0543_
rlabel metal2 42952 56392 42952 56392 0 _0544_
rlabel metal2 43624 57344 43624 57344 0 _0545_
rlabel metal2 44968 58408 44968 58408 0 _0546_
rlabel metal3 42728 59304 42728 59304 0 _0547_
rlabel metal2 42616 58744 42616 58744 0 _0548_
rlabel metal3 42280 59192 42280 59192 0 _0549_
rlabel metal3 40712 60536 40712 60536 0 _0550_
rlabel metal2 40824 59472 40824 59472 0 _0551_
rlabel metal2 41496 59640 41496 59640 0 _0552_
rlabel metal3 43820 62328 43820 62328 0 _0553_
rlabel metal3 42896 61432 42896 61432 0 _0554_
rlabel metal2 43008 62328 43008 62328 0 _0555_
rlabel metal2 42504 62272 42504 62272 0 _0556_
rlabel metal2 43288 63056 43288 63056 0 _0557_
rlabel metal2 45528 62664 45528 62664 0 _0558_
rlabel metal2 44744 62720 44744 62720 0 _0559_
rlabel metal2 44744 62328 44744 62328 0 _0560_
rlabel metal3 45360 62328 45360 62328 0 _0561_
rlabel metal2 46536 62440 46536 62440 0 _0562_
rlabel metal2 45192 63560 45192 63560 0 _0563_
rlabel metal2 47208 62608 47208 62608 0 _0564_
rlabel metal3 50680 64120 50680 64120 0 _0565_
rlabel metal2 55048 62664 55048 62664 0 _0566_
rlabel metal2 54656 63336 54656 63336 0 _0567_
rlabel metal2 53592 63616 53592 63616 0 _0568_
rlabel metal3 54712 63672 54712 63672 0 _0569_
rlabel metal2 56560 59192 56560 59192 0 _0570_
rlabel metal2 57176 61600 57176 61600 0 _0571_
rlabel metal3 57512 60536 57512 60536 0 _0572_
rlabel metal2 52864 51576 52864 51576 0 _0573_
rlabel metal2 51688 54208 51688 54208 0 _0574_
rlabel metal2 54712 48720 54712 48720 0 _0575_
rlabel metal2 54824 48552 54824 48552 0 _0576_
rlabel metal2 56728 51968 56728 51968 0 _0577_
rlabel metal2 55160 55720 55160 55720 0 _0578_
rlabel metal2 55608 56280 55608 56280 0 _0579_
rlabel metal2 56056 54320 56056 54320 0 _0580_
rlabel metal2 51016 50456 51016 50456 0 _0581_
rlabel metal2 53032 49280 53032 49280 0 _0582_
rlabel metal2 54488 53592 54488 53592 0 _0583_
rlabel metal2 53256 49896 53256 49896 0 _0584_
rlabel metal2 47656 50960 47656 50960 0 _0585_
rlabel metal2 47320 49952 47320 49952 0 _0586_
rlabel metal2 44968 47600 44968 47600 0 _0587_
rlabel metal2 45528 51408 45528 51408 0 _0588_
rlabel metal3 51688 53648 51688 53648 0 _0589_
rlabel metal2 51240 53984 51240 53984 0 _0590_
rlabel metal2 48776 51520 48776 51520 0 _0591_
rlabel metal2 43848 52472 43848 52472 0 _0592_
rlabel metal2 47208 55776 47208 55776 0 _0593_
rlabel metal2 46648 55328 46648 55328 0 _0594_
rlabel metal2 48776 56224 48776 56224 0 _0595_
rlabel metal2 51464 62104 51464 62104 0 _0596_
rlabel metal3 50232 63112 50232 63112 0 _0597_
rlabel metal3 48888 59304 48888 59304 0 _0598_
rlabel metal2 49672 61040 49672 61040 0 _0599_
rlabel metal2 50400 64120 50400 64120 0 _0600_
rlabel metal2 51688 63896 51688 63896 0 _0601_
rlabel metal2 52024 59136 52024 59136 0 _0602_
rlabel metal3 52416 56504 52416 56504 0 _0603_
rlabel metal2 31360 24920 31360 24920 0 _0604_
rlabel metal2 18648 16856 18648 16856 0 _0605_
rlabel metal2 24136 22680 24136 22680 0 _0606_
rlabel metal2 24920 23744 24920 23744 0 _0607_
rlabel metal2 24584 25648 24584 25648 0 _0608_
rlabel metal2 25424 22232 25424 22232 0 _0609_
rlabel metal3 31080 21784 31080 21784 0 _0610_
rlabel metal2 40936 19264 40936 19264 0 _0611_
rlabel metal2 42280 20888 42280 20888 0 _0612_
rlabel metal2 41832 22512 41832 22512 0 _0613_
rlabel metal2 24248 18480 24248 18480 0 _0614_
rlabel metal2 40264 18648 40264 18648 0 _0615_
rlabel metal2 42168 19656 42168 19656 0 _0616_
rlabel metal2 39592 18704 39592 18704 0 _0617_
rlabel metal3 42000 18424 42000 18424 0 _0618_
rlabel metal2 39704 18872 39704 18872 0 _0619_
rlabel metal2 21560 17696 21560 17696 0 _0620_
rlabel metal2 37800 19208 37800 19208 0 _0621_
rlabel metal3 33656 25256 33656 25256 0 _0622_
rlabel metal2 22680 21952 22680 21952 0 _0623_
rlabel metal3 34496 18648 34496 18648 0 _0624_
rlabel metal3 35280 21560 35280 21560 0 _0625_
rlabel metal2 25368 23576 25368 23576 0 _0626_
rlabel metal2 26376 22736 26376 22736 0 _0627_
rlabel metal2 26824 23464 26824 23464 0 _0628_
rlabel metal2 26768 20104 26768 20104 0 _0629_
rlabel metal3 29680 19992 29680 19992 0 _0630_
rlabel metal3 28896 15960 28896 15960 0 _0631_
rlabel metal2 18312 17136 18312 17136 0 _0632_
rlabel metal2 28280 16800 28280 16800 0 _0633_
rlabel metal2 18760 20832 18760 20832 0 _0634_
rlabel metal2 28504 19376 28504 19376 0 _0635_
rlabel metal2 30072 19992 30072 19992 0 _0636_
rlabel metal3 19936 24024 19936 24024 0 _0637_
rlabel via2 24472 18312 24472 18312 0 _0638_
rlabel metal3 27888 18424 27888 18424 0 _0639_
rlabel metal2 31472 17416 31472 17416 0 _0640_
rlabel metal3 31864 20104 31864 20104 0 _0641_
rlabel metal3 22680 21784 22680 21784 0 _0642_
rlabel metal2 18312 21224 18312 21224 0 _0643_
rlabel metal2 20104 21224 20104 21224 0 _0644_
rlabel metal2 19208 16968 19208 16968 0 _0645_
rlabel metal2 22456 17976 22456 17976 0 _0646_
rlabel metal2 18200 17640 18200 17640 0 _0647_
rlabel metal2 21784 19600 21784 19600 0 _0648_
rlabel metal2 18536 20272 18536 20272 0 _0649_
rlabel metal2 18536 18648 18536 18648 0 _0650_
rlabel metal2 21896 17976 21896 17976 0 _0651_
rlabel metal2 22904 25256 22904 25256 0 _0652_
rlabel metal3 21336 20664 21336 20664 0 _0653_
rlabel metal2 14840 28560 14840 28560 0 _0654_
rlabel metal2 25368 26656 25368 26656 0 _0655_
rlabel metal2 26376 26152 26376 26152 0 _0656_
rlabel metal2 26600 26096 26600 26096 0 _0657_
rlabel metal3 25872 26264 25872 26264 0 _0658_
rlabel metal2 26488 26712 26488 26712 0 _0659_
rlabel metal3 28392 27048 28392 27048 0 _0660_
rlabel metal2 29960 29792 29960 29792 0 _0661_
rlabel metal2 28840 29344 28840 29344 0 _0662_
rlabel metal2 31304 28336 31304 28336 0 _0663_
rlabel metal2 31192 29568 31192 29568 0 _0664_
rlabel metal2 25256 29456 25256 29456 0 _0665_
rlabel metal2 29624 30184 29624 30184 0 _0666_
rlabel metal3 28112 29512 28112 29512 0 _0667_
rlabel metal2 26264 25536 26264 25536 0 _0668_
rlabel metal2 25928 25424 25928 25424 0 _0669_
rlabel metal3 25424 25592 25424 25592 0 _0670_
rlabel metal2 24584 28336 24584 28336 0 _0671_
rlabel metal2 22344 30576 22344 30576 0 _0672_
rlabel metal3 23072 29512 23072 29512 0 _0673_
rlabel metal2 24584 30520 24584 30520 0 _0674_
rlabel metal2 22008 30240 22008 30240 0 _0675_
rlabel metal2 21112 29288 21112 29288 0 _0676_
rlabel metal3 22288 31192 22288 31192 0 _0677_
rlabel metal3 21840 29512 21840 29512 0 _0678_
rlabel metal2 26152 26600 26152 26600 0 _0679_
rlabel metal2 25592 26600 25592 26600 0 _0680_
rlabel metal3 20552 26488 20552 26488 0 _0681_
rlabel metal2 14448 28392 14448 28392 0 _0682_
rlabel metal3 13328 26936 13328 26936 0 _0683_
rlabel metal2 15008 28056 15008 28056 0 _0684_
rlabel metal2 14504 28112 14504 28112 0 _0685_
rlabel metal3 13720 28560 13720 28560 0 _0686_
rlabel metal2 14392 25704 14392 25704 0 _0687_
rlabel metal2 14280 24752 14280 24752 0 _0688_
rlabel metal2 27272 25816 27272 25816 0 _0689_
rlabel metal2 17752 25984 17752 25984 0 _0690_
rlabel metal3 17024 25480 17024 25480 0 _0691_
rlabel metal2 17360 26376 17360 26376 0 _0692_
rlabel metal3 16800 30072 16800 30072 0 _0693_
rlabel metal2 17864 25368 17864 25368 0 _0694_
rlabel metal2 19264 24920 19264 24920 0 _0695_
rlabel metal2 17416 28672 17416 28672 0 _0696_
rlabel metal2 16296 25144 16296 25144 0 _0697_
rlabel metal2 22288 23128 22288 23128 0 _0698_
rlabel metal2 22344 24696 22344 24696 0 _0699_
rlabel metal3 23632 23128 23632 23128 0 _0700_
rlabel metal2 29120 24024 29120 24024 0 _0701_
rlabel metal2 38472 25984 38472 25984 0 _0702_
rlabel metal2 38696 27776 38696 27776 0 _0703_
rlabel metal3 37968 25368 37968 25368 0 _0704_
rlabel metal2 37912 29064 37912 29064 0 _0705_
rlabel metal2 38920 28616 38920 28616 0 _0706_
rlabel metal3 38752 27944 38752 27944 0 _0707_
rlabel metal2 23352 36176 23352 36176 0 _0708_
rlabel metal2 29288 40488 29288 40488 0 _0709_
rlabel metal2 25368 37744 25368 37744 0 _0710_
rlabel metal2 26040 37576 26040 37576 0 _0711_
rlabel metal2 27160 37632 27160 37632 0 _0712_
rlabel metal2 26600 37632 26600 37632 0 _0713_
rlabel metal2 27608 40320 27608 40320 0 _0714_
rlabel metal2 24360 40880 24360 40880 0 _0715_
rlabel metal3 26040 39592 26040 39592 0 _0716_
rlabel metal2 22232 39872 22232 39872 0 _0717_
rlabel metal2 25032 39592 25032 39592 0 _0718_
rlabel metal2 28952 40488 28952 40488 0 _0719_
rlabel metal2 27944 39200 27944 39200 0 _0720_
rlabel metal2 27776 42728 27776 42728 0 _0721_
rlabel metal2 31192 40376 31192 40376 0 _0722_
rlabel metal3 25368 38920 25368 38920 0 _0723_
rlabel metal3 24752 37240 24752 37240 0 _0724_
rlabel metal2 27048 38976 27048 38976 0 _0725_
rlabel metal2 23016 40320 23016 40320 0 _0726_
rlabel metal2 27832 40544 27832 40544 0 _0727_
rlabel metal2 28056 40488 28056 40488 0 _0728_
rlabel metal3 36456 31752 36456 31752 0 _0729_
rlabel metal2 38696 33152 38696 33152 0 _0730_
rlabel metal2 32592 35672 32592 35672 0 _0731_
rlabel metal2 33880 33656 33880 33656 0 _0732_
rlabel metal2 35112 30240 35112 30240 0 _0733_
rlabel metal2 49000 31360 49000 31360 0 _0734_
rlabel metal2 34104 35728 34104 35728 0 _0735_
rlabel metal2 37240 36904 37240 36904 0 _0736_
rlabel metal2 37464 35336 37464 35336 0 _0737_
rlabel metal3 37632 32536 37632 32536 0 _0738_
rlabel metal3 42728 32480 42728 32480 0 _0739_
rlabel metal3 34552 37240 34552 37240 0 _0740_
rlabel metal2 36064 34104 36064 34104 0 _0741_
rlabel metal3 36288 33992 36288 33992 0 _0742_
rlabel metal2 34608 40376 34608 40376 0 _0743_
rlabel metal2 34552 32872 34552 32872 0 _0744_
rlabel metal2 31976 34440 31976 34440 0 _0745_
rlabel metal2 36064 34888 36064 34888 0 _0746_
rlabel metal3 32368 38696 32368 38696 0 _0747_
rlabel metal2 34944 39592 34944 39592 0 _0748_
rlabel metal2 35896 41104 35896 41104 0 _0749_
rlabel metal3 19824 40488 19824 40488 0 _0750_
rlabel metal2 17528 41272 17528 41272 0 _0751_
rlabel metal2 18872 37688 18872 37688 0 _0752_
rlabel metal2 17640 37184 17640 37184 0 _0753_
rlabel metal3 17136 35672 17136 35672 0 _0754_
rlabel metal2 16184 34160 16184 34160 0 _0755_
rlabel metal2 16296 34720 16296 34720 0 _0756_
rlabel metal2 16520 37688 16520 37688 0 _0757_
rlabel metal2 21280 38808 21280 38808 0 _0758_
rlabel metal2 14504 37632 14504 37632 0 _0759_
rlabel metal2 15064 36792 15064 36792 0 _0760_
rlabel metal2 19768 38416 19768 38416 0 _0761_
rlabel metal2 20440 35616 20440 35616 0 _0762_
rlabel metal2 17976 40432 17976 40432 0 _0763_
rlabel metal2 15848 38864 15848 38864 0 _0764_
rlabel metal2 15960 34944 15960 34944 0 _0765_
rlabel metal2 12600 38416 12600 38416 0 _0766_
rlabel metal2 7336 28000 7336 28000 0 _0767_
rlabel metal2 7896 27440 7896 27440 0 _0768_
rlabel metal2 7896 29232 7896 29232 0 _0769_
rlabel metal2 10696 32256 10696 32256 0 _0770_
rlabel metal2 9800 29848 9800 29848 0 _0771_
rlabel metal2 8904 30856 8904 30856 0 _0772_
rlabel metal2 11760 30968 11760 30968 0 _0773_
rlabel metal2 12376 30184 12376 30184 0 _0774_
rlabel metal2 8568 28448 8568 28448 0 _0775_
rlabel metal2 11592 31332 11592 31332 0 _0776_
rlabel metal2 12152 27664 12152 27664 0 _0777_
rlabel metal2 8120 30744 8120 30744 0 _0778_
rlabel metal3 9240 31864 9240 31864 0 _0779_
rlabel metal3 7616 31864 7616 31864 0 _0780_
rlabel metal2 12320 28504 12320 28504 0 _0781_
rlabel metal2 11592 32480 11592 32480 0 _0782_
rlabel metal2 13272 28896 13272 28896 0 _0783_
rlabel metal2 12656 37240 12656 37240 0 _0784_
rlabel metal2 12880 41944 12880 41944 0 _0785_
rlabel metal2 28616 40824 28616 40824 0 _0786_
rlabel metal2 36904 41888 36904 41888 0 _0787_
rlabel metal3 36792 41160 36792 41160 0 _0788_
rlabel metal2 37128 40432 37128 40432 0 _0789_
rlabel metal2 37240 42224 37240 42224 0 _0790_
rlabel metal2 37128 43232 37128 43232 0 _0791_
rlabel metal3 25424 38696 25424 38696 0 _0792_
rlabel metal2 25704 39256 25704 39256 0 _0793_
rlabel metal2 38024 39648 38024 39648 0 _0794_
rlabel metal2 31640 31080 31640 31080 0 _0795_
rlabel metal2 37688 37184 37688 37184 0 _0796_
rlabel metal2 38752 35896 38752 35896 0 _0797_
rlabel metal2 36568 36960 36568 36960 0 _0798_
rlabel metal2 37352 38024 37352 38024 0 _0799_
rlabel metal2 37072 36456 37072 36456 0 _0800_
rlabel metal2 43736 39928 43736 39928 0 _0801_
rlabel metal2 38808 41216 38808 41216 0 _0802_
rlabel metal2 19208 41160 19208 41160 0 _0803_
rlabel metal2 18200 26656 18200 26656 0 _0804_
rlabel metal2 20328 41440 20328 41440 0 _0805_
rlabel metal2 14056 37856 14056 37856 0 _0806_
rlabel metal2 20608 42504 20608 42504 0 _0807_
rlabel metal2 14392 41104 14392 41104 0 _0808_
rlabel metal2 17528 43568 17528 43568 0 _0809_
rlabel metal3 14896 40376 14896 40376 0 _0810_
rlabel metal3 11928 42056 11928 42056 0 _0811_
rlabel metal2 14728 27888 14728 27888 0 _0812_
rlabel metal3 13720 35560 13720 35560 0 _0813_
rlabel metal2 12824 28840 12824 28840 0 _0814_
rlabel metal3 14504 27104 14504 27104 0 _0815_
rlabel metal2 12376 31696 12376 31696 0 _0816_
rlabel metal3 13552 33432 13552 33432 0 _0817_
rlabel metal2 14224 37240 14224 37240 0 _0818_
rlabel metal2 37912 43876 37912 43876 0 _0819_
rlabel metal2 39032 42336 39032 42336 0 _0820_
rlabel metal3 38304 46648 38304 46648 0 _0821_
rlabel metal2 38864 37016 38864 37016 0 _0822_
rlabel metal2 37744 39032 37744 39032 0 _0823_
rlabel metal3 37072 46648 37072 46648 0 _0824_
rlabel metal2 8512 27272 8512 27272 0 _0825_
rlabel metal3 13664 40376 13664 40376 0 _0826_
rlabel metal2 13720 41888 13720 41888 0 _0827_
rlabel metal2 14616 40656 14616 40656 0 _0828_
rlabel metal2 15848 47264 15848 47264 0 _0829_
rlabel metal3 17024 47432 17024 47432 0 _0830_
rlabel metal2 9072 34104 9072 34104 0 _0831_
rlabel metal3 8624 36232 8624 36232 0 _0832_
rlabel metal2 7056 26936 7056 26936 0 _0833_
rlabel metal2 8008 34384 8008 34384 0 _0834_
rlabel metal2 8120 35056 8120 35056 0 _0835_
rlabel metal2 11480 33600 11480 33600 0 _0836_
rlabel metal3 11760 36232 11760 36232 0 _0837_
rlabel metal3 13160 36456 13160 36456 0 _0838_
rlabel metal2 11872 38024 11872 38024 0 _0839_
rlabel metal2 18760 40320 18760 40320 0 _0840_
rlabel metal2 20664 37408 20664 37408 0 _0841_
rlabel metal2 21224 40936 21224 40936 0 _0842_
rlabel metal2 19992 42000 19992 42000 0 _0843_
rlabel metal2 15736 40768 15736 40768 0 _0844_
rlabel metal2 21672 40600 21672 40600 0 _0845_
rlabel metal2 17864 40432 17864 40432 0 _0846_
rlabel metal3 16688 43400 16688 43400 0 _0847_
rlabel metal2 17976 44912 17976 44912 0 _0848_
rlabel metal2 35112 37296 35112 37296 0 _0849_
rlabel metal2 36344 33264 36344 33264 0 _0850_
rlabel metal3 33096 41272 33096 41272 0 _0851_
rlabel metal2 31304 37352 31304 37352 0 _0852_
rlabel metal2 32088 34552 32088 34552 0 _0853_
rlabel metal2 32536 38724 32536 38724 0 _0854_
rlabel metal2 35168 41160 35168 41160 0 _0855_
rlabel via2 25144 41384 25144 41384 0 _0856_
rlabel metal2 27664 41720 27664 41720 0 _0857_
rlabel metal2 26936 41552 26936 41552 0 _0858_
rlabel metal2 25928 41552 25928 41552 0 _0859_
rlabel metal2 28112 41160 28112 41160 0 _0860_
rlabel metal3 28168 42728 28168 42728 0 _0861_
rlabel metal2 24808 44688 24808 44688 0 _0862_
rlabel metal3 21504 46648 21504 46648 0 _0863_
rlabel metal2 35784 46536 35784 46536 0 _0864_
rlabel metal2 36120 47096 36120 47096 0 _0865_
rlabel metal2 36456 47152 36456 47152 0 _0866_
rlabel metal2 37688 47320 37688 47320 0 _0867_
rlabel metal2 18312 47264 18312 47264 0 _0868_
rlabel metal2 31416 44240 31416 44240 0 _0869_
rlabel metal2 24472 44520 24472 44520 0 _0870_
rlabel metal2 24136 45976 24136 45976 0 _0871_
rlabel metal3 30072 46816 30072 46816 0 _0872_
rlabel metal2 35112 34048 35112 34048 0 _0873_
rlabel metal2 32424 34328 32424 34328 0 _0874_
rlabel metal2 33656 34440 33656 34440 0 _0875_
rlabel metal3 28840 45080 28840 45080 0 _0876_
rlabel metal2 27496 40768 27496 40768 0 _0877_
rlabel metal2 24472 40544 24472 40544 0 _0878_
rlabel metal3 27048 38808 27048 38808 0 _0879_
rlabel metal2 26712 40040 26712 40040 0 _0880_
rlabel metal2 27496 46256 27496 46256 0 _0881_
rlabel metal2 27384 47152 27384 47152 0 _0882_
rlabel metal3 14280 32312 14280 32312 0 _0883_
rlabel metal2 13776 33096 13776 33096 0 _0884_
rlabel metal2 14504 45248 14504 45248 0 _0885_
rlabel metal2 15568 44184 15568 44184 0 _0886_
rlabel metal2 18368 42728 18368 42728 0 _0887_
rlabel metal2 20440 41272 20440 41272 0 _0888_
rlabel metal2 14616 43960 14616 43960 0 _0889_
rlabel metal2 26040 46592 26040 46592 0 _0890_
rlabel metal2 15400 44800 15400 44800 0 _0891_
rlabel metal3 14840 45696 14840 45696 0 _0892_
rlabel metal3 16464 45864 16464 45864 0 _0893_
rlabel metal2 27496 47208 27496 47208 0 _0894_
rlabel metal2 35000 47096 35000 47096 0 _0895_
rlabel metal2 36680 47880 36680 47880 0 _0896_
rlabel metal2 35336 47040 35336 47040 0 _0897_
rlabel metal2 37240 49000 37240 49000 0 _0898_
rlabel metal2 27216 48216 27216 48216 0 _0899_
rlabel metal2 29400 47992 29400 47992 0 _0900_
rlabel metal2 27272 47040 27272 47040 0 _0901_
rlabel metal2 27944 48104 27944 48104 0 _0902_
rlabel metal2 27384 48944 27384 48944 0 _0903_
rlabel metal2 28392 43120 28392 43120 0 _0904_
rlabel metal2 31416 49000 31416 49000 0 _0905_
rlabel metal2 30072 38920 30072 38920 0 _0906_
rlabel metal2 32256 49000 32256 49000 0 _0907_
rlabel metal2 32760 49448 32760 49448 0 _0908_
rlabel metal2 14392 45808 14392 45808 0 _0909_
rlabel metal2 10752 50456 10752 50456 0 _0910_
rlabel metal2 15064 49392 15064 49392 0 _0911_
rlabel metal2 16072 46872 16072 46872 0 _0912_
rlabel metal2 13496 47096 13496 47096 0 _0913_
rlabel metal2 11144 48552 11144 48552 0 _0914_
rlabel metal2 16632 47768 16632 47768 0 _0915_
rlabel metal2 16296 47824 16296 47824 0 _0916_
rlabel metal2 33768 49392 33768 49392 0 _0917_
rlabel metal2 35168 49784 35168 49784 0 _0918_
rlabel metal2 38696 50512 38696 50512 0 _0919_
rlabel metal2 38696 51800 38696 51800 0 _0920_
rlabel metal2 35504 50008 35504 50008 0 _0921_
rlabel metal2 36008 53424 36008 53424 0 _0922_
rlabel metal3 31556 49672 31556 49672 0 _0923_
rlabel metal2 28336 49896 28336 49896 0 _0924_
rlabel metal2 33320 49896 33320 49896 0 _0925_
rlabel metal2 35672 52248 35672 52248 0 _0926_
rlabel metal2 28056 42056 28056 42056 0 _0927_
rlabel metal2 30800 50344 30800 50344 0 _0928_
rlabel metal2 30408 39256 30408 39256 0 _0929_
rlabel metal2 32200 40824 32200 40824 0 _0930_
rlabel metal2 33768 52472 33768 52472 0 _0931_
rlabel metal3 14728 51464 14728 51464 0 _0932_
rlabel metal2 15064 51912 15064 51912 0 _0933_
rlabel metal2 14840 37688 14840 37688 0 _0934_
rlabel metal3 13664 51576 13664 51576 0 _0935_
rlabel metal2 10248 37184 10248 37184 0 _0936_
rlabel metal2 9576 35112 9576 35112 0 _0937_
rlabel metal2 8568 37296 8568 37296 0 _0938_
rlabel metal2 9688 51520 9688 51520 0 _0939_
rlabel metal3 14896 52136 14896 52136 0 _0940_
rlabel metal3 15960 52192 15960 52192 0 _0941_
rlabel metal2 15960 52360 15960 52360 0 _0942_
rlabel metal2 16520 52416 16520 52416 0 _0943_
rlabel metal3 36400 52920 36400 52920 0 _0944_
rlabel metal2 36232 53424 36232 53424 0 _0945_
rlabel metal2 42056 54152 42056 54152 0 _0946_
rlabel metal2 30968 32256 30968 32256 0 _0947_
rlabel metal2 29792 34104 29792 34104 0 _0948_
rlabel metal2 29736 35336 29736 35336 0 _0949_
rlabel metal2 31416 34944 31416 34944 0 _0950_
rlabel metal2 30968 50232 30968 50232 0 _0951_
rlabel metal2 26824 37296 26824 37296 0 _0952_
rlabel metal2 29232 40936 29232 40936 0 _0953_
rlabel metal2 29064 41552 29064 41552 0 _0954_
rlabel metal2 28616 42000 28616 42000 0 _0955_
rlabel metal2 29008 42504 29008 42504 0 _0956_
rlabel metal2 29288 45864 29288 45864 0 _0957_
rlabel metal3 32704 55160 32704 55160 0 _0958_
rlabel metal2 18088 44408 18088 44408 0 _0959_
rlabel metal2 21672 42112 21672 42112 0 _0960_
rlabel metal2 18648 44352 18648 44352 0 _0961_
rlabel metal2 11592 51912 11592 51912 0 _0962_
rlabel metal3 11928 37352 11928 37352 0 _0963_
rlabel metal2 8176 34328 8176 34328 0 _0964_
rlabel metal2 9184 37128 9184 37128 0 _0965_
rlabel metal2 7840 38360 7840 38360 0 _0966_
rlabel metal3 15008 54488 15008 54488 0 _0967_
rlabel metal2 12936 52584 12936 52584 0 _0968_
rlabel metal2 15008 54488 15008 54488 0 _0969_
rlabel metal3 20160 54320 20160 54320 0 _0970_
rlabel metal2 34328 55272 34328 55272 0 _0971_
rlabel metal3 20664 53648 20664 53648 0 _0972_
rlabel metal3 28840 54376 28840 54376 0 _0973_
rlabel metal2 32760 52416 32760 52416 0 _0974_
rlabel metal2 33656 54152 33656 54152 0 _0975_
rlabel metal3 35672 56728 35672 56728 0 _0976_
rlabel metal2 36120 53088 36120 53088 0 _0977_
rlabel metal2 36456 53424 36456 53424 0 _0978_
rlabel metal3 38836 56056 38836 56056 0 _0979_
rlabel metal2 42168 57232 42168 57232 0 _0980_
rlabel metal2 36008 56168 36008 56168 0 _0981_
rlabel metal2 36344 57344 36344 57344 0 _0982_
rlabel metal2 30744 55104 30744 55104 0 _0983_
rlabel metal2 24808 53872 24808 53872 0 _0984_
rlabel metal2 31752 55720 31752 55720 0 _0985_
rlabel metal2 32312 55776 32312 55776 0 _0986_
rlabel metal3 34104 56168 34104 56168 0 _0987_
rlabel metal2 11704 36960 11704 36960 0 _0988_
rlabel metal2 13160 52248 13160 52248 0 _0989_
rlabel metal2 15288 39648 15288 39648 0 _0990_
rlabel metal3 15288 55048 15288 55048 0 _0991_
rlabel metal3 13720 56168 13720 56168 0 _0992_
rlabel metal2 6776 59192 6776 59192 0 _0993_
rlabel metal3 12096 60760 12096 60760 0 _0994_
rlabel metal2 13944 56672 13944 56672 0 _0995_
rlabel metal2 14280 56000 14280 56000 0 _0996_
rlabel metal2 11032 55048 11032 55048 0 _0997_
rlabel metal2 6216 56056 6216 56056 0 _0998_
rlabel metal3 12432 55272 12432 55272 0 _0999_
rlabel metal2 14280 54656 14280 54656 0 _1000_
rlabel metal2 14616 54656 14616 54656 0 _1001_
rlabel metal2 26488 57512 26488 57512 0 _1002_
rlabel metal2 23688 41776 23688 41776 0 _1003_
rlabel metal2 25816 56840 25816 56840 0 _1004_
rlabel metal2 30576 38808 30576 38808 0 _1005_
rlabel metal2 25704 57344 25704 57344 0 _1006_
rlabel metal2 26992 56728 26992 56728 0 _1007_
rlabel metal2 27048 58072 27048 58072 0 _1008_
rlabel metal2 36288 58296 36288 58296 0 _1009_
rlabel metal2 39480 58408 39480 58408 0 _1010_
rlabel metal2 35672 60424 35672 60424 0 _1011_
rlabel metal2 36568 57736 36568 57736 0 _1012_
rlabel metal3 38584 62328 38584 62328 0 _1013_
rlabel metal2 23632 55384 23632 55384 0 _1014_
rlabel metal2 25368 58072 25368 58072 0 _1015_
rlabel metal3 26208 58408 26208 58408 0 _1016_
rlabel metal2 34552 61264 34552 61264 0 _1017_
rlabel metal2 31752 46312 31752 46312 0 _1018_
rlabel metal2 27888 60088 27888 60088 0 _1019_
rlabel metal2 27384 49672 27384 49672 0 _1020_
rlabel metal2 28392 60480 28392 60480 0 _1021_
rlabel metal2 25480 60424 25480 60424 0 _1022_
rlabel metal3 28448 59976 28448 59976 0 _1023_
rlabel metal3 28448 60760 28448 60760 0 _1024_
rlabel metal3 15232 57736 15232 57736 0 _1025_
rlabel metal2 13776 59864 13776 59864 0 _1026_
rlabel metal2 12936 53256 12936 53256 0 _1027_
rlabel metal2 8232 52752 8232 52752 0 _1028_
rlabel metal2 4312 53312 4312 53312 0 _1029_
rlabel metal2 12376 52864 12376 52864 0 _1030_
rlabel metal2 12600 51912 12600 51912 0 _1031_
rlabel metal2 5544 50960 5544 50960 0 _1032_
rlabel metal2 12544 52248 12544 52248 0 _1033_
rlabel metal2 13216 52696 13216 52696 0 _1034_
rlabel metal3 14728 56728 14728 56728 0 _1035_
rlabel metal2 15064 57568 15064 57568 0 _1036_
rlabel metal2 15736 60312 15736 60312 0 _1037_
rlabel metal2 34440 61264 34440 61264 0 _1038_
rlabel metal3 38920 62216 38920 62216 0 _1039_
rlabel metal2 41944 62664 41944 62664 0 _1040_
rlabel metal2 35112 60144 35112 60144 0 _1041_
rlabel metal3 36008 59192 36008 59192 0 _1042_
rlabel metal2 37240 60200 37240 60200 0 _1043_
rlabel metal2 34216 60256 34216 60256 0 _1044_
rlabel metal2 36848 43680 36848 43680 0 _1045_
rlabel metal2 31080 49896 31080 49896 0 _1046_
rlabel metal2 33096 59976 33096 59976 0 _1047_
rlabel metal2 26264 56812 26264 56812 0 _1048_
rlabel metal2 15960 59080 15960 59080 0 _1049_
rlabel metal2 16296 60368 16296 60368 0 _1050_
rlabel metal2 18144 60872 18144 60872 0 _1051_
rlabel metal2 16408 61992 16408 61992 0 _1052_
rlabel metal3 17864 59304 17864 59304 0 _1053_
rlabel metal2 16744 59976 16744 59976 0 _1054_
rlabel metal2 7896 62272 7896 62272 0 _1055_
rlabel metal2 13832 57064 13832 57064 0 _1056_
rlabel metal2 14168 58072 14168 58072 0 _1057_
rlabel metal2 17192 59752 17192 59752 0 _1058_
rlabel metal3 20160 60256 20160 60256 0 _1059_
rlabel metal2 34328 60648 34328 60648 0 _1060_
rlabel metal2 37576 61152 37576 61152 0 _1061_
rlabel metal3 46256 62888 46256 62888 0 _1062_
rlabel metal2 32536 63224 32536 63224 0 _1063_
rlabel metal2 24696 58688 24696 58688 0 _1064_
rlabel metal2 32536 60760 32536 60760 0 _1065_
rlabel metal2 32872 60704 32872 60704 0 _1066_
rlabel metal2 37800 61040 37800 61040 0 _1067_
rlabel metal2 17752 59976 17752 59976 0 _1068_
rlabel metal2 25144 60088 25144 60088 0 _1069_
rlabel metal2 38752 62328 38752 62328 0 _1070_
rlabel metal2 34776 60368 34776 60368 0 _1071_
rlabel metal2 38416 62216 38416 62216 0 _1072_
rlabel metal2 53256 62776 53256 62776 0 _1073_
rlabel metal2 39928 61040 39928 61040 0 _1074_
rlabel metal2 51632 57848 51632 57848 0 _1075_
rlabel metal2 52192 51352 52192 51352 0 _1076_
rlabel metal2 54488 49616 54488 49616 0 _1077_
rlabel metal3 51464 51128 51464 51128 0 _1078_
rlabel metal2 51688 53704 51688 53704 0 _1079_
rlabel metal3 30352 9576 30352 9576 0 _1080_
rlabel metal2 40712 25424 40712 25424 0 _1081_
rlabel metal2 39760 26376 39760 26376 0 _1082_
rlabel metal2 29512 25704 29512 25704 0 _1083_
rlabel metal2 26936 25816 26936 25816 0 _1084_
rlabel metal2 24416 23352 24416 23352 0 _1085_
rlabel metal2 34216 24752 34216 24752 0 _1086_
rlabel metal2 32984 19908 32984 19908 0 _1087_
rlabel metal2 31024 5880 31024 5880 0 _1088_
rlabel metal2 31528 10136 31528 10136 0 _1089_
rlabel metal2 30744 10136 30744 10136 0 _1090_
rlabel metal2 35784 24696 35784 24696 0 _1091_
rlabel metal3 24416 29624 24416 29624 0 _1092_
rlabel metal2 46424 21952 46424 21952 0 _1093_
rlabel metal2 57288 11648 57288 11648 0 _1094_
rlabel metal2 18648 24472 18648 24472 0 _1095_
rlabel metal3 46592 19992 46592 19992 0 _1096_
rlabel metal3 24696 19208 24696 19208 0 _1097_
rlabel metal3 23632 9912 23632 9912 0 _1098_
rlabel metal2 42168 8680 42168 8680 0 _1099_
rlabel metal3 31416 8120 31416 8120 0 _1100_
rlabel metal2 14504 25144 14504 25144 0 _1101_
rlabel metal2 42392 18536 42392 18536 0 _1102_
rlabel metal2 30744 5320 30744 5320 0 _1103_
rlabel metal2 14560 24808 14560 24808 0 _1104_
rlabel metal2 45416 20720 45416 20720 0 _1105_
rlabel metal2 31416 6160 31416 6160 0 _1106_
rlabel metal3 47880 4536 47880 4536 0 _1107_
rlabel metal3 39928 25368 39928 25368 0 _1108_
rlabel metal3 40320 26264 40320 26264 0 _1109_
rlabel metal2 40824 24584 40824 24584 0 _1110_
rlabel metal2 43008 6664 43008 6664 0 _1111_
rlabel metal2 43680 7672 43680 7672 0 _1112_
rlabel metal3 46816 5992 46816 5992 0 _1113_
rlabel metal2 46088 8232 46088 8232 0 _1114_
rlabel metal3 45472 17416 45472 17416 0 _1115_
rlabel metal2 45864 4872 45864 4872 0 _1116_
rlabel metal2 43512 6776 43512 6776 0 _1117_
rlabel metal3 48328 21784 48328 21784 0 _1118_
rlabel metal2 39816 25872 39816 25872 0 _1119_
rlabel metal2 44632 23688 44632 23688 0 _1120_
rlabel metal2 45640 22792 45640 22792 0 _1121_
rlabel metal2 47544 19880 47544 19880 0 _1122_
rlabel metal2 47096 22008 47096 22008 0 _1123_
rlabel metal2 47096 18872 47096 18872 0 _1124_
rlabel metal2 46200 19320 46200 19320 0 _1125_
rlabel metal2 7504 38136 7504 38136 0 _1126_
rlabel metal2 40376 41776 40376 41776 0 _1127_
rlabel metal2 46480 22344 46480 22344 0 _1128_
rlabel metal2 41384 40488 41384 40488 0 _1129_
rlabel metal3 49672 45752 49672 45752 0 _1130_
rlabel metal2 48888 39144 48888 39144 0 _1131_
rlabel metal2 24808 12768 24808 12768 0 _1132_
rlabel metal3 39984 38584 39984 38584 0 _1133_
rlabel metal2 40880 36680 40880 36680 0 _1134_
rlabel metal2 39144 37688 39144 37688 0 _1135_
rlabel metal2 39984 37464 39984 37464 0 _1136_
rlabel metal3 36568 42392 36568 42392 0 _1137_
rlabel metal2 22288 44184 22288 44184 0 _1138_
rlabel metal2 22792 43848 22792 43848 0 _1139_
rlabel metal3 50176 46648 50176 46648 0 _1140_
rlabel metal3 46200 47040 46200 47040 0 _1141_
rlabel metal2 22456 52472 22456 52472 0 _1142_
rlabel metal2 22008 44968 22008 44968 0 _1143_
rlabel metal2 23352 45192 23352 45192 0 _1144_
rlabel metal2 22904 46872 22904 46872 0 _1145_
rlabel metal2 22120 49000 22120 49000 0 _1146_
rlabel metal2 24360 47768 24360 47768 0 _1147_
rlabel metal3 24136 47432 24136 47432 0 _1148_
rlabel metal2 21560 48216 21560 48216 0 _1149_
rlabel metal2 20328 49112 20328 49112 0 _1150_
rlabel metal2 20104 48832 20104 48832 0 _1151_
rlabel metal3 21056 48888 21056 48888 0 _1152_
rlabel metal2 19376 49560 19376 49560 0 _1153_
rlabel metal2 21224 49672 21224 49672 0 _1154_
rlabel metal2 19656 53032 19656 53032 0 _1155_
rlabel metal2 18592 53480 18592 53480 0 _1156_
rlabel metal3 4256 52136 4256 52136 0 _1157_
rlabel metal2 17864 53760 17864 53760 0 _1158_
rlabel metal2 20216 52864 20216 52864 0 _1159_
rlabel metal2 20440 53032 20440 53032 0 _1160_
rlabel metal2 23128 52528 23128 52528 0 _1161_
rlabel metal2 22568 52752 22568 52752 0 _1162_
rlabel metal2 23912 53256 23912 53256 0 _1163_
rlabel metal2 24024 53424 24024 53424 0 _1164_
rlabel metal2 23016 56112 23016 56112 0 _1165_
rlabel metal2 22680 56840 22680 56840 0 _1166_
rlabel metal2 23800 56448 23800 56448 0 _1167_
rlabel metal2 24696 57344 24696 57344 0 _1168_
rlabel metal2 24024 59920 24024 59920 0 _1169_
rlabel metal2 23184 59864 23184 59864 0 _1170_
rlabel metal2 2520 46536 2520 46536 0 _1171_
rlabel metal2 25480 61152 25480 61152 0 _1172_
rlabel metal2 26264 60368 26264 60368 0 _1173_
rlabel metal2 25928 60088 25928 60088 0 _1174_
rlabel metal2 20776 57960 20776 57960 0 _1175_
rlabel metal2 18480 55944 18480 55944 0 _1176_
rlabel metal3 19880 57624 19880 57624 0 _1177_
rlabel metal2 20104 57288 20104 57288 0 _1178_
rlabel metal2 3640 37744 3640 37744 0 _1179_
rlabel metal3 3472 37240 3472 37240 0 _1180_
rlabel metal2 4032 41160 4032 41160 0 _1181_
rlabel metal2 2912 39368 2912 39368 0 _1182_
rlabel metal3 4928 39816 4928 39816 0 _1183_
rlabel metal2 5376 41160 5376 41160 0 _1184_
rlabel metal2 3640 41888 3640 41888 0 _1185_
rlabel metal2 4536 44352 4536 44352 0 _1186_
rlabel metal2 5096 44072 5096 44072 0 _1187_
rlabel metal2 3528 44464 3528 44464 0 _1188_
rlabel metal2 2912 42840 2912 42840 0 _1189_
rlabel metal2 4984 44016 4984 44016 0 _1190_
rlabel metal2 4200 45528 4200 45528 0 _1191_
rlabel metal3 3136 46536 3136 46536 0 _1192_
rlabel metal2 5432 47656 5432 47656 0 _1193_
rlabel metal2 5880 48216 5880 48216 0 _1194_
rlabel metal3 4368 50456 4368 50456 0 _1195_
rlabel metal2 5096 51072 5096 51072 0 _1196_
rlabel metal3 4368 51128 4368 51128 0 _1197_
rlabel metal2 4704 50456 4704 50456 0 _1198_
rlabel metal3 4648 50568 4648 50568 0 _1199_
rlabel metal2 5768 51072 5768 51072 0 _1200_
rlabel metal2 5432 53032 5432 53032 0 _1201_
rlabel metal2 3080 55272 3080 55272 0 _1202_
rlabel metal2 4536 55356 4536 55356 0 _1203_
rlabel metal2 3752 55272 3752 55272 0 _1204_
rlabel metal2 4648 53816 4648 53816 0 _1205_
rlabel metal2 5096 54936 5096 54936 0 _1206_
rlabel metal2 4648 56896 4648 56896 0 _1207_
rlabel metal2 4984 58016 4984 58016 0 _1208_
rlabel metal2 4424 56952 4424 56952 0 _1209_
rlabel metal2 48328 45472 48328 45472 0 _1210_
rlabel metal3 7896 59304 7896 59304 0 _1211_
rlabel metal2 6328 57904 6328 57904 0 _1212_
rlabel metal2 6104 57176 6104 57176 0 _1213_
rlabel metal2 7112 59864 7112 59864 0 _1214_
rlabel metal2 7840 59304 7840 59304 0 _1215_
rlabel metal2 6552 60536 6552 60536 0 _1216_
rlabel metal2 7448 60648 7448 60648 0 _1217_
rlabel metal3 6944 62328 6944 62328 0 _1218_
rlabel metal2 8120 62720 8120 62720 0 _1219_
rlabel metal3 7112 63000 7112 63000 0 _1220_
rlabel metal2 7224 62776 7224 62776 0 _1221_
rlabel metal2 8344 62328 8344 62328 0 _1222_
rlabel metal2 9128 62328 9128 62328 0 _1223_
rlabel metal3 14952 62440 14952 62440 0 _1224_
rlabel metal2 18984 60816 18984 60816 0 _1225_
rlabel metal2 19432 62832 19432 62832 0 _1226_
rlabel metal3 43064 24696 43064 24696 0 _1227_
rlabel metal2 20440 62272 20440 62272 0 _1228_
rlabel metal2 19824 62552 19824 62552 0 _1229_
rlabel metal3 10080 38808 10080 38808 0 _1230_
rlabel metal2 6496 38024 6496 38024 0 _1231_
rlabel metal3 9352 41160 9352 41160 0 _1232_
rlabel metal2 8512 40936 8512 40936 0 _1233_
rlabel metal3 9296 42728 9296 42728 0 _1234_
rlabel metal2 9912 42056 9912 42056 0 _1235_
rlabel metal2 10136 44016 10136 44016 0 _1236_
rlabel metal2 8120 45024 8120 45024 0 _1237_
rlabel metal2 9128 52696 9128 52696 0 _1238_
rlabel metal2 8008 44184 8008 44184 0 _1239_
rlabel metal2 9128 46312 9128 46312 0 _1240_
rlabel metal2 9632 45304 9632 45304 0 _1241_
rlabel metal3 10416 47432 10416 47432 0 _1242_
rlabel metal2 12544 46760 12544 46760 0 _1243_
rlabel metal2 11256 48160 11256 48160 0 _1244_
rlabel metal3 12824 47432 12824 47432 0 _1245_
rlabel metal2 9576 48272 9576 48272 0 _1246_
rlabel metal2 8680 48944 8680 48944 0 _1247_
rlabel metal2 8568 48720 8568 48720 0 _1248_
rlabel metal2 8456 48608 8456 48608 0 _1249_
rlabel metal2 9912 49784 9912 49784 0 _1250_
rlabel metal2 9912 50484 9912 50484 0 _1251_
rlabel metal2 7896 53648 7896 53648 0 _1252_
rlabel metal2 7336 52528 7336 52528 0 _1253_
rlabel metal2 7672 53368 7672 53368 0 _1254_
rlabel metal2 8792 52752 8792 52752 0 _1255_
rlabel metal2 8680 53704 8680 53704 0 _1256_
rlabel metal3 8960 57624 8960 57624 0 _1257_
rlabel metal2 8232 57008 8232 57008 0 _1258_
rlabel metal2 30184 44240 30184 44240 0 clknet_0_wb_clk_i
rlabel metal2 21504 4312 21504 4312 0 clknet_4_0_0_wb_clk_i
rlabel metal2 5096 53928 5096 53928 0 clknet_4_10_0_wb_clk_i
rlabel metal2 25368 53424 25368 53424 0 clknet_4_11_0_wb_clk_i
rlabel metal2 44856 47488 44856 47488 0 clknet_4_12_0_wb_clk_i
rlabel metal2 49672 49336 49672 49336 0 clknet_4_13_0_wb_clk_i
rlabel metal2 44408 65408 44408 65408 0 clknet_4_14_0_wb_clk_i
rlabel metal2 55272 53424 55272 53424 0 clknet_4_15_0_wb_clk_i
rlabel metal3 24976 10584 24976 10584 0 clknet_4_1_0_wb_clk_i
rlabel metal2 4760 28224 4760 28224 0 clknet_4_2_0_wb_clk_i
rlabel metal2 19712 24696 19712 24696 0 clknet_4_3_0_wb_clk_i
rlabel metal2 41048 16520 41048 16520 0 clknet_4_4_0_wb_clk_i
rlabel metal2 53368 4648 53368 4648 0 clknet_4_5_0_wb_clk_i
rlabel metal2 41272 22736 41272 22736 0 clknet_4_6_0_wb_clk_i
rlabel metal2 47992 22736 47992 22736 0 clknet_4_7_0_wb_clk_i
rlabel metal2 1848 49000 1848 49000 0 clknet_4_8_0_wb_clk_i
rlabel metal2 25480 50512 25480 50512 0 clknet_4_9_0_wb_clk_i
rlabel metal3 58730 59192 58730 59192 0 custom_settings[0]
rlabel metal2 58184 65800 58184 65800 0 custom_settings[1]
rlabel metal2 58184 3976 58184 3976 0 io_in_1[0]
rlabel metal3 58730 10584 58730 10584 0 io_in_1[1]
rlabel metal3 58730 17528 58730 17528 0 io_in_1[2]
rlabel metal2 58184 24920 58184 24920 0 io_in_1[3]
rlabel metal2 58184 31248 58184 31248 0 io_in_1[4]
rlabel metal3 57904 38696 57904 38696 0 io_in_1[5]
rlabel metal3 58730 45304 58730 45304 0 io_in_1[6]
rlabel metal2 58184 52584 58184 52584 0 io_in_1[7]
rlabel metal3 1246 58296 1246 58296 0 io_in_2
rlabel metal2 22904 67802 22904 67802 0 io_out[10]
rlabel metal3 25536 66472 25536 66472 0 io_out[11]
rlabel metal2 26936 68222 26936 68222 0 io_out[12]
rlabel metal2 37016 67802 37016 67802 0 io_out[17]
rlabel metal3 39928 66472 39928 66472 0 io_out[18]
rlabel metal3 41888 65464 41888 65464 0 io_out[19]
rlabel metal2 43848 66808 43848 66808 0 io_out[20]
rlabel metal3 46760 66472 46760 66472 0 io_out[21]
rlabel metal2 47096 68222 47096 68222 0 io_out[22]
rlabel metal3 50680 66472 50680 66472 0 io_out[23]
rlabel metal3 51128 65520 51128 65520 0 io_out[24]
rlabel metal2 53144 67858 53144 67858 0 io_out[25]
rlabel metal2 55160 66514 55160 66514 0 io_out[26]
rlabel metal2 55384 63112 55384 63112 0 io_out[27]
rlabel metal2 18872 67802 18872 67802 0 io_out[8]
rlabel metal2 20888 68222 20888 68222 0 io_out[9]
rlabel metal2 57792 41944 57792 41944 0 net1
rlabel metal2 52864 47992 52864 47992 0 net10
rlabel metal2 2296 29092 2296 29092 0 net11
rlabel metal2 49784 47712 49784 47712 0 net12
rlabel metal2 23016 64624 23016 64624 0 net13
rlabel metal2 24696 65800 24696 65800 0 net14
rlabel metal2 30296 65128 30296 65128 0 net15
rlabel metal2 51688 49504 51688 49504 0 net16
rlabel metal2 39592 65800 39592 65800 0 net17
rlabel metal2 41384 64736 41384 64736 0 net18
rlabel metal2 46200 64512 46200 64512 0 net19
rlabel metal2 57680 44184 57680 44184 0 net2
rlabel metal2 47432 64204 47432 64204 0 net20
rlabel metal2 49448 63504 49448 63504 0 net21
rlabel metal2 51016 63056 51016 63056 0 net22
rlabel metal3 50456 63896 50456 63896 0 net23
rlabel metal2 50680 63336 50680 63336 0 net24
rlabel metal2 52808 61152 52808 61152 0 net25
rlabel metal3 54040 60760 54040 60760 0 net26
rlabel metal2 17416 65800 17416 65800 0 net27
rlabel metal2 20776 64400 20776 64400 0 net28
rlabel metal2 2744 68222 2744 68222 0 net29
rlabel metal2 54040 5376 54040 5376 0 net3
rlabel metal2 5544 66472 5544 66472 0 net30
rlabel metal2 6776 68222 6776 68222 0 net31
rlabel metal2 9352 66472 9352 66472 0 net32
rlabel metal2 10808 68222 10808 68222 0 net33
rlabel metal2 12824 68222 12824 68222 0 net34
rlabel metal2 14840 68222 14840 68222 0 net35
rlabel metal2 16856 68222 16856 68222 0 net36
rlabel metal2 28952 68222 28952 68222 0 net37
rlabel metal2 30968 68222 30968 68222 0 net38
rlabel metal2 32984 68222 32984 68222 0 net39
rlabel metal2 57624 11256 57624 11256 0 net4
rlabel metal2 35000 68222 35000 68222 0 net40
rlabel metal2 32648 42616 32648 42616 0 net41
rlabel metal2 21504 41944 21504 41944 0 net42
rlabel metal2 14840 39816 14840 39816 0 net43
rlabel metal2 54376 63000 54376 63000 0 net44
rlabel metal3 57176 60872 57176 60872 0 net45
rlabel metal2 15848 44744 15848 44744 0 net46
rlabel metal2 12824 33824 12824 33824 0 net47
rlabel metal2 12600 34944 12600 34944 0 net48
rlabel metal2 39816 42672 39816 42672 0 net49
rlabel metal2 38696 27216 38696 27216 0 net5
rlabel metal2 6552 40712 6552 40712 0 net50
rlabel metal3 5432 39704 5432 39704 0 net51
rlabel metal2 19544 40320 19544 40320 0 net52
rlabel metal2 15624 47320 15624 47320 0 net53
rlabel metal2 10360 35392 10360 35392 0 net54
rlabel metal2 38024 51632 38024 51632 0 net55
rlabel metal2 27832 58128 27832 58128 0 net56
rlabel metal2 9688 41944 9688 41944 0 net57
rlabel metal2 19096 47488 19096 47488 0 net58
rlabel metal2 18872 39592 18872 39592 0 net59
rlabel metal2 57848 25032 57848 25032 0 net6
rlabel metal2 13832 39536 13832 39536 0 net60
rlabel metal3 41048 26488 41048 26488 0 net7
rlabel metal2 35000 25536 35000 25536 0 net8
rlabel metal3 56952 44408 56952 44408 0 net9
rlabel metal3 1302 35000 1302 35000 0 rst_n
rlabel metal3 19880 31752 19880 31752 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
rlabel metal2 19208 25928 19208 25928 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
rlabel metal2 20776 34664 20776 34664 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
rlabel metal2 13832 23856 13832 23856 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
rlabel metal2 19432 34048 19432 34048 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.in
rlabel metal2 7224 29344 7224 29344 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
rlabel metal2 7560 27776 7560 27776 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
rlabel metal2 11368 30576 11368 30576 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
rlabel metal2 13496 26656 13496 26656 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
rlabel metal2 7448 27496 7448 27496 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.in
rlabel metal2 24360 36400 24360 36400 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
rlabel metal2 24024 35336 24024 35336 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
rlabel metal3 24080 37128 24080 37128 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
rlabel metal2 22624 40600 22624 40600 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
rlabel metal2 25480 34776 25480 34776 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.in
rlabel metal3 33768 31752 33768 31752 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
rlabel metal2 31864 32592 31864 32592 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
rlabel metal2 31192 31472 31192 31472 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
rlabel metal2 35224 31808 35224 31808 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
rlabel metal2 41496 32200 41496 32200 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.in
rlabel metal2 56560 39704 56560 39704 0 tt_um_rejunity_sn76489.clk_counter\[0\]
rlabel metal2 55720 46872 55720 46872 0 tt_um_rejunity_sn76489.clk_counter\[1\]
rlabel metal2 55272 45528 55272 45528 0 tt_um_rejunity_sn76489.clk_counter\[2\]
rlabel metal2 55496 44184 55496 44184 0 tt_um_rejunity_sn76489.clk_counter\[3\]
rlabel metal2 51912 44632 51912 44632 0 tt_um_rejunity_sn76489.clk_counter\[4\]
rlabel metal2 52024 42168 52024 42168 0 tt_um_rejunity_sn76489.clk_counter\[5\]
rlabel metal2 53144 39928 53144 39928 0 tt_um_rejunity_sn76489.clk_counter\[6\]
rlabel metal2 38248 25480 38248 25480 0 tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
rlabel metal2 39872 30296 39872 30296 0 tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
rlabel metal2 41496 29008 41496 29008 0 tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
rlabel metal3 29288 9688 29288 9688 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
rlabel metal3 29736 7336 29736 7336 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
rlabel metal2 25144 6440 25144 6440 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
rlabel metal2 21784 5712 21784 5712 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
rlabel metal2 18984 7980 18984 7980 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
rlabel metal2 16856 16912 16856 16912 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
rlabel metal2 18760 19992 18760 19992 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
rlabel metal2 18312 14868 18312 14868 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
rlabel metal2 22792 14420 22792 14420 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
rlabel metal2 22008 20216 22008 20216 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
rlabel metal2 49896 5544 49896 5544 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
rlabel metal3 46984 8232 46984 8232 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
rlabel metal3 47824 4200 47824 4200 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
rlabel metal3 42000 7560 42000 7560 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
rlabel metal2 29512 15512 29512 15512 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
rlabel metal2 30072 13776 30072 13776 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
rlabel metal3 30632 18984 30632 18984 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
rlabel metal2 28728 17864 28728 17864 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
rlabel metal2 32536 16296 32536 16296 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
rlabel metal2 33544 19544 33544 19544 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
rlabel metal2 50904 22456 50904 22456 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
rlabel metal2 49952 19320 49952 19320 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
rlabel metal2 47880 18312 47880 18312 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
rlabel metal2 48216 22736 48216 22736 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
rlabel metal2 44184 22176 44184 22176 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
rlabel metal2 44744 19208 44744 19208 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
rlabel metal2 44296 17808 44296 17808 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
rlabel metal2 40712 16520 40712 16520 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
rlabel metal2 39144 16016 39144 16016 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
rlabel metal2 36456 22512 36456 22512 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
rlabel metal3 7224 38584 7224 38584 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\]
rlabel metal2 9576 42168 9576 42168 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\]
rlabel metal2 8904 45864 8904 45864 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\]
rlabel metal3 10304 48328 10304 48328 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\]
rlabel metal2 8904 48720 8904 48720 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\]
rlabel metal2 8008 52080 8008 52080 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\]
rlabel metal2 10248 57848 10248 57848 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\]
rlabel metal2 11256 60032 11256 60032 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\]
rlabel metal3 11816 64008 11816 64008 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\]
rlabel metal2 16408 63392 16408 63392 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\]
rlabel metal2 3864 36904 3864 36904 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\]
rlabel metal2 5768 40208 5768 40208 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\]
rlabel metal2 4928 45192 4928 45192 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\]
rlabel metal2 5768 47432 5768 47432 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\]
rlabel metal2 4984 50624 4984 50624 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\]
rlabel metal2 4648 54432 4648 54432 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\]
rlabel metal2 5656 57232 5656 57232 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\]
rlabel metal2 6328 60760 6328 60760 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\]
rlabel metal2 8568 64400 8568 64400 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\]
rlabel metal2 20216 60200 20216 60200 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\]
rlabel metal3 41384 40376 41384 40376 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\]
rlabel metal2 39704 37240 39704 37240 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\]
rlabel metal2 21784 45136 21784 45136 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\]
rlabel metal2 24472 48608 24472 48608 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\]
rlabel metal2 19656 50428 19656 50428 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\]
rlabel metal2 20328 52472 20328 52472 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\]
rlabel metal3 23744 53592 23744 53592 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\]
rlabel metal2 24248 56560 24248 56560 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\]
rlabel metal2 24920 60648 24920 60648 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\]
rlabel metal2 20216 56392 20216 56392 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\]
rlabel metal2 45808 38024 45808 38024 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\]
rlabel metal2 47544 39984 47544 39984 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\]
rlabel metal2 31192 44240 31192 44240 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\]
rlabel metal2 29848 46368 29848 46368 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\]
rlabel metal2 28448 50680 28448 50680 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\]
rlabel metal2 28952 54096 28952 54096 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\]
rlabel metal2 30632 57736 30632 57736 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\]
rlabel metal2 27496 64344 27496 64344 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\]
rlabel metal2 31304 63056 31304 63056 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\]
rlabel metal2 33544 64344 33544 64344 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\]
rlabel metal2 23464 24640 23464 24640 0 tt_um_rejunity_sn76489.latch_control_reg\[0\]
rlabel metal2 24472 22736 24472 22736 0 tt_um_rejunity_sn76489.latch_control_reg\[1\]
rlabel metal2 27720 24864 27720 24864 0 tt_um_rejunity_sn76489.latch_control_reg\[2\]
rlabel metal3 45528 25480 45528 25480 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
rlabel metal2 45304 25760 45304 25760 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
rlabel metal3 43736 28392 43736 28392 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
rlabel metal3 44744 31752 44744 31752 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
rlabel metal2 41272 33712 41272 33712 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
rlabel metal2 42728 35000 42728 35000 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
rlabel metal2 45976 33824 45976 33824 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
rlabel metal2 57624 32480 57624 32480 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
rlabel metal2 57960 35896 57960 35896 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
rlabel metal2 56392 35672 56392 35672 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
rlabel metal2 55608 33096 55608 33096 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
rlabel metal2 51240 33096 51240 33096 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
rlabel metal2 50176 29960 50176 29960 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
rlabel metal2 54264 27328 54264 27328 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
rlabel metal2 52584 26152 52584 26152 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
rlabel metal2 53704 23912 53704 23912 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
rlabel metal3 53200 23240 53200 23240 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
rlabel metal2 57848 21504 57848 21504 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
rlabel metal3 55944 23352 55944 23352 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
rlabel metal2 56616 25704 56616 25704 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
rlabel metal3 57568 29624 57568 29624 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
rlabel metal3 49168 28728 49168 28728 0 tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
rlabel metal2 52528 35672 52528 35672 0 tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
rlabel metal3 47544 43400 47544 43400 0 tt_um_rejunity_sn76489.pwm.accumulator\[0\]
rlabel metal3 54600 63224 54600 63224 0 tt_um_rejunity_sn76489.pwm.accumulator\[10\]
rlabel metal2 55272 60592 55272 60592 0 tt_um_rejunity_sn76489.pwm.accumulator\[11\]
rlabel metal2 44072 44296 44072 44296 0 tt_um_rejunity_sn76489.pwm.accumulator\[1\]
rlabel metal2 44856 46928 44856 46928 0 tt_um_rejunity_sn76489.pwm.accumulator\[2\]
rlabel metal2 42616 47712 42616 47712 0 tt_um_rejunity_sn76489.pwm.accumulator\[3\]
rlabel metal3 38192 49896 38192 49896 0 tt_um_rejunity_sn76489.pwm.accumulator\[4\]
rlabel metal2 41496 55160 41496 55160 0 tt_um_rejunity_sn76489.pwm.accumulator\[5\]
rlabel metal2 43176 58352 43176 58352 0 tt_um_rejunity_sn76489.pwm.accumulator\[6\]
rlabel metal2 41384 58800 41384 58800 0 tt_um_rejunity_sn76489.pwm.accumulator\[7\]
rlabel metal3 44632 63000 44632 63000 0 tt_um_rejunity_sn76489.pwm.accumulator\[8\]
rlabel metal2 46536 64232 46536 64232 0 tt_um_rejunity_sn76489.pwm.accumulator\[9\]
rlabel metal2 53704 53144 53704 53144 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\]
rlabel metal2 55384 50120 55384 50120 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
rlabel metal2 57064 51464 57064 51464 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
rlabel metal2 55160 54264 55160 54264 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\]
rlabel metal2 54936 53984 54936 53984 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
rlabel metal2 46816 49112 46816 49112 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
rlabel metal2 54264 59528 54264 59528 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 53984 52920 53984 52920 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 46928 51352 46928 51352 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\]
rlabel metal2 47712 52248 47712 52248 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 46648 53816 46648 53816 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal2 47768 54880 47768 54880 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 48104 56728 48104 56728 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 49896 59640 49896 59640 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal3 50904 62216 50904 62216 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 50792 63896 50792 63896 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 51800 61544 51800 61544 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 24360 7924 24360 7924 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
rlabel metal2 26040 6440 26040 6440 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
rlabel metal2 24472 5432 24472 5432 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
rlabel metal3 21616 5880 21616 5880 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
rlabel metal2 18872 7672 18872 7672 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
rlabel metal3 18984 9800 18984 9800 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
rlabel metal2 18760 11424 18760 11424 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
rlabel metal2 20328 12488 20328 12488 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
rlabel metal2 21672 10416 21672 10416 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
rlabel metal3 26152 14616 26152 14616 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
rlabel metal3 50904 8232 50904 8232 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
rlabel metal2 51464 7112 51464 7112 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
rlabel metal2 51240 6328 51240 6328 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
rlabel metal2 43848 5320 43848 5320 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
rlabel metal2 37128 9464 37128 9464 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
rlabel metal2 35112 5824 35112 5824 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
rlabel metal2 34552 6328 34552 6328 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
rlabel metal2 33320 11704 33320 11704 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
rlabel metal2 38136 11984 38136 11984 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
rlabel metal2 37800 15568 37800 15568 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
rlabel metal2 52136 12432 52136 12432 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
rlabel metal2 53144 18200 53144 18200 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
rlabel metal2 53536 17640 53536 17640 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
rlabel metal2 53592 14784 53592 14784 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
rlabel metal2 52136 14056 52136 14056 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
rlabel metal2 47096 15148 47096 15148 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
rlabel metal2 45696 15288 45696 15288 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
rlabel metal3 45696 15176 45696 15176 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
rlabel metal3 44744 13272 44744 13272 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
rlabel metal3 43232 22456 43232 22456 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
rlabel metal3 1862 11704 1862 11704 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 60000 70000
<< end >>
