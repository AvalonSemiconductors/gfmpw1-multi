VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_ay8913
  CLASS BLOCK ;
  FOREIGN wrapped_ay8913 ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 210.560 250.000 211.120 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 235.200 250.000 235.760 ;
    END
  END custom_settings[1]
  PIN io_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 13.440 250.000 14.000 ;
    END
  END io_in_1[0]
  PIN io_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 38.080 250.000 38.640 ;
    END
  END io_in_1[1]
  PIN io_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 62.720 250.000 63.280 ;
    END
  END io_in_1[2]
  PIN io_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 87.360 250.000 87.920 ;
    END
  END io_in_1[3]
  PIN io_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 112.000 250.000 112.560 ;
    END
  END io_in_1[4]
  PIN io_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 136.640 250.000 137.200 ;
    END
  END io_in_1[5]
  PIN io_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 161.280 250.000 161.840 ;
    END
  END io_in_1[6]
  PIN io_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 185.920 250.000 186.480 ;
    END
  END io_in_1[7]
  PIN io_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 246.000 155.120 250.000 ;
    END
  END io_in_2[0]
  PIN io_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 246.000 216.720 250.000 ;
    END
  END io_in_2[1]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 0.000 18.480 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 0.000 143.920 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 0.000 206.640 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 0.000 222.320 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 246.000 93.520 250.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 246.000 31.920 250.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 229.245 243.470 231.710 ;
        RECT 6.290 229.120 107.905 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 243.470 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 62.200 225.600 ;
        RECT 6.290 221.405 243.470 225.475 ;
        RECT 6.290 221.280 47.640 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 243.470 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 33.425 217.760 ;
        RECT 6.290 213.565 243.470 217.635 ;
        RECT 6.290 213.440 71.505 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 243.470 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 34.545 209.920 ;
        RECT 6.290 205.725 243.470 209.795 ;
        RECT 6.290 205.600 118.200 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 243.470 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 17.960 202.080 ;
        RECT 6.290 197.885 243.470 201.955 ;
        RECT 6.290 197.760 37.905 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 243.470 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 17.960 194.240 ;
        RECT 6.290 190.045 243.470 194.115 ;
        RECT 6.290 189.920 75.985 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 243.470 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 28.945 186.400 ;
        RECT 6.290 182.205 243.470 186.275 ;
        RECT 6.290 182.080 17.960 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 243.470 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 63.880 178.560 ;
        RECT 6.290 174.365 243.470 178.435 ;
        RECT 6.290 174.240 47.465 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 243.470 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 12.705 170.720 ;
        RECT 6.290 166.525 243.470 170.595 ;
        RECT 6.290 166.400 77.320 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 243.470 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 55.825 162.880 ;
        RECT 6.290 158.685 243.470 162.755 ;
        RECT 6.290 158.560 12.705 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 243.470 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 22.225 155.040 ;
        RECT 6.290 150.845 243.470 154.915 ;
        RECT 6.290 150.720 12.705 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 243.470 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 12.705 147.200 ;
        RECT 6.290 143.005 243.470 147.075 ;
        RECT 6.290 142.880 120.225 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 243.470 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 58.625 139.360 ;
        RECT 6.290 135.165 243.470 139.235 ;
        RECT 6.290 135.040 12.705 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 243.470 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 17.960 131.520 ;
        RECT 6.290 127.325 243.470 131.395 ;
        RECT 6.290 127.200 71.505 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 243.470 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 12.705 123.680 ;
        RECT 6.290 119.485 243.470 123.555 ;
        RECT 6.290 119.360 59.400 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 243.470 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 146.760 115.840 ;
        RECT 6.290 111.645 243.470 115.715 ;
        RECT 6.290 111.520 12.705 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 243.470 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 57.505 108.000 ;
        RECT 6.290 103.805 243.470 107.875 ;
        RECT 6.290 103.680 12.705 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 243.470 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 186.305 100.160 ;
        RECT 6.290 95.965 243.470 100.035 ;
        RECT 6.290 95.840 12.705 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 243.470 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 30.625 92.320 ;
        RECT 6.290 88.125 243.470 92.195 ;
        RECT 6.290 88.000 12.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 243.470 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 34.545 84.480 ;
        RECT 6.290 80.285 243.470 84.355 ;
        RECT 6.290 80.160 130.305 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 243.470 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 12.705 76.640 ;
        RECT 6.290 72.445 243.470 76.515 ;
        RECT 6.290 72.320 83.265 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 243.470 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 12.705 68.800 ;
        RECT 6.290 64.605 243.470 68.675 ;
        RECT 6.290 64.480 45.745 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 243.470 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 12.705 60.960 ;
        RECT 6.290 56.765 243.470 60.835 ;
        RECT 6.290 56.640 40.705 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 243.470 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 17.960 53.120 ;
        RECT 6.290 48.925 243.470 52.995 ;
        RECT 6.290 48.800 32.305 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 243.470 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 61.985 45.280 ;
        RECT 6.290 41.085 243.470 45.155 ;
        RECT 6.290 40.960 12.705 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 243.470 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 31.185 37.440 ;
        RECT 6.290 33.245 243.470 37.315 ;
        RECT 6.290 33.120 12.705 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 243.470 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 112.385 29.600 ;
        RECT 6.290 25.405 243.470 29.475 ;
        RECT 6.290 25.280 37.905 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 243.470 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 25.025 21.760 ;
        RECT 6.290 17.565 243.470 21.635 ;
        RECT 6.290 17.440 165.025 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 243.470 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 8.550 243.040 232.250 ;
      LAYER Metal2 ;
        RECT 8.540 245.700 31.060 246.000 ;
        RECT 32.220 245.700 92.660 246.000 ;
        RECT 93.820 245.700 154.260 246.000 ;
        RECT 155.420 245.700 215.860 246.000 ;
        RECT 217.020 245.700 242.900 246.000 ;
        RECT 8.540 4.300 242.900 245.700 ;
        RECT 8.540 3.500 17.620 4.300 ;
        RECT 18.780 3.500 25.460 4.300 ;
        RECT 26.620 3.500 33.300 4.300 ;
        RECT 34.460 3.500 41.140 4.300 ;
        RECT 42.300 3.500 48.980 4.300 ;
        RECT 50.140 3.500 56.820 4.300 ;
        RECT 57.980 3.500 64.660 4.300 ;
        RECT 65.820 3.500 72.500 4.300 ;
        RECT 73.660 3.500 80.340 4.300 ;
        RECT 81.500 3.500 88.180 4.300 ;
        RECT 89.340 3.500 96.020 4.300 ;
        RECT 97.180 3.500 103.860 4.300 ;
        RECT 105.020 3.500 111.700 4.300 ;
        RECT 112.860 3.500 119.540 4.300 ;
        RECT 120.700 3.500 127.380 4.300 ;
        RECT 128.540 3.500 135.220 4.300 ;
        RECT 136.380 3.500 143.060 4.300 ;
        RECT 144.220 3.500 150.900 4.300 ;
        RECT 152.060 3.500 158.740 4.300 ;
        RECT 159.900 3.500 166.580 4.300 ;
        RECT 167.740 3.500 174.420 4.300 ;
        RECT 175.580 3.500 182.260 4.300 ;
        RECT 183.420 3.500 190.100 4.300 ;
        RECT 191.260 3.500 197.940 4.300 ;
        RECT 199.100 3.500 205.780 4.300 ;
        RECT 206.940 3.500 213.620 4.300 ;
        RECT 214.780 3.500 221.460 4.300 ;
        RECT 222.620 3.500 229.300 4.300 ;
        RECT 230.460 3.500 242.900 4.300 ;
      LAYER Metal3 ;
        RECT 8.490 234.900 245.700 235.620 ;
        RECT 8.490 211.420 246.000 234.900 ;
        RECT 8.490 210.260 245.700 211.420 ;
        RECT 8.490 186.780 246.000 210.260 ;
        RECT 8.490 185.620 245.700 186.780 ;
        RECT 8.490 162.140 246.000 185.620 ;
        RECT 8.490 160.980 245.700 162.140 ;
        RECT 8.490 137.500 246.000 160.980 ;
        RECT 8.490 136.340 245.700 137.500 ;
        RECT 8.490 112.860 246.000 136.340 ;
        RECT 8.490 111.700 245.700 112.860 ;
        RECT 8.490 88.220 246.000 111.700 ;
        RECT 8.490 87.060 245.700 88.220 ;
        RECT 8.490 63.580 246.000 87.060 ;
        RECT 8.490 62.420 245.700 63.580 ;
        RECT 8.490 38.940 246.000 62.420 ;
        RECT 8.490 37.780 245.700 38.940 ;
        RECT 8.490 14.300 246.000 37.780 ;
        RECT 8.490 13.140 245.700 14.300 ;
        RECT 8.490 8.540 246.000 13.140 ;
      LAYER Metal4 ;
        RECT 80.220 22.490 98.740 220.550 ;
        RECT 100.940 22.490 175.540 220.550 ;
        RECT 177.740 22.490 235.620 220.550 ;
  END
END wrapped_ay8913
END LIBRARY

